magic
tech sky130A
magscale 1 2
timestamp 1607998557
<< obsli1 >>
rect 1104 2159 158884 157777
<< obsm1 >>
rect 658 1844 159330 157956
<< metal2 >>
rect 662 159200 718 160000
rect 1950 159200 2006 160000
rect 3238 159200 3294 160000
rect 4618 159200 4674 160000
rect 5906 159200 5962 160000
rect 7194 159200 7250 160000
rect 8574 159200 8630 160000
rect 9862 159200 9918 160000
rect 11150 159200 11206 160000
rect 12530 159200 12586 160000
rect 13818 159200 13874 160000
rect 15198 159200 15254 160000
rect 16486 159200 16542 160000
rect 17774 159200 17830 160000
rect 19154 159200 19210 160000
rect 20442 159200 20498 160000
rect 21730 159200 21786 160000
rect 23110 159200 23166 160000
rect 24398 159200 24454 160000
rect 25778 159200 25834 160000
rect 27066 159200 27122 160000
rect 28354 159200 28410 160000
rect 29734 159200 29790 160000
rect 31022 159200 31078 160000
rect 32310 159200 32366 160000
rect 33690 159200 33746 160000
rect 34978 159200 35034 160000
rect 36358 159200 36414 160000
rect 37646 159200 37702 160000
rect 38934 159200 38990 160000
rect 40314 159200 40370 160000
rect 41602 159200 41658 160000
rect 42890 159200 42946 160000
rect 44270 159200 44326 160000
rect 45558 159200 45614 160000
rect 46938 159200 46994 160000
rect 48226 159200 48282 160000
rect 49514 159200 49570 160000
rect 50894 159200 50950 160000
rect 52182 159200 52238 160000
rect 53470 159200 53526 160000
rect 54850 159200 54906 160000
rect 56138 159200 56194 160000
rect 57426 159200 57482 160000
rect 58806 159200 58862 160000
rect 60094 159200 60150 160000
rect 61474 159200 61530 160000
rect 62762 159200 62818 160000
rect 64050 159200 64106 160000
rect 65430 159200 65486 160000
rect 66718 159200 66774 160000
rect 68006 159200 68062 160000
rect 69386 159200 69442 160000
rect 70674 159200 70730 160000
rect 72054 159200 72110 160000
rect 73342 159200 73398 160000
rect 74630 159200 74686 160000
rect 76010 159200 76066 160000
rect 77298 159200 77354 160000
rect 78586 159200 78642 160000
rect 79966 159200 80022 160000
rect 81254 159200 81310 160000
rect 82634 159200 82690 160000
rect 83922 159200 83978 160000
rect 85210 159200 85266 160000
rect 86590 159200 86646 160000
rect 87878 159200 87934 160000
rect 89166 159200 89222 160000
rect 90546 159200 90602 160000
rect 91834 159200 91890 160000
rect 93214 159200 93270 160000
rect 94502 159200 94558 160000
rect 95790 159200 95846 160000
rect 97170 159200 97226 160000
rect 98458 159200 98514 160000
rect 99746 159200 99802 160000
rect 101126 159200 101182 160000
rect 102414 159200 102470 160000
rect 103794 159200 103850 160000
rect 105082 159200 105138 160000
rect 106370 159200 106426 160000
rect 107750 159200 107806 160000
rect 109038 159200 109094 160000
rect 110326 159200 110382 160000
rect 111706 159200 111762 160000
rect 112994 159200 113050 160000
rect 114282 159200 114338 160000
rect 115662 159200 115718 160000
rect 116950 159200 117006 160000
rect 118330 159200 118386 160000
rect 119618 159200 119674 160000
rect 120906 159200 120962 160000
rect 122286 159200 122342 160000
rect 123574 159200 123630 160000
rect 124862 159200 124918 160000
rect 126242 159200 126298 160000
rect 127530 159200 127586 160000
rect 128910 159200 128966 160000
rect 130198 159200 130254 160000
rect 131486 159200 131542 160000
rect 132866 159200 132922 160000
rect 134154 159200 134210 160000
rect 135442 159200 135498 160000
rect 136822 159200 136878 160000
rect 138110 159200 138166 160000
rect 139490 159200 139546 160000
rect 140778 159200 140834 160000
rect 142066 159200 142122 160000
rect 143446 159200 143502 160000
rect 144734 159200 144790 160000
rect 146022 159200 146078 160000
rect 147402 159200 147458 160000
rect 148690 159200 148746 160000
rect 150070 159200 150126 160000
rect 151358 159200 151414 160000
rect 152646 159200 152702 160000
rect 154026 159200 154082 160000
rect 155314 159200 155370 160000
rect 156602 159200 156658 160000
rect 157982 159200 158038 160000
rect 159270 159200 159326 160000
rect 110 0 166 800
rect 386 0 442 800
rect 662 0 718 800
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 1950 0 2006 800
rect 2318 0 2374 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 19062 0 19118 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24766 0 24822 800
rect 25134 0 25190 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37002 0 37058 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42430 0 42486 800
rect 42798 0 42854 800
rect 43074 0 43130 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 44086 0 44142 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 46018 0 46074 800
rect 46294 0 46350 800
rect 46662 0 46718 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48226 0 48282 800
rect 48594 0 48650 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49882 0 49938 800
rect 50158 0 50214 800
rect 50526 0 50582 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51814 0 51870 800
rect 52090 0 52146 800
rect 52458 0 52514 800
rect 52734 0 52790 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53746 0 53802 800
rect 54022 0 54078 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 55954 0 56010 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57610 0 57666 800
rect 57886 0 57942 800
rect 58254 0 58310 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59174 0 59230 800
rect 59542 0 59598 800
rect 59818 0 59874 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60738 0 60794 800
rect 61106 0 61162 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62670 0 62726 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65246 0 65302 800
rect 65614 0 65670 800
rect 65890 0 65946 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 67822 0 67878 800
rect 68190 0 68246 800
rect 68466 0 68522 800
rect 68834 0 68890 800
rect 69110 0 69166 800
rect 69478 0 69534 800
rect 69754 0 69810 800
rect 70122 0 70178 800
rect 70398 0 70454 800
rect 70766 0 70822 800
rect 71042 0 71098 800
rect 71410 0 71466 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 72974 0 73030 800
rect 73342 0 73398 800
rect 73618 0 73674 800
rect 73986 0 74042 800
rect 74262 0 74318 800
rect 74630 0 74686 800
rect 74906 0 74962 800
rect 75274 0 75330 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76562 0 76618 800
rect 76838 0 76894 800
rect 77206 0 77262 800
rect 77482 0 77538 800
rect 77850 0 77906 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78770 0 78826 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79782 0 79838 800
rect 80058 0 80114 800
rect 80334 0 80390 800
rect 80702 0 80758 800
rect 80978 0 81034 800
rect 81346 0 81402 800
rect 81622 0 81678 800
rect 81990 0 82046 800
rect 82266 0 82322 800
rect 82634 0 82690 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83554 0 83610 800
rect 83922 0 83978 800
rect 84198 0 84254 800
rect 84566 0 84622 800
rect 84842 0 84898 800
rect 85210 0 85266 800
rect 85486 0 85542 800
rect 85854 0 85910 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86774 0 86830 800
rect 87142 0 87198 800
rect 87418 0 87474 800
rect 87786 0 87842 800
rect 88062 0 88118 800
rect 88430 0 88486 800
rect 88706 0 88762 800
rect 89074 0 89130 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 89994 0 90050 800
rect 90362 0 90418 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91282 0 91338 800
rect 91650 0 91706 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92570 0 92626 800
rect 92938 0 92994 800
rect 93214 0 93270 800
rect 93582 0 93638 800
rect 93858 0 93914 800
rect 94226 0 94282 800
rect 94502 0 94558 800
rect 94870 0 94926 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 96158 0 96214 800
rect 96434 0 96490 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100298 0 100354 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101218 0 101274 800
rect 101586 0 101642 800
rect 101862 0 101918 800
rect 102230 0 102286 800
rect 102506 0 102562 800
rect 102874 0 102930 800
rect 103150 0 103206 800
rect 103518 0 103574 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105726 0 105782 800
rect 106094 0 106150 800
rect 106370 0 106426 800
rect 106738 0 106794 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107658 0 107714 800
rect 108026 0 108082 800
rect 108302 0 108358 800
rect 108670 0 108726 800
rect 108946 0 109002 800
rect 109314 0 109370 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110878 0 110934 800
rect 111246 0 111302 800
rect 111522 0 111578 800
rect 111890 0 111946 800
rect 112166 0 112222 800
rect 112534 0 112590 800
rect 112810 0 112866 800
rect 113178 0 113234 800
rect 113454 0 113510 800
rect 113822 0 113878 800
rect 114098 0 114154 800
rect 114466 0 114522 800
rect 114742 0 114798 800
rect 115110 0 115166 800
rect 115386 0 115442 800
rect 115754 0 115810 800
rect 116030 0 116086 800
rect 116398 0 116454 800
rect 116674 0 116730 800
rect 117042 0 117098 800
rect 117318 0 117374 800
rect 117686 0 117742 800
rect 117962 0 118018 800
rect 118330 0 118386 800
rect 118606 0 118662 800
rect 118974 0 119030 800
rect 119250 0 119306 800
rect 119618 0 119674 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120814 0 120870 800
rect 121182 0 121238 800
rect 121458 0 121514 800
rect 121826 0 121882 800
rect 122102 0 122158 800
rect 122470 0 122526 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123390 0 123446 800
rect 123758 0 123814 800
rect 124034 0 124090 800
rect 124402 0 124458 800
rect 124678 0 124734 800
rect 125046 0 125102 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127254 0 127310 800
rect 127622 0 127678 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128542 0 128598 800
rect 128910 0 128966 800
rect 129186 0 129242 800
rect 129554 0 129610 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131118 0 131174 800
rect 131486 0 131542 800
rect 131762 0 131818 800
rect 132130 0 132186 800
rect 132406 0 132462 800
rect 132774 0 132830 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133694 0 133750 800
rect 134062 0 134118 800
rect 134338 0 134394 800
rect 134706 0 134762 800
rect 134982 0 135038 800
rect 135350 0 135406 800
rect 135626 0 135682 800
rect 135994 0 136050 800
rect 136270 0 136326 800
rect 136638 0 136694 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 138846 0 138902 800
rect 139214 0 139270 800
rect 139490 0 139546 800
rect 139858 0 139914 800
rect 140134 0 140190 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141054 0 141110 800
rect 141422 0 141478 800
rect 141698 0 141754 800
rect 142066 0 142122 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143630 0 143686 800
rect 143998 0 144054 800
rect 144274 0 144330 800
rect 144642 0 144698 800
rect 144918 0 144974 800
rect 145286 0 145342 800
rect 145562 0 145618 800
rect 145930 0 145986 800
rect 146206 0 146262 800
rect 146574 0 146630 800
rect 146850 0 146906 800
rect 147218 0 147274 800
rect 147494 0 147550 800
rect 147862 0 147918 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148782 0 148838 800
rect 149150 0 149206 800
rect 149426 0 149482 800
rect 149794 0 149850 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151358 0 151414 800
rect 151726 0 151782 800
rect 152002 0 152058 800
rect 152370 0 152426 800
rect 152646 0 152702 800
rect 153014 0 153070 800
rect 153290 0 153346 800
rect 153658 0 153714 800
rect 153934 0 153990 800
rect 154302 0 154358 800
rect 154578 0 154634 800
rect 154946 0 155002 800
rect 155222 0 155278 800
rect 155590 0 155646 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156510 0 156566 800
rect 156878 0 156934 800
rect 157154 0 157210 800
rect 157522 0 157578 800
rect 157798 0 157854 800
rect 158166 0 158222 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159086 0 159142 800
rect 159454 0 159510 800
rect 159730 0 159786 800
<< obsm2 >>
rect 110 159144 606 159202
rect 774 159144 1894 159202
rect 2062 159144 3182 159202
rect 3350 159144 4562 159202
rect 4730 159144 5850 159202
rect 6018 159144 7138 159202
rect 7306 159144 8518 159202
rect 8686 159144 9806 159202
rect 9974 159144 11094 159202
rect 11262 159144 12474 159202
rect 12642 159144 13762 159202
rect 13930 159144 15142 159202
rect 15310 159144 16430 159202
rect 16598 159144 17718 159202
rect 17886 159144 19098 159202
rect 19266 159144 20386 159202
rect 20554 159144 21674 159202
rect 21842 159144 23054 159202
rect 23222 159144 24342 159202
rect 24510 159144 25722 159202
rect 25890 159144 27010 159202
rect 27178 159144 28298 159202
rect 28466 159144 29678 159202
rect 29846 159144 30966 159202
rect 31134 159144 32254 159202
rect 32422 159144 33634 159202
rect 33802 159144 34922 159202
rect 35090 159144 36302 159202
rect 36470 159144 37590 159202
rect 37758 159144 38878 159202
rect 39046 159144 40258 159202
rect 40426 159144 41546 159202
rect 41714 159144 42834 159202
rect 43002 159144 44214 159202
rect 44382 159144 45502 159202
rect 45670 159144 46882 159202
rect 47050 159144 48170 159202
rect 48338 159144 49458 159202
rect 49626 159144 50838 159202
rect 51006 159144 52126 159202
rect 52294 159144 53414 159202
rect 53582 159144 54794 159202
rect 54962 159144 56082 159202
rect 56250 159144 57370 159202
rect 57538 159144 58750 159202
rect 58918 159144 60038 159202
rect 60206 159144 61418 159202
rect 61586 159144 62706 159202
rect 62874 159144 63994 159202
rect 64162 159144 65374 159202
rect 65542 159144 66662 159202
rect 66830 159144 67950 159202
rect 68118 159144 69330 159202
rect 69498 159144 70618 159202
rect 70786 159144 71998 159202
rect 72166 159144 73286 159202
rect 73454 159144 74574 159202
rect 74742 159144 75954 159202
rect 76122 159144 77242 159202
rect 77410 159144 78530 159202
rect 78698 159144 79910 159202
rect 80078 159144 81198 159202
rect 81366 159144 82578 159202
rect 82746 159144 83866 159202
rect 84034 159144 85154 159202
rect 85322 159144 86534 159202
rect 86702 159144 87822 159202
rect 87990 159144 89110 159202
rect 89278 159144 90490 159202
rect 90658 159144 91778 159202
rect 91946 159144 93158 159202
rect 93326 159144 94446 159202
rect 94614 159144 95734 159202
rect 95902 159144 97114 159202
rect 97282 159144 98402 159202
rect 98570 159144 99690 159202
rect 99858 159144 101070 159202
rect 101238 159144 102358 159202
rect 102526 159144 103738 159202
rect 103906 159144 105026 159202
rect 105194 159144 106314 159202
rect 106482 159144 107694 159202
rect 107862 159144 108982 159202
rect 109150 159144 110270 159202
rect 110438 159144 111650 159202
rect 111818 159144 112938 159202
rect 113106 159144 114226 159202
rect 114394 159144 115606 159202
rect 115774 159144 116894 159202
rect 117062 159144 118274 159202
rect 118442 159144 119562 159202
rect 119730 159144 120850 159202
rect 121018 159144 122230 159202
rect 122398 159144 123518 159202
rect 123686 159144 124806 159202
rect 124974 159144 126186 159202
rect 126354 159144 127474 159202
rect 127642 159144 128854 159202
rect 129022 159144 130142 159202
rect 130310 159144 131430 159202
rect 131598 159144 132810 159202
rect 132978 159144 134098 159202
rect 134266 159144 135386 159202
rect 135554 159144 136766 159202
rect 136934 159144 138054 159202
rect 138222 159144 139434 159202
rect 139602 159144 140722 159202
rect 140890 159144 142010 159202
rect 142178 159144 143390 159202
rect 143558 159144 144678 159202
rect 144846 159144 145966 159202
rect 146134 159144 147346 159202
rect 147514 159144 148634 159202
rect 148802 159144 150014 159202
rect 150182 159144 151302 159202
rect 151470 159144 152590 159202
rect 152758 159144 153970 159202
rect 154138 159144 155258 159202
rect 155426 159144 156546 159202
rect 156714 159144 157926 159202
rect 158094 159144 159214 159202
rect 110 856 159324 159144
rect 222 800 330 856
rect 498 800 606 856
rect 774 800 974 856
rect 1142 800 1250 856
rect 1418 800 1618 856
rect 1786 800 1894 856
rect 2062 800 2262 856
rect 2430 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3182 856
rect 3350 800 3550 856
rect 3718 800 3826 856
rect 3994 800 4194 856
rect 4362 800 4470 856
rect 4638 800 4838 856
rect 5006 800 5114 856
rect 5282 800 5482 856
rect 5650 800 5758 856
rect 5926 800 6126 856
rect 6294 800 6402 856
rect 6570 800 6770 856
rect 6938 800 7046 856
rect 7214 800 7414 856
rect 7582 800 7690 856
rect 7858 800 8058 856
rect 8226 800 8334 856
rect 8502 800 8702 856
rect 8870 800 8978 856
rect 9146 800 9346 856
rect 9514 800 9622 856
rect 9790 800 9990 856
rect 10158 800 10266 856
rect 10434 800 10634 856
rect 10802 800 10910 856
rect 11078 800 11278 856
rect 11446 800 11554 856
rect 11722 800 11922 856
rect 12090 800 12198 856
rect 12366 800 12566 856
rect 12734 800 12842 856
rect 13010 800 13210 856
rect 13378 800 13486 856
rect 13654 800 13854 856
rect 14022 800 14130 856
rect 14298 800 14498 856
rect 14666 800 14774 856
rect 14942 800 15142 856
rect 15310 800 15418 856
rect 15586 800 15786 856
rect 15954 800 16062 856
rect 16230 800 16430 856
rect 16598 800 16706 856
rect 16874 800 17074 856
rect 17242 800 17350 856
rect 17518 800 17718 856
rect 17886 800 17994 856
rect 18162 800 18362 856
rect 18530 800 18638 856
rect 18806 800 19006 856
rect 19174 800 19282 856
rect 19450 800 19650 856
rect 19818 800 19926 856
rect 20094 800 20202 856
rect 20370 800 20570 856
rect 20738 800 20846 856
rect 21014 800 21214 856
rect 21382 800 21490 856
rect 21658 800 21858 856
rect 22026 800 22134 856
rect 22302 800 22502 856
rect 22670 800 22778 856
rect 22946 800 23146 856
rect 23314 800 23422 856
rect 23590 800 23790 856
rect 23958 800 24066 856
rect 24234 800 24434 856
rect 24602 800 24710 856
rect 24878 800 25078 856
rect 25246 800 25354 856
rect 25522 800 25722 856
rect 25890 800 25998 856
rect 26166 800 26366 856
rect 26534 800 26642 856
rect 26810 800 27010 856
rect 27178 800 27286 856
rect 27454 800 27654 856
rect 27822 800 27930 856
rect 28098 800 28298 856
rect 28466 800 28574 856
rect 28742 800 28942 856
rect 29110 800 29218 856
rect 29386 800 29586 856
rect 29754 800 29862 856
rect 30030 800 30230 856
rect 30398 800 30506 856
rect 30674 800 30874 856
rect 31042 800 31150 856
rect 31318 800 31518 856
rect 31686 800 31794 856
rect 31962 800 32162 856
rect 32330 800 32438 856
rect 32606 800 32806 856
rect 32974 800 33082 856
rect 33250 800 33450 856
rect 33618 800 33726 856
rect 33894 800 34094 856
rect 34262 800 34370 856
rect 34538 800 34738 856
rect 34906 800 35014 856
rect 35182 800 35382 856
rect 35550 800 35658 856
rect 35826 800 36026 856
rect 36194 800 36302 856
rect 36470 800 36670 856
rect 36838 800 36946 856
rect 37114 800 37314 856
rect 37482 800 37590 856
rect 37758 800 37958 856
rect 38126 800 38234 856
rect 38402 800 38602 856
rect 38770 800 38878 856
rect 39046 800 39246 856
rect 39414 800 39522 856
rect 39690 800 39890 856
rect 40058 800 40166 856
rect 40334 800 40442 856
rect 40610 800 40810 856
rect 40978 800 41086 856
rect 41254 800 41454 856
rect 41622 800 41730 856
rect 41898 800 42098 856
rect 42266 800 42374 856
rect 42542 800 42742 856
rect 42910 800 43018 856
rect 43186 800 43386 856
rect 43554 800 43662 856
rect 43830 800 44030 856
rect 44198 800 44306 856
rect 44474 800 44674 856
rect 44842 800 44950 856
rect 45118 800 45318 856
rect 45486 800 45594 856
rect 45762 800 45962 856
rect 46130 800 46238 856
rect 46406 800 46606 856
rect 46774 800 46882 856
rect 47050 800 47250 856
rect 47418 800 47526 856
rect 47694 800 47894 856
rect 48062 800 48170 856
rect 48338 800 48538 856
rect 48706 800 48814 856
rect 48982 800 49182 856
rect 49350 800 49458 856
rect 49626 800 49826 856
rect 49994 800 50102 856
rect 50270 800 50470 856
rect 50638 800 50746 856
rect 50914 800 51114 856
rect 51282 800 51390 856
rect 51558 800 51758 856
rect 51926 800 52034 856
rect 52202 800 52402 856
rect 52570 800 52678 856
rect 52846 800 53046 856
rect 53214 800 53322 856
rect 53490 800 53690 856
rect 53858 800 53966 856
rect 54134 800 54334 856
rect 54502 800 54610 856
rect 54778 800 54978 856
rect 55146 800 55254 856
rect 55422 800 55622 856
rect 55790 800 55898 856
rect 56066 800 56266 856
rect 56434 800 56542 856
rect 56710 800 56910 856
rect 57078 800 57186 856
rect 57354 800 57554 856
rect 57722 800 57830 856
rect 57998 800 58198 856
rect 58366 800 58474 856
rect 58642 800 58842 856
rect 59010 800 59118 856
rect 59286 800 59486 856
rect 59654 800 59762 856
rect 59930 800 60038 856
rect 60206 800 60406 856
rect 60574 800 60682 856
rect 60850 800 61050 856
rect 61218 800 61326 856
rect 61494 800 61694 856
rect 61862 800 61970 856
rect 62138 800 62338 856
rect 62506 800 62614 856
rect 62782 800 62982 856
rect 63150 800 63258 856
rect 63426 800 63626 856
rect 63794 800 63902 856
rect 64070 800 64270 856
rect 64438 800 64546 856
rect 64714 800 64914 856
rect 65082 800 65190 856
rect 65358 800 65558 856
rect 65726 800 65834 856
rect 66002 800 66202 856
rect 66370 800 66478 856
rect 66646 800 66846 856
rect 67014 800 67122 856
rect 67290 800 67490 856
rect 67658 800 67766 856
rect 67934 800 68134 856
rect 68302 800 68410 856
rect 68578 800 68778 856
rect 68946 800 69054 856
rect 69222 800 69422 856
rect 69590 800 69698 856
rect 69866 800 70066 856
rect 70234 800 70342 856
rect 70510 800 70710 856
rect 70878 800 70986 856
rect 71154 800 71354 856
rect 71522 800 71630 856
rect 71798 800 71998 856
rect 72166 800 72274 856
rect 72442 800 72642 856
rect 72810 800 72918 856
rect 73086 800 73286 856
rect 73454 800 73562 856
rect 73730 800 73930 856
rect 74098 800 74206 856
rect 74374 800 74574 856
rect 74742 800 74850 856
rect 75018 800 75218 856
rect 75386 800 75494 856
rect 75662 800 75862 856
rect 76030 800 76138 856
rect 76306 800 76506 856
rect 76674 800 76782 856
rect 76950 800 77150 856
rect 77318 800 77426 856
rect 77594 800 77794 856
rect 77962 800 78070 856
rect 78238 800 78438 856
rect 78606 800 78714 856
rect 78882 800 79082 856
rect 79250 800 79358 856
rect 79526 800 79726 856
rect 79894 800 80002 856
rect 80170 800 80278 856
rect 80446 800 80646 856
rect 80814 800 80922 856
rect 81090 800 81290 856
rect 81458 800 81566 856
rect 81734 800 81934 856
rect 82102 800 82210 856
rect 82378 800 82578 856
rect 82746 800 82854 856
rect 83022 800 83222 856
rect 83390 800 83498 856
rect 83666 800 83866 856
rect 84034 800 84142 856
rect 84310 800 84510 856
rect 84678 800 84786 856
rect 84954 800 85154 856
rect 85322 800 85430 856
rect 85598 800 85798 856
rect 85966 800 86074 856
rect 86242 800 86442 856
rect 86610 800 86718 856
rect 86886 800 87086 856
rect 87254 800 87362 856
rect 87530 800 87730 856
rect 87898 800 88006 856
rect 88174 800 88374 856
rect 88542 800 88650 856
rect 88818 800 89018 856
rect 89186 800 89294 856
rect 89462 800 89662 856
rect 89830 800 89938 856
rect 90106 800 90306 856
rect 90474 800 90582 856
rect 90750 800 90950 856
rect 91118 800 91226 856
rect 91394 800 91594 856
rect 91762 800 91870 856
rect 92038 800 92238 856
rect 92406 800 92514 856
rect 92682 800 92882 856
rect 93050 800 93158 856
rect 93326 800 93526 856
rect 93694 800 93802 856
rect 93970 800 94170 856
rect 94338 800 94446 856
rect 94614 800 94814 856
rect 94982 800 95090 856
rect 95258 800 95458 856
rect 95626 800 95734 856
rect 95902 800 96102 856
rect 96270 800 96378 856
rect 96546 800 96746 856
rect 96914 800 97022 856
rect 97190 800 97390 856
rect 97558 800 97666 856
rect 97834 800 98034 856
rect 98202 800 98310 856
rect 98478 800 98678 856
rect 98846 800 98954 856
rect 99122 800 99322 856
rect 99490 800 99598 856
rect 99766 800 99966 856
rect 100134 800 100242 856
rect 100410 800 100518 856
rect 100686 800 100886 856
rect 101054 800 101162 856
rect 101330 800 101530 856
rect 101698 800 101806 856
rect 101974 800 102174 856
rect 102342 800 102450 856
rect 102618 800 102818 856
rect 102986 800 103094 856
rect 103262 800 103462 856
rect 103630 800 103738 856
rect 103906 800 104106 856
rect 104274 800 104382 856
rect 104550 800 104750 856
rect 104918 800 105026 856
rect 105194 800 105394 856
rect 105562 800 105670 856
rect 105838 800 106038 856
rect 106206 800 106314 856
rect 106482 800 106682 856
rect 106850 800 106958 856
rect 107126 800 107326 856
rect 107494 800 107602 856
rect 107770 800 107970 856
rect 108138 800 108246 856
rect 108414 800 108614 856
rect 108782 800 108890 856
rect 109058 800 109258 856
rect 109426 800 109534 856
rect 109702 800 109902 856
rect 110070 800 110178 856
rect 110346 800 110546 856
rect 110714 800 110822 856
rect 110990 800 111190 856
rect 111358 800 111466 856
rect 111634 800 111834 856
rect 112002 800 112110 856
rect 112278 800 112478 856
rect 112646 800 112754 856
rect 112922 800 113122 856
rect 113290 800 113398 856
rect 113566 800 113766 856
rect 113934 800 114042 856
rect 114210 800 114410 856
rect 114578 800 114686 856
rect 114854 800 115054 856
rect 115222 800 115330 856
rect 115498 800 115698 856
rect 115866 800 115974 856
rect 116142 800 116342 856
rect 116510 800 116618 856
rect 116786 800 116986 856
rect 117154 800 117262 856
rect 117430 800 117630 856
rect 117798 800 117906 856
rect 118074 800 118274 856
rect 118442 800 118550 856
rect 118718 800 118918 856
rect 119086 800 119194 856
rect 119362 800 119562 856
rect 119730 800 119838 856
rect 120006 800 120114 856
rect 120282 800 120482 856
rect 120650 800 120758 856
rect 120926 800 121126 856
rect 121294 800 121402 856
rect 121570 800 121770 856
rect 121938 800 122046 856
rect 122214 800 122414 856
rect 122582 800 122690 856
rect 122858 800 123058 856
rect 123226 800 123334 856
rect 123502 800 123702 856
rect 123870 800 123978 856
rect 124146 800 124346 856
rect 124514 800 124622 856
rect 124790 800 124990 856
rect 125158 800 125266 856
rect 125434 800 125634 856
rect 125802 800 125910 856
rect 126078 800 126278 856
rect 126446 800 126554 856
rect 126722 800 126922 856
rect 127090 800 127198 856
rect 127366 800 127566 856
rect 127734 800 127842 856
rect 128010 800 128210 856
rect 128378 800 128486 856
rect 128654 800 128854 856
rect 129022 800 129130 856
rect 129298 800 129498 856
rect 129666 800 129774 856
rect 129942 800 130142 856
rect 130310 800 130418 856
rect 130586 800 130786 856
rect 130954 800 131062 856
rect 131230 800 131430 856
rect 131598 800 131706 856
rect 131874 800 132074 856
rect 132242 800 132350 856
rect 132518 800 132718 856
rect 132886 800 132994 856
rect 133162 800 133362 856
rect 133530 800 133638 856
rect 133806 800 134006 856
rect 134174 800 134282 856
rect 134450 800 134650 856
rect 134818 800 134926 856
rect 135094 800 135294 856
rect 135462 800 135570 856
rect 135738 800 135938 856
rect 136106 800 136214 856
rect 136382 800 136582 856
rect 136750 800 136858 856
rect 137026 800 137226 856
rect 137394 800 137502 856
rect 137670 800 137870 856
rect 138038 800 138146 856
rect 138314 800 138514 856
rect 138682 800 138790 856
rect 138958 800 139158 856
rect 139326 800 139434 856
rect 139602 800 139802 856
rect 139970 800 140078 856
rect 140246 800 140354 856
rect 140522 800 140722 856
rect 140890 800 140998 856
rect 141166 800 141366 856
rect 141534 800 141642 856
rect 141810 800 142010 856
rect 142178 800 142286 856
rect 142454 800 142654 856
rect 142822 800 142930 856
rect 143098 800 143298 856
rect 143466 800 143574 856
rect 143742 800 143942 856
rect 144110 800 144218 856
rect 144386 800 144586 856
rect 144754 800 144862 856
rect 145030 800 145230 856
rect 145398 800 145506 856
rect 145674 800 145874 856
rect 146042 800 146150 856
rect 146318 800 146518 856
rect 146686 800 146794 856
rect 146962 800 147162 856
rect 147330 800 147438 856
rect 147606 800 147806 856
rect 147974 800 148082 856
rect 148250 800 148450 856
rect 148618 800 148726 856
rect 148894 800 149094 856
rect 149262 800 149370 856
rect 149538 800 149738 856
rect 149906 800 150014 856
rect 150182 800 150382 856
rect 150550 800 150658 856
rect 150826 800 151026 856
rect 151194 800 151302 856
rect 151470 800 151670 856
rect 151838 800 151946 856
rect 152114 800 152314 856
rect 152482 800 152590 856
rect 152758 800 152958 856
rect 153126 800 153234 856
rect 153402 800 153602 856
rect 153770 800 153878 856
rect 154046 800 154246 856
rect 154414 800 154522 856
rect 154690 800 154890 856
rect 155058 800 155166 856
rect 155334 800 155534 856
rect 155702 800 155810 856
rect 155978 800 156178 856
rect 156346 800 156454 856
rect 156622 800 156822 856
rect 156990 800 157098 856
rect 157266 800 157466 856
rect 157634 800 157742 856
rect 157910 800 158110 856
rect 158278 800 158386 856
rect 158554 800 158754 856
rect 158922 800 159030 856
rect 159198 800 159324 856
<< metal3 >>
rect 0 151784 800 151904
rect 159200 146616 160000 146736
rect 0 135736 800 135856
rect 0 119824 800 119944
rect 159200 119960 160000 120080
rect 0 103776 800 103896
rect 159200 93304 160000 93424
rect 0 87864 800 87984
rect 0 71816 800 71936
rect 159200 66648 160000 66768
rect 0 55768 800 55888
rect 0 39856 800 39976
rect 159200 39992 160000 40112
rect 0 23808 800 23928
rect 159200 13336 160000 13456
rect 0 7896 800 8016
<< obsm3 >>
rect 105 151984 159200 157793
rect 880 151704 159200 151984
rect 105 146816 159200 151704
rect 105 146536 159120 146816
rect 105 135936 159200 146536
rect 880 135656 159200 135936
rect 105 120160 159200 135656
rect 105 120024 159120 120160
rect 880 119880 159120 120024
rect 880 119744 159200 119880
rect 105 103976 159200 119744
rect 880 103696 159200 103976
rect 105 93504 159200 103696
rect 105 93224 159120 93504
rect 105 88064 159200 93224
rect 880 87784 159200 88064
rect 105 72016 159200 87784
rect 880 71736 159200 72016
rect 105 66848 159200 71736
rect 105 66568 159120 66848
rect 105 55968 159200 66568
rect 880 55688 159200 55968
rect 105 40192 159200 55688
rect 105 40056 159120 40192
rect 880 39912 159120 40056
rect 880 39776 159200 39912
rect 105 24008 159200 39776
rect 880 23728 159200 24008
rect 105 13536 159200 23728
rect 105 13256 159120 13536
rect 105 8096 159200 13256
rect 880 7816 159200 8096
rect 105 2143 159200 7816
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
<< obsm4 >>
rect 26371 2128 158128 157808
<< labels >>
rlabel metal2 s 151358 159200 151414 160000 6 analog_io[0]
port 1 nsew default bidirectional
rlabel metal2 s 158166 0 158222 800 6 analog_io[10]
port 2 nsew default bidirectional
rlabel metal3 s 159200 39992 160000 40112 6 analog_io[11]
port 3 nsew default bidirectional
rlabel metal2 s 155314 159200 155370 160000 6 analog_io[12]
port 4 nsew default bidirectional
rlabel metal2 s 158442 0 158498 800 6 analog_io[13]
port 5 nsew default bidirectional
rlabel metal3 s 159200 66648 160000 66768 6 analog_io[14]
port 6 nsew default bidirectional
rlabel metal2 s 158810 0 158866 800 6 analog_io[15]
port 7 nsew default bidirectional
rlabel metal2 s 156602 159200 156658 160000 6 analog_io[16]
port 8 nsew default bidirectional
rlabel metal2 s 159086 0 159142 800 6 analog_io[17]
port 9 nsew default bidirectional
rlabel metal2 s 159454 0 159510 800 6 analog_io[18]
port 10 nsew default bidirectional
rlabel metal3 s 0 71816 800 71936 6 analog_io[19]
port 11 nsew default bidirectional
rlabel metal3 s 0 7896 800 8016 6 analog_io[1]
port 12 nsew default bidirectional
rlabel metal3 s 159200 93304 160000 93424 6 analog_io[20]
port 13 nsew default bidirectional
rlabel metal2 s 159730 0 159786 800 6 analog_io[21]
port 14 nsew default bidirectional
rlabel metal2 s 157982 159200 158038 160000 6 analog_io[22]
port 15 nsew default bidirectional
rlabel metal3 s 0 87864 800 87984 6 analog_io[23]
port 16 nsew default bidirectional
rlabel metal2 s 159270 159200 159326 160000 6 analog_io[24]
port 17 nsew default bidirectional
rlabel metal3 s 159200 119960 160000 120080 6 analog_io[25]
port 18 nsew default bidirectional
rlabel metal3 s 0 103776 800 103896 6 analog_io[26]
port 19 nsew default bidirectional
rlabel metal3 s 0 119824 800 119944 6 analog_io[27]
port 20 nsew default bidirectional
rlabel metal3 s 159200 146616 160000 146736 6 analog_io[28]
port 21 nsew default bidirectional
rlabel metal3 s 0 135736 800 135856 6 analog_io[29]
port 22 nsew default bidirectional
rlabel metal3 s 159200 13336 160000 13456 6 analog_io[2]
port 23 nsew default bidirectional
rlabel metal3 s 0 151784 800 151904 6 analog_io[30]
port 24 nsew default bidirectional
rlabel metal2 s 157522 0 157578 800 6 analog_io[3]
port 25 nsew default bidirectional
rlabel metal3 s 0 23808 800 23928 6 analog_io[4]
port 26 nsew default bidirectional
rlabel metal2 s 152646 159200 152702 160000 6 analog_io[5]
port 27 nsew default bidirectional
rlabel metal3 s 0 39856 800 39976 6 analog_io[6]
port 28 nsew default bidirectional
rlabel metal2 s 157798 0 157854 800 6 analog_io[7]
port 29 nsew default bidirectional
rlabel metal3 s 0 55768 800 55888 6 analog_io[8]
port 30 nsew default bidirectional
rlabel metal2 s 154026 159200 154082 160000 6 analog_io[9]
port 31 nsew default bidirectional
rlabel metal2 s 662 159200 718 160000 6 io_in[0]
port 32 nsew default input
rlabel metal2 s 40314 159200 40370 160000 6 io_in[10]
port 33 nsew default input
rlabel metal2 s 44270 159200 44326 160000 6 io_in[11]
port 34 nsew default input
rlabel metal2 s 48226 159200 48282 160000 6 io_in[12]
port 35 nsew default input
rlabel metal2 s 52182 159200 52238 160000 6 io_in[13]
port 36 nsew default input
rlabel metal2 s 56138 159200 56194 160000 6 io_in[14]
port 37 nsew default input
rlabel metal2 s 60094 159200 60150 160000 6 io_in[15]
port 38 nsew default input
rlabel metal2 s 64050 159200 64106 160000 6 io_in[16]
port 39 nsew default input
rlabel metal2 s 68006 159200 68062 160000 6 io_in[17]
port 40 nsew default input
rlabel metal2 s 72054 159200 72110 160000 6 io_in[18]
port 41 nsew default input
rlabel metal2 s 76010 159200 76066 160000 6 io_in[19]
port 42 nsew default input
rlabel metal2 s 4618 159200 4674 160000 6 io_in[1]
port 43 nsew default input
rlabel metal2 s 79966 159200 80022 160000 6 io_in[20]
port 44 nsew default input
rlabel metal2 s 83922 159200 83978 160000 6 io_in[21]
port 45 nsew default input
rlabel metal2 s 87878 159200 87934 160000 6 io_in[22]
port 46 nsew default input
rlabel metal2 s 91834 159200 91890 160000 6 io_in[23]
port 47 nsew default input
rlabel metal2 s 95790 159200 95846 160000 6 io_in[24]
port 48 nsew default input
rlabel metal2 s 99746 159200 99802 160000 6 io_in[25]
port 49 nsew default input
rlabel metal2 s 103794 159200 103850 160000 6 io_in[26]
port 50 nsew default input
rlabel metal2 s 107750 159200 107806 160000 6 io_in[27]
port 51 nsew default input
rlabel metal2 s 111706 159200 111762 160000 6 io_in[28]
port 52 nsew default input
rlabel metal2 s 115662 159200 115718 160000 6 io_in[29]
port 53 nsew default input
rlabel metal2 s 8574 159200 8630 160000 6 io_in[2]
port 54 nsew default input
rlabel metal2 s 119618 159200 119674 160000 6 io_in[30]
port 55 nsew default input
rlabel metal2 s 123574 159200 123630 160000 6 io_in[31]
port 56 nsew default input
rlabel metal2 s 127530 159200 127586 160000 6 io_in[32]
port 57 nsew default input
rlabel metal2 s 131486 159200 131542 160000 6 io_in[33]
port 58 nsew default input
rlabel metal2 s 135442 159200 135498 160000 6 io_in[34]
port 59 nsew default input
rlabel metal2 s 139490 159200 139546 160000 6 io_in[35]
port 60 nsew default input
rlabel metal2 s 143446 159200 143502 160000 6 io_in[36]
port 61 nsew default input
rlabel metal2 s 147402 159200 147458 160000 6 io_in[37]
port 62 nsew default input
rlabel metal2 s 12530 159200 12586 160000 6 io_in[3]
port 63 nsew default input
rlabel metal2 s 16486 159200 16542 160000 6 io_in[4]
port 64 nsew default input
rlabel metal2 s 20442 159200 20498 160000 6 io_in[5]
port 65 nsew default input
rlabel metal2 s 24398 159200 24454 160000 6 io_in[6]
port 66 nsew default input
rlabel metal2 s 28354 159200 28410 160000 6 io_in[7]
port 67 nsew default input
rlabel metal2 s 32310 159200 32366 160000 6 io_in[8]
port 68 nsew default input
rlabel metal2 s 36358 159200 36414 160000 6 io_in[9]
port 69 nsew default input
rlabel metal2 s 1950 159200 2006 160000 6 io_oeb[0]
port 70 nsew default output
rlabel metal2 s 41602 159200 41658 160000 6 io_oeb[10]
port 71 nsew default output
rlabel metal2 s 45558 159200 45614 160000 6 io_oeb[11]
port 72 nsew default output
rlabel metal2 s 49514 159200 49570 160000 6 io_oeb[12]
port 73 nsew default output
rlabel metal2 s 53470 159200 53526 160000 6 io_oeb[13]
port 74 nsew default output
rlabel metal2 s 57426 159200 57482 160000 6 io_oeb[14]
port 75 nsew default output
rlabel metal2 s 61474 159200 61530 160000 6 io_oeb[15]
port 76 nsew default output
rlabel metal2 s 65430 159200 65486 160000 6 io_oeb[16]
port 77 nsew default output
rlabel metal2 s 69386 159200 69442 160000 6 io_oeb[17]
port 78 nsew default output
rlabel metal2 s 73342 159200 73398 160000 6 io_oeb[18]
port 79 nsew default output
rlabel metal2 s 77298 159200 77354 160000 6 io_oeb[19]
port 80 nsew default output
rlabel metal2 s 5906 159200 5962 160000 6 io_oeb[1]
port 81 nsew default output
rlabel metal2 s 81254 159200 81310 160000 6 io_oeb[20]
port 82 nsew default output
rlabel metal2 s 85210 159200 85266 160000 6 io_oeb[21]
port 83 nsew default output
rlabel metal2 s 89166 159200 89222 160000 6 io_oeb[22]
port 84 nsew default output
rlabel metal2 s 93214 159200 93270 160000 6 io_oeb[23]
port 85 nsew default output
rlabel metal2 s 97170 159200 97226 160000 6 io_oeb[24]
port 86 nsew default output
rlabel metal2 s 101126 159200 101182 160000 6 io_oeb[25]
port 87 nsew default output
rlabel metal2 s 105082 159200 105138 160000 6 io_oeb[26]
port 88 nsew default output
rlabel metal2 s 109038 159200 109094 160000 6 io_oeb[27]
port 89 nsew default output
rlabel metal2 s 112994 159200 113050 160000 6 io_oeb[28]
port 90 nsew default output
rlabel metal2 s 116950 159200 117006 160000 6 io_oeb[29]
port 91 nsew default output
rlabel metal2 s 9862 159200 9918 160000 6 io_oeb[2]
port 92 nsew default output
rlabel metal2 s 120906 159200 120962 160000 6 io_oeb[30]
port 93 nsew default output
rlabel metal2 s 124862 159200 124918 160000 6 io_oeb[31]
port 94 nsew default output
rlabel metal2 s 128910 159200 128966 160000 6 io_oeb[32]
port 95 nsew default output
rlabel metal2 s 132866 159200 132922 160000 6 io_oeb[33]
port 96 nsew default output
rlabel metal2 s 136822 159200 136878 160000 6 io_oeb[34]
port 97 nsew default output
rlabel metal2 s 140778 159200 140834 160000 6 io_oeb[35]
port 98 nsew default output
rlabel metal2 s 144734 159200 144790 160000 6 io_oeb[36]
port 99 nsew default output
rlabel metal2 s 148690 159200 148746 160000 6 io_oeb[37]
port 100 nsew default output
rlabel metal2 s 13818 159200 13874 160000 6 io_oeb[3]
port 101 nsew default output
rlabel metal2 s 17774 159200 17830 160000 6 io_oeb[4]
port 102 nsew default output
rlabel metal2 s 21730 159200 21786 160000 6 io_oeb[5]
port 103 nsew default output
rlabel metal2 s 25778 159200 25834 160000 6 io_oeb[6]
port 104 nsew default output
rlabel metal2 s 29734 159200 29790 160000 6 io_oeb[7]
port 105 nsew default output
rlabel metal2 s 33690 159200 33746 160000 6 io_oeb[8]
port 106 nsew default output
rlabel metal2 s 37646 159200 37702 160000 6 io_oeb[9]
port 107 nsew default output
rlabel metal2 s 3238 159200 3294 160000 6 io_out[0]
port 108 nsew default output
rlabel metal2 s 42890 159200 42946 160000 6 io_out[10]
port 109 nsew default output
rlabel metal2 s 46938 159200 46994 160000 6 io_out[11]
port 110 nsew default output
rlabel metal2 s 50894 159200 50950 160000 6 io_out[12]
port 111 nsew default output
rlabel metal2 s 54850 159200 54906 160000 6 io_out[13]
port 112 nsew default output
rlabel metal2 s 58806 159200 58862 160000 6 io_out[14]
port 113 nsew default output
rlabel metal2 s 62762 159200 62818 160000 6 io_out[15]
port 114 nsew default output
rlabel metal2 s 66718 159200 66774 160000 6 io_out[16]
port 115 nsew default output
rlabel metal2 s 70674 159200 70730 160000 6 io_out[17]
port 116 nsew default output
rlabel metal2 s 74630 159200 74686 160000 6 io_out[18]
port 117 nsew default output
rlabel metal2 s 78586 159200 78642 160000 6 io_out[19]
port 118 nsew default output
rlabel metal2 s 7194 159200 7250 160000 6 io_out[1]
port 119 nsew default output
rlabel metal2 s 82634 159200 82690 160000 6 io_out[20]
port 120 nsew default output
rlabel metal2 s 86590 159200 86646 160000 6 io_out[21]
port 121 nsew default output
rlabel metal2 s 90546 159200 90602 160000 6 io_out[22]
port 122 nsew default output
rlabel metal2 s 94502 159200 94558 160000 6 io_out[23]
port 123 nsew default output
rlabel metal2 s 98458 159200 98514 160000 6 io_out[24]
port 124 nsew default output
rlabel metal2 s 102414 159200 102470 160000 6 io_out[25]
port 125 nsew default output
rlabel metal2 s 106370 159200 106426 160000 6 io_out[26]
port 126 nsew default output
rlabel metal2 s 110326 159200 110382 160000 6 io_out[27]
port 127 nsew default output
rlabel metal2 s 114282 159200 114338 160000 6 io_out[28]
port 128 nsew default output
rlabel metal2 s 118330 159200 118386 160000 6 io_out[29]
port 129 nsew default output
rlabel metal2 s 11150 159200 11206 160000 6 io_out[2]
port 130 nsew default output
rlabel metal2 s 122286 159200 122342 160000 6 io_out[30]
port 131 nsew default output
rlabel metal2 s 126242 159200 126298 160000 6 io_out[31]
port 132 nsew default output
rlabel metal2 s 130198 159200 130254 160000 6 io_out[32]
port 133 nsew default output
rlabel metal2 s 134154 159200 134210 160000 6 io_out[33]
port 134 nsew default output
rlabel metal2 s 138110 159200 138166 160000 6 io_out[34]
port 135 nsew default output
rlabel metal2 s 142066 159200 142122 160000 6 io_out[35]
port 136 nsew default output
rlabel metal2 s 146022 159200 146078 160000 6 io_out[36]
port 137 nsew default output
rlabel metal2 s 150070 159200 150126 160000 6 io_out[37]
port 138 nsew default output
rlabel metal2 s 15198 159200 15254 160000 6 io_out[3]
port 139 nsew default output
rlabel metal2 s 19154 159200 19210 160000 6 io_out[4]
port 140 nsew default output
rlabel metal2 s 23110 159200 23166 160000 6 io_out[5]
port 141 nsew default output
rlabel metal2 s 27066 159200 27122 160000 6 io_out[6]
port 142 nsew default output
rlabel metal2 s 31022 159200 31078 160000 6 io_out[7]
port 143 nsew default output
rlabel metal2 s 34978 159200 35034 160000 6 io_out[8]
port 144 nsew default output
rlabel metal2 s 38934 159200 38990 160000 6 io_out[9]
port 145 nsew default output
rlabel metal2 s 34150 0 34206 800 6 la_data_in[0]
port 146 nsew default input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[100]
port 147 nsew default input
rlabel metal2 s 131486 0 131542 800 6 la_data_in[101]
port 148 nsew default input
rlabel metal2 s 132406 0 132462 800 6 la_data_in[102]
port 149 nsew default input
rlabel metal2 s 133418 0 133474 800 6 la_data_in[103]
port 150 nsew default input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[104]
port 151 nsew default input
rlabel metal2 s 135350 0 135406 800 6 la_data_in[105]
port 152 nsew default input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[106]
port 153 nsew default input
rlabel metal2 s 137282 0 137338 800 6 la_data_in[107]
port 154 nsew default input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[108]
port 155 nsew default input
rlabel metal2 s 139214 0 139270 800 6 la_data_in[109]
port 156 nsew default input
rlabel metal2 s 43718 0 43774 800 6 la_data_in[10]
port 157 nsew default input
rlabel metal2 s 140134 0 140190 800 6 la_data_in[110]
port 158 nsew default input
rlabel metal2 s 141054 0 141110 800 6 la_data_in[111]
port 159 nsew default input
rlabel metal2 s 142066 0 142122 800 6 la_data_in[112]
port 160 nsew default input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[113]
port 161 nsew default input
rlabel metal2 s 143998 0 144054 800 6 la_data_in[114]
port 162 nsew default input
rlabel metal2 s 144918 0 144974 800 6 la_data_in[115]
port 163 nsew default input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[116]
port 164 nsew default input
rlabel metal2 s 146850 0 146906 800 6 la_data_in[117]
port 165 nsew default input
rlabel metal2 s 147862 0 147918 800 6 la_data_in[118]
port 166 nsew default input
rlabel metal2 s 148782 0 148838 800 6 la_data_in[119]
port 167 nsew default input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[11]
port 168 nsew default input
rlabel metal2 s 149794 0 149850 800 6 la_data_in[120]
port 169 nsew default input
rlabel metal2 s 150714 0 150770 800 6 la_data_in[121]
port 170 nsew default input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[122]
port 171 nsew default input
rlabel metal2 s 152646 0 152702 800 6 la_data_in[123]
port 172 nsew default input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[124]
port 173 nsew default input
rlabel metal2 s 154578 0 154634 800 6 la_data_in[125]
port 174 nsew default input
rlabel metal2 s 155590 0 155646 800 6 la_data_in[126]
port 175 nsew default input
rlabel metal2 s 156510 0 156566 800 6 la_data_in[127]
port 176 nsew default input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[12]
port 177 nsew default input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[13]
port 178 nsew default input
rlabel metal2 s 47582 0 47638 800 6 la_data_in[14]
port 179 nsew default input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[15]
port 180 nsew default input
rlabel metal2 s 49514 0 49570 800 6 la_data_in[16]
port 181 nsew default input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[17]
port 182 nsew default input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[18]
port 183 nsew default input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[19]
port 184 nsew default input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[1]
port 185 nsew default input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[20]
port 186 nsew default input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[21]
port 187 nsew default input
rlabel metal2 s 55310 0 55366 800 6 la_data_in[22]
port 188 nsew default input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[23]
port 189 nsew default input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[24]
port 190 nsew default input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[25]
port 191 nsew default input
rlabel metal2 s 59174 0 59230 800 6 la_data_in[26]
port 192 nsew default input
rlabel metal2 s 60094 0 60150 800 6 la_data_in[27]
port 193 nsew default input
rlabel metal2 s 61106 0 61162 800 6 la_data_in[28]
port 194 nsew default input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[29]
port 195 nsew default input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[2]
port 196 nsew default input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[30]
port 197 nsew default input
rlabel metal2 s 63958 0 64014 800 6 la_data_in[31]
port 198 nsew default input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[32]
port 199 nsew default input
rlabel metal2 s 65890 0 65946 800 6 la_data_in[33]
port 200 nsew default input
rlabel metal2 s 66902 0 66958 800 6 la_data_in[34]
port 201 nsew default input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[35]
port 202 nsew default input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[36]
port 203 nsew default input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[37]
port 204 nsew default input
rlabel metal2 s 70766 0 70822 800 6 la_data_in[38]
port 205 nsew default input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[39]
port 206 nsew default input
rlabel metal2 s 37002 0 37058 800 6 la_data_in[3]
port 207 nsew default input
rlabel metal2 s 72698 0 72754 800 6 la_data_in[40]
port 208 nsew default input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[41]
port 209 nsew default input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[42]
port 210 nsew default input
rlabel metal2 s 75550 0 75606 800 6 la_data_in[43]
port 211 nsew default input
rlabel metal2 s 76562 0 76618 800 6 la_data_in[44]
port 212 nsew default input
rlabel metal2 s 77482 0 77538 800 6 la_data_in[45]
port 213 nsew default input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[46]
port 214 nsew default input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[47]
port 215 nsew default input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[48]
port 216 nsew default input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[49]
port 217 nsew default input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[4]
port 218 nsew default input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[50]
port 219 nsew default input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[51]
port 220 nsew default input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[52]
port 221 nsew default input
rlabel metal2 s 85210 0 85266 800 6 la_data_in[53]
port 222 nsew default input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[54]
port 223 nsew default input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[55]
port 224 nsew default input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[56]
port 225 nsew default input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[57]
port 226 nsew default input
rlabel metal2 s 89994 0 90050 800 6 la_data_in[58]
port 227 nsew default input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[59]
port 228 nsew default input
rlabel metal2 s 38934 0 38990 800 6 la_data_in[5]
port 229 nsew default input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[60]
port 230 nsew default input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[61]
port 231 nsew default input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[62]
port 232 nsew default input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[63]
port 233 nsew default input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[64]
port 234 nsew default input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[65]
port 235 nsew default input
rlabel metal2 s 97722 0 97778 800 6 la_data_in[66]
port 236 nsew default input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[67]
port 237 nsew default input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[68]
port 238 nsew default input
rlabel metal2 s 100574 0 100630 800 6 la_data_in[69]
port 239 nsew default input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[6]
port 240 nsew default input
rlabel metal2 s 101586 0 101642 800 6 la_data_in[70]
port 241 nsew default input
rlabel metal2 s 102506 0 102562 800 6 la_data_in[71]
port 242 nsew default input
rlabel metal2 s 103518 0 103574 800 6 la_data_in[72]
port 243 nsew default input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[73]
port 244 nsew default input
rlabel metal2 s 105450 0 105506 800 6 la_data_in[74]
port 245 nsew default input
rlabel metal2 s 106370 0 106426 800 6 la_data_in[75]
port 246 nsew default input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[76]
port 247 nsew default input
rlabel metal2 s 108302 0 108358 800 6 la_data_in[77]
port 248 nsew default input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[78]
port 249 nsew default input
rlabel metal2 s 110234 0 110290 800 6 la_data_in[79]
port 250 nsew default input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[7]
port 251 nsew default input
rlabel metal2 s 111246 0 111302 800 6 la_data_in[80]
port 252 nsew default input
rlabel metal2 s 112166 0 112222 800 6 la_data_in[81]
port 253 nsew default input
rlabel metal2 s 113178 0 113234 800 6 la_data_in[82]
port 254 nsew default input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[83]
port 255 nsew default input
rlabel metal2 s 115110 0 115166 800 6 la_data_in[84]
port 256 nsew default input
rlabel metal2 s 116030 0 116086 800 6 la_data_in[85]
port 257 nsew default input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[86]
port 258 nsew default input
rlabel metal2 s 117962 0 118018 800 6 la_data_in[87]
port 259 nsew default input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[88]
port 260 nsew default input
rlabel metal2 s 119894 0 119950 800 6 la_data_in[89]
port 261 nsew default input
rlabel metal2 s 41786 0 41842 800 6 la_data_in[8]
port 262 nsew default input
rlabel metal2 s 120814 0 120870 800 6 la_data_in[90]
port 263 nsew default input
rlabel metal2 s 121826 0 121882 800 6 la_data_in[91]
port 264 nsew default input
rlabel metal2 s 122746 0 122802 800 6 la_data_in[92]
port 265 nsew default input
rlabel metal2 s 123758 0 123814 800 6 la_data_in[93]
port 266 nsew default input
rlabel metal2 s 124678 0 124734 800 6 la_data_in[94]
port 267 nsew default input
rlabel metal2 s 125690 0 125746 800 6 la_data_in[95]
port 268 nsew default input
rlabel metal2 s 126610 0 126666 800 6 la_data_in[96]
port 269 nsew default input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[97]
port 270 nsew default input
rlabel metal2 s 128542 0 128598 800 6 la_data_in[98]
port 271 nsew default input
rlabel metal2 s 129554 0 129610 800 6 la_data_in[99]
port 272 nsew default input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[9]
port 273 nsew default input
rlabel metal2 s 34426 0 34482 800 6 la_data_out[0]
port 274 nsew default output
rlabel metal2 s 130842 0 130898 800 6 la_data_out[100]
port 275 nsew default output
rlabel metal2 s 131762 0 131818 800 6 la_data_out[101]
port 276 nsew default output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[102]
port 277 nsew default output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[103]
port 278 nsew default output
rlabel metal2 s 134706 0 134762 800 6 la_data_out[104]
port 279 nsew default output
rlabel metal2 s 135626 0 135682 800 6 la_data_out[105]
port 280 nsew default output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[106]
port 281 nsew default output
rlabel metal2 s 137558 0 137614 800 6 la_data_out[107]
port 282 nsew default output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[108]
port 283 nsew default output
rlabel metal2 s 139490 0 139546 800 6 la_data_out[109]
port 284 nsew default output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[10]
port 285 nsew default output
rlabel metal2 s 140410 0 140466 800 6 la_data_out[110]
port 286 nsew default output
rlabel metal2 s 141422 0 141478 800 6 la_data_out[111]
port 287 nsew default output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[112]
port 288 nsew default output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[113]
port 289 nsew default output
rlabel metal2 s 144274 0 144330 800 6 la_data_out[114]
port 290 nsew default output
rlabel metal2 s 145286 0 145342 800 6 la_data_out[115]
port 291 nsew default output
rlabel metal2 s 146206 0 146262 800 6 la_data_out[116]
port 292 nsew default output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[117]
port 293 nsew default output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[118]
port 294 nsew default output
rlabel metal2 s 149150 0 149206 800 6 la_data_out[119]
port 295 nsew default output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[11]
port 296 nsew default output
rlabel metal2 s 150070 0 150126 800 6 la_data_out[120]
port 297 nsew default output
rlabel metal2 s 151082 0 151138 800 6 la_data_out[121]
port 298 nsew default output
rlabel metal2 s 152002 0 152058 800 6 la_data_out[122]
port 299 nsew default output
rlabel metal2 s 153014 0 153070 800 6 la_data_out[123]
port 300 nsew default output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[124]
port 301 nsew default output
rlabel metal2 s 154946 0 155002 800 6 la_data_out[125]
port 302 nsew default output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[126]
port 303 nsew default output
rlabel metal2 s 156878 0 156934 800 6 la_data_out[127]
port 304 nsew default output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[12]
port 305 nsew default output
rlabel metal2 s 46938 0 46994 800 6 la_data_out[13]
port 306 nsew default output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[14]
port 307 nsew default output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[15]
port 308 nsew default output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[16]
port 309 nsew default output
rlabel metal2 s 50802 0 50858 800 6 la_data_out[17]
port 310 nsew default output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[18]
port 311 nsew default output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[19]
port 312 nsew default output
rlabel metal2 s 35438 0 35494 800 6 la_data_out[1]
port 313 nsew default output
rlabel metal2 s 53746 0 53802 800 6 la_data_out[20]
port 314 nsew default output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[21]
port 315 nsew default output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[22]
port 316 nsew default output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[23]
port 317 nsew default output
rlabel metal2 s 57610 0 57666 800 6 la_data_out[24]
port 318 nsew default output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[25]
port 319 nsew default output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[26]
port 320 nsew default output
rlabel metal2 s 60462 0 60518 800 6 la_data_out[27]
port 321 nsew default output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[28]
port 322 nsew default output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[29]
port 323 nsew default output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[2]
port 324 nsew default output
rlabel metal2 s 63314 0 63370 800 6 la_data_out[30]
port 325 nsew default output
rlabel metal2 s 64326 0 64382 800 6 la_data_out[31]
port 326 nsew default output
rlabel metal2 s 65246 0 65302 800 6 la_data_out[32]
port 327 nsew default output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[33]
port 328 nsew default output
rlabel metal2 s 67178 0 67234 800 6 la_data_out[34]
port 329 nsew default output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[35]
port 330 nsew default output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[36]
port 331 nsew default output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[37]
port 332 nsew default output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[38]
port 333 nsew default output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[39]
port 334 nsew default output
rlabel metal2 s 37370 0 37426 800 6 la_data_out[3]
port 335 nsew default output
rlabel metal2 s 72974 0 73030 800 6 la_data_out[40]
port 336 nsew default output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[41]
port 337 nsew default output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[42]
port 338 nsew default output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[43]
port 339 nsew default output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[44]
port 340 nsew default output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[45]
port 341 nsew default output
rlabel metal2 s 78770 0 78826 800 6 la_data_out[46]
port 342 nsew default output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[47]
port 343 nsew default output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[48]
port 344 nsew default output
rlabel metal2 s 81622 0 81678 800 6 la_data_out[49]
port 345 nsew default output
rlabel metal2 s 38290 0 38346 800 6 la_data_out[4]
port 346 nsew default output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[50]
port 347 nsew default output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[51]
port 348 nsew default output
rlabel metal2 s 84566 0 84622 800 6 la_data_out[52]
port 349 nsew default output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[53]
port 350 nsew default output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[54]
port 351 nsew default output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[55]
port 352 nsew default output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[56]
port 353 nsew default output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[57]
port 354 nsew default output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[58]
port 355 nsew default output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[59]
port 356 nsew default output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[5]
port 357 nsew default output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[60]
port 358 nsew default output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[61]
port 359 nsew default output
rlabel metal2 s 94226 0 94282 800 6 la_data_out[62]
port 360 nsew default output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[63]
port 361 nsew default output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[64]
port 362 nsew default output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[65]
port 363 nsew default output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[66]
port 364 nsew default output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[67]
port 365 nsew default output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[68]
port 366 nsew default output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[69]
port 367 nsew default output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[6]
port 368 nsew default output
rlabel metal2 s 101862 0 101918 800 6 la_data_out[70]
port 369 nsew default output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[71]
port 370 nsew default output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[72]
port 371 nsew default output
rlabel metal2 s 104806 0 104862 800 6 la_data_out[73]
port 372 nsew default output
rlabel metal2 s 105726 0 105782 800 6 la_data_out[74]
port 373 nsew default output
rlabel metal2 s 106738 0 106794 800 6 la_data_out[75]
port 374 nsew default output
rlabel metal2 s 107658 0 107714 800 6 la_data_out[76]
port 375 nsew default output
rlabel metal2 s 108670 0 108726 800 6 la_data_out[77]
port 376 nsew default output
rlabel metal2 s 109590 0 109646 800 6 la_data_out[78]
port 377 nsew default output
rlabel metal2 s 110602 0 110658 800 6 la_data_out[79]
port 378 nsew default output
rlabel metal2 s 41142 0 41198 800 6 la_data_out[7]
port 379 nsew default output
rlabel metal2 s 111522 0 111578 800 6 la_data_out[80]
port 380 nsew default output
rlabel metal2 s 112534 0 112590 800 6 la_data_out[81]
port 381 nsew default output
rlabel metal2 s 113454 0 113510 800 6 la_data_out[82]
port 382 nsew default output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[83]
port 383 nsew default output
rlabel metal2 s 115386 0 115442 800 6 la_data_out[84]
port 384 nsew default output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[85]
port 385 nsew default output
rlabel metal2 s 117318 0 117374 800 6 la_data_out[86]
port 386 nsew default output
rlabel metal2 s 118330 0 118386 800 6 la_data_out[87]
port 387 nsew default output
rlabel metal2 s 119250 0 119306 800 6 la_data_out[88]
port 388 nsew default output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[89]
port 389 nsew default output
rlabel metal2 s 42154 0 42210 800 6 la_data_out[8]
port 390 nsew default output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[90]
port 391 nsew default output
rlabel metal2 s 122102 0 122158 800 6 la_data_out[91]
port 392 nsew default output
rlabel metal2 s 123114 0 123170 800 6 la_data_out[92]
port 393 nsew default output
rlabel metal2 s 124034 0 124090 800 6 la_data_out[93]
port 394 nsew default output
rlabel metal2 s 125046 0 125102 800 6 la_data_out[94]
port 395 nsew default output
rlabel metal2 s 125966 0 126022 800 6 la_data_out[95]
port 396 nsew default output
rlabel metal2 s 126978 0 127034 800 6 la_data_out[96]
port 397 nsew default output
rlabel metal2 s 127898 0 127954 800 6 la_data_out[97]
port 398 nsew default output
rlabel metal2 s 128910 0 128966 800 6 la_data_out[98]
port 399 nsew default output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[99]
port 400 nsew default output
rlabel metal2 s 43074 0 43130 800 6 la_data_out[9]
port 401 nsew default output
rlabel metal2 s 34794 0 34850 800 6 la_oen[0]
port 402 nsew default input
rlabel metal2 s 131118 0 131174 800 6 la_oen[100]
port 403 nsew default input
rlabel metal2 s 132130 0 132186 800 6 la_oen[101]
port 404 nsew default input
rlabel metal2 s 133050 0 133106 800 6 la_oen[102]
port 405 nsew default input
rlabel metal2 s 134062 0 134118 800 6 la_oen[103]
port 406 nsew default input
rlabel metal2 s 134982 0 135038 800 6 la_oen[104]
port 407 nsew default input
rlabel metal2 s 135994 0 136050 800 6 la_oen[105]
port 408 nsew default input
rlabel metal2 s 136914 0 136970 800 6 la_oen[106]
port 409 nsew default input
rlabel metal2 s 137926 0 137982 800 6 la_oen[107]
port 410 nsew default input
rlabel metal2 s 138846 0 138902 800 6 la_oen[108]
port 411 nsew default input
rlabel metal2 s 139858 0 139914 800 6 la_oen[109]
port 412 nsew default input
rlabel metal2 s 44362 0 44418 800 6 la_oen[10]
port 413 nsew default input
rlabel metal2 s 140778 0 140834 800 6 la_oen[110]
port 414 nsew default input
rlabel metal2 s 141698 0 141754 800 6 la_oen[111]
port 415 nsew default input
rlabel metal2 s 142710 0 142766 800 6 la_oen[112]
port 416 nsew default input
rlabel metal2 s 143630 0 143686 800 6 la_oen[113]
port 417 nsew default input
rlabel metal2 s 144642 0 144698 800 6 la_oen[114]
port 418 nsew default input
rlabel metal2 s 145562 0 145618 800 6 la_oen[115]
port 419 nsew default input
rlabel metal2 s 146574 0 146630 800 6 la_oen[116]
port 420 nsew default input
rlabel metal2 s 147494 0 147550 800 6 la_oen[117]
port 421 nsew default input
rlabel metal2 s 148506 0 148562 800 6 la_oen[118]
port 422 nsew default input
rlabel metal2 s 149426 0 149482 800 6 la_oen[119]
port 423 nsew default input
rlabel metal2 s 45374 0 45430 800 6 la_oen[11]
port 424 nsew default input
rlabel metal2 s 150438 0 150494 800 6 la_oen[120]
port 425 nsew default input
rlabel metal2 s 151358 0 151414 800 6 la_oen[121]
port 426 nsew default input
rlabel metal2 s 152370 0 152426 800 6 la_oen[122]
port 427 nsew default input
rlabel metal2 s 153290 0 153346 800 6 la_oen[123]
port 428 nsew default input
rlabel metal2 s 154302 0 154358 800 6 la_oen[124]
port 429 nsew default input
rlabel metal2 s 155222 0 155278 800 6 la_oen[125]
port 430 nsew default input
rlabel metal2 s 156234 0 156290 800 6 la_oen[126]
port 431 nsew default input
rlabel metal2 s 157154 0 157210 800 6 la_oen[127]
port 432 nsew default input
rlabel metal2 s 46294 0 46350 800 6 la_oen[12]
port 433 nsew default input
rlabel metal2 s 47306 0 47362 800 6 la_oen[13]
port 434 nsew default input
rlabel metal2 s 48226 0 48282 800 6 la_oen[14]
port 435 nsew default input
rlabel metal2 s 49238 0 49294 800 6 la_oen[15]
port 436 nsew default input
rlabel metal2 s 50158 0 50214 800 6 la_oen[16]
port 437 nsew default input
rlabel metal2 s 51170 0 51226 800 6 la_oen[17]
port 438 nsew default input
rlabel metal2 s 52090 0 52146 800 6 la_oen[18]
port 439 nsew default input
rlabel metal2 s 53102 0 53158 800 6 la_oen[19]
port 440 nsew default input
rlabel metal2 s 35714 0 35770 800 6 la_oen[1]
port 441 nsew default input
rlabel metal2 s 54022 0 54078 800 6 la_oen[20]
port 442 nsew default input
rlabel metal2 s 55034 0 55090 800 6 la_oen[21]
port 443 nsew default input
rlabel metal2 s 55954 0 56010 800 6 la_oen[22]
port 444 nsew default input
rlabel metal2 s 56966 0 57022 800 6 la_oen[23]
port 445 nsew default input
rlabel metal2 s 57886 0 57942 800 6 la_oen[24]
port 446 nsew default input
rlabel metal2 s 58898 0 58954 800 6 la_oen[25]
port 447 nsew default input
rlabel metal2 s 59818 0 59874 800 6 la_oen[26]
port 448 nsew default input
rlabel metal2 s 60738 0 60794 800 6 la_oen[27]
port 449 nsew default input
rlabel metal2 s 61750 0 61806 800 6 la_oen[28]
port 450 nsew default input
rlabel metal2 s 62670 0 62726 800 6 la_oen[29]
port 451 nsew default input
rlabel metal2 s 36726 0 36782 800 6 la_oen[2]
port 452 nsew default input
rlabel metal2 s 63682 0 63738 800 6 la_oen[30]
port 453 nsew default input
rlabel metal2 s 64602 0 64658 800 6 la_oen[31]
port 454 nsew default input
rlabel metal2 s 65614 0 65670 800 6 la_oen[32]
port 455 nsew default input
rlabel metal2 s 66534 0 66590 800 6 la_oen[33]
port 456 nsew default input
rlabel metal2 s 67546 0 67602 800 6 la_oen[34]
port 457 nsew default input
rlabel metal2 s 68466 0 68522 800 6 la_oen[35]
port 458 nsew default input
rlabel metal2 s 69478 0 69534 800 6 la_oen[36]
port 459 nsew default input
rlabel metal2 s 70398 0 70454 800 6 la_oen[37]
port 460 nsew default input
rlabel metal2 s 71410 0 71466 800 6 la_oen[38]
port 461 nsew default input
rlabel metal2 s 72330 0 72386 800 6 la_oen[39]
port 462 nsew default input
rlabel metal2 s 37646 0 37702 800 6 la_oen[3]
port 463 nsew default input
rlabel metal2 s 73342 0 73398 800 6 la_oen[40]
port 464 nsew default input
rlabel metal2 s 74262 0 74318 800 6 la_oen[41]
port 465 nsew default input
rlabel metal2 s 75274 0 75330 800 6 la_oen[42]
port 466 nsew default input
rlabel metal2 s 76194 0 76250 800 6 la_oen[43]
port 467 nsew default input
rlabel metal2 s 77206 0 77262 800 6 la_oen[44]
port 468 nsew default input
rlabel metal2 s 78126 0 78182 800 6 la_oen[45]
port 469 nsew default input
rlabel metal2 s 79138 0 79194 800 6 la_oen[46]
port 470 nsew default input
rlabel metal2 s 80058 0 80114 800 6 la_oen[47]
port 471 nsew default input
rlabel metal2 s 80978 0 81034 800 6 la_oen[48]
port 472 nsew default input
rlabel metal2 s 81990 0 82046 800 6 la_oen[49]
port 473 nsew default input
rlabel metal2 s 38658 0 38714 800 6 la_oen[4]
port 474 nsew default input
rlabel metal2 s 82910 0 82966 800 6 la_oen[50]
port 475 nsew default input
rlabel metal2 s 83922 0 83978 800 6 la_oen[51]
port 476 nsew default input
rlabel metal2 s 84842 0 84898 800 6 la_oen[52]
port 477 nsew default input
rlabel metal2 s 85854 0 85910 800 6 la_oen[53]
port 478 nsew default input
rlabel metal2 s 86774 0 86830 800 6 la_oen[54]
port 479 nsew default input
rlabel metal2 s 87786 0 87842 800 6 la_oen[55]
port 480 nsew default input
rlabel metal2 s 88706 0 88762 800 6 la_oen[56]
port 481 nsew default input
rlabel metal2 s 89718 0 89774 800 6 la_oen[57]
port 482 nsew default input
rlabel metal2 s 90638 0 90694 800 6 la_oen[58]
port 483 nsew default input
rlabel metal2 s 91650 0 91706 800 6 la_oen[59]
port 484 nsew default input
rlabel metal2 s 39578 0 39634 800 6 la_oen[5]
port 485 nsew default input
rlabel metal2 s 92570 0 92626 800 6 la_oen[60]
port 486 nsew default input
rlabel metal2 s 93582 0 93638 800 6 la_oen[61]
port 487 nsew default input
rlabel metal2 s 94502 0 94558 800 6 la_oen[62]
port 488 nsew default input
rlabel metal2 s 95514 0 95570 800 6 la_oen[63]
port 489 nsew default input
rlabel metal2 s 96434 0 96490 800 6 la_oen[64]
port 490 nsew default input
rlabel metal2 s 97446 0 97502 800 6 la_oen[65]
port 491 nsew default input
rlabel metal2 s 98366 0 98422 800 6 la_oen[66]
port 492 nsew default input
rlabel metal2 s 99378 0 99434 800 6 la_oen[67]
port 493 nsew default input
rlabel metal2 s 100298 0 100354 800 6 la_oen[68]
port 494 nsew default input
rlabel metal2 s 101218 0 101274 800 6 la_oen[69]
port 495 nsew default input
rlabel metal2 s 40498 0 40554 800 6 la_oen[6]
port 496 nsew default input
rlabel metal2 s 102230 0 102286 800 6 la_oen[70]
port 497 nsew default input
rlabel metal2 s 103150 0 103206 800 6 la_oen[71]
port 498 nsew default input
rlabel metal2 s 104162 0 104218 800 6 la_oen[72]
port 499 nsew default input
rlabel metal2 s 105082 0 105138 800 6 la_oen[73]
port 500 nsew default input
rlabel metal2 s 106094 0 106150 800 6 la_oen[74]
port 501 nsew default input
rlabel metal2 s 107014 0 107070 800 6 la_oen[75]
port 502 nsew default input
rlabel metal2 s 108026 0 108082 800 6 la_oen[76]
port 503 nsew default input
rlabel metal2 s 108946 0 109002 800 6 la_oen[77]
port 504 nsew default input
rlabel metal2 s 109958 0 110014 800 6 la_oen[78]
port 505 nsew default input
rlabel metal2 s 110878 0 110934 800 6 la_oen[79]
port 506 nsew default input
rlabel metal2 s 41510 0 41566 800 6 la_oen[7]
port 507 nsew default input
rlabel metal2 s 111890 0 111946 800 6 la_oen[80]
port 508 nsew default input
rlabel metal2 s 112810 0 112866 800 6 la_oen[81]
port 509 nsew default input
rlabel metal2 s 113822 0 113878 800 6 la_oen[82]
port 510 nsew default input
rlabel metal2 s 114742 0 114798 800 6 la_oen[83]
port 511 nsew default input
rlabel metal2 s 115754 0 115810 800 6 la_oen[84]
port 512 nsew default input
rlabel metal2 s 116674 0 116730 800 6 la_oen[85]
port 513 nsew default input
rlabel metal2 s 117686 0 117742 800 6 la_oen[86]
port 514 nsew default input
rlabel metal2 s 118606 0 118662 800 6 la_oen[87]
port 515 nsew default input
rlabel metal2 s 119618 0 119674 800 6 la_oen[88]
port 516 nsew default input
rlabel metal2 s 120538 0 120594 800 6 la_oen[89]
port 517 nsew default input
rlabel metal2 s 42430 0 42486 800 6 la_oen[8]
port 518 nsew default input
rlabel metal2 s 121458 0 121514 800 6 la_oen[90]
port 519 nsew default input
rlabel metal2 s 122470 0 122526 800 6 la_oen[91]
port 520 nsew default input
rlabel metal2 s 123390 0 123446 800 6 la_oen[92]
port 521 nsew default input
rlabel metal2 s 124402 0 124458 800 6 la_oen[93]
port 522 nsew default input
rlabel metal2 s 125322 0 125378 800 6 la_oen[94]
port 523 nsew default input
rlabel metal2 s 126334 0 126390 800 6 la_oen[95]
port 524 nsew default input
rlabel metal2 s 127254 0 127310 800 6 la_oen[96]
port 525 nsew default input
rlabel metal2 s 128266 0 128322 800 6 la_oen[97]
port 526 nsew default input
rlabel metal2 s 129186 0 129242 800 6 la_oen[98]
port 527 nsew default input
rlabel metal2 s 130198 0 130254 800 6 la_oen[99]
port 528 nsew default input
rlabel metal2 s 43442 0 43498 800 6 la_oen[9]
port 529 nsew default input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 530 nsew default input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 531 nsew default input
rlabel metal2 s 662 0 718 800 6 wbs_ack_o
port 532 nsew default output
rlabel metal2 s 1950 0 2006 800 6 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 13910 0 13966 800 6 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 18694 0 18750 800 6 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 20626 0 20682 800 6 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 3238 0 3294 800 6 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 23478 0 23534 800 6 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 25410 0 25466 800 6 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 28354 0 28410 800 6 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 30286 0 30342 800 6 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 32218 0 32274 800 6 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 33138 0 33194 800 6 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 7102 0 7158 800 6 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 1030 0 1086 800 6 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_o[0]
port 598 nsew default output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[10]
port 599 nsew default output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[11]
port 600 nsew default output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[12]
port 601 nsew default output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[13]
port 602 nsew default output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[14]
port 603 nsew default output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[15]
port 604 nsew default output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[16]
port 605 nsew default output
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_o[17]
port 606 nsew default output
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_o[18]
port 607 nsew default output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[19]
port 608 nsew default output
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[1]
port 609 nsew default output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[20]
port 610 nsew default output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[21]
port 611 nsew default output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[22]
port 612 nsew default output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[23]
port 613 nsew default output
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_o[24]
port 614 nsew default output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[25]
port 615 nsew default output
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_o[26]
port 616 nsew default output
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_o[27]
port 617 nsew default output
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_o[28]
port 618 nsew default output
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_o[29]
port 619 nsew default output
rlabel metal2 s 5170 0 5226 800 6 wbs_dat_o[2]
port 620 nsew default output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[30]
port 621 nsew default output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[31]
port 622 nsew default output
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_o[3]
port 623 nsew default output
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_o[4]
port 624 nsew default output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[5]
port 625 nsew default output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[6]
port 626 nsew default output
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_o[7]
port 627 nsew default output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[8]
port 628 nsew default output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[9]
port 629 nsew default output
rlabel metal2 s 2962 0 3018 800 6 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 4250 0 4306 800 6 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 5538 0 5594 800 6 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 6826 0 6882 800 6 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 1306 0 1362 800 6 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 1674 0 1730 800 6 wbs_we_i
port 635 nsew default input
rlabel metal4 s 4208 2128 4528 157808 6 VPWR
port 636 nsew power input
rlabel metal4 s 19568 2128 19888 157808 6 VGND
port 637 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 160000 160000
string LEFview TRUE
<< end >>
