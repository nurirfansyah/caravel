magic
tech sky130A
magscale 1 2
timestamp 1608026852
<< obsli1 >>
rect 1104 2159 158884 157777
<< obsm1 >>
rect 750 1640 158884 157808
<< metal2 >>
rect 662 159200 718 160000
rect 1950 159200 2006 160000
rect 3238 159200 3294 160000
rect 4526 159200 4582 160000
rect 5814 159200 5870 160000
rect 7102 159200 7158 160000
rect 8390 159200 8446 160000
rect 9678 159200 9734 160000
rect 10966 159200 11022 160000
rect 12254 159200 12310 160000
rect 13542 159200 13598 160000
rect 14830 159200 14886 160000
rect 16118 159200 16174 160000
rect 17406 159200 17462 160000
rect 18694 159200 18750 160000
rect 19982 159200 20038 160000
rect 21270 159200 21326 160000
rect 22558 159200 22614 160000
rect 23846 159200 23902 160000
rect 25134 159200 25190 160000
rect 26422 159200 26478 160000
rect 27710 159200 27766 160000
rect 28998 159200 29054 160000
rect 30286 159200 30342 160000
rect 31574 159200 31630 160000
rect 32862 159200 32918 160000
rect 34150 159200 34206 160000
rect 35438 159200 35494 160000
rect 36726 159200 36782 160000
rect 38014 159200 38070 160000
rect 39302 159200 39358 160000
rect 40590 159200 40646 160000
rect 41878 159200 41934 160000
rect 43166 159200 43222 160000
rect 44454 159200 44510 160000
rect 45742 159200 45798 160000
rect 47030 159200 47086 160000
rect 48318 159200 48374 160000
rect 49606 159200 49662 160000
rect 50894 159200 50950 160000
rect 52182 159200 52238 160000
rect 53470 159200 53526 160000
rect 54850 159200 54906 160000
rect 56138 159200 56194 160000
rect 57426 159200 57482 160000
rect 58714 159200 58770 160000
rect 60002 159200 60058 160000
rect 61290 159200 61346 160000
rect 62578 159200 62634 160000
rect 63866 159200 63922 160000
rect 65154 159200 65210 160000
rect 66442 159200 66498 160000
rect 67730 159200 67786 160000
rect 69018 159200 69074 160000
rect 70306 159200 70362 160000
rect 71594 159200 71650 160000
rect 72882 159200 72938 160000
rect 74170 159200 74226 160000
rect 75458 159200 75514 160000
rect 76746 159200 76802 160000
rect 78034 159200 78090 160000
rect 79322 159200 79378 160000
rect 80610 159200 80666 160000
rect 81898 159200 81954 160000
rect 83186 159200 83242 160000
rect 84474 159200 84530 160000
rect 85762 159200 85818 160000
rect 87050 159200 87106 160000
rect 88338 159200 88394 160000
rect 89626 159200 89682 160000
rect 90914 159200 90970 160000
rect 92202 159200 92258 160000
rect 93490 159200 93546 160000
rect 94778 159200 94834 160000
rect 96066 159200 96122 160000
rect 97354 159200 97410 160000
rect 98642 159200 98698 160000
rect 99930 159200 99986 160000
rect 101218 159200 101274 160000
rect 102506 159200 102562 160000
rect 103794 159200 103850 160000
rect 105082 159200 105138 160000
rect 106370 159200 106426 160000
rect 107750 159200 107806 160000
rect 109038 159200 109094 160000
rect 110326 159200 110382 160000
rect 111614 159200 111670 160000
rect 112902 159200 112958 160000
rect 114190 159200 114246 160000
rect 115478 159200 115534 160000
rect 116766 159200 116822 160000
rect 118054 159200 118110 160000
rect 119342 159200 119398 160000
rect 120630 159200 120686 160000
rect 121918 159200 121974 160000
rect 123206 159200 123262 160000
rect 124494 159200 124550 160000
rect 125782 159200 125838 160000
rect 127070 159200 127126 160000
rect 128358 159200 128414 160000
rect 129646 159200 129702 160000
rect 130934 159200 130990 160000
rect 132222 159200 132278 160000
rect 133510 159200 133566 160000
rect 134798 159200 134854 160000
rect 136086 159200 136142 160000
rect 137374 159200 137430 160000
rect 138662 159200 138718 160000
rect 139950 159200 140006 160000
rect 141238 159200 141294 160000
rect 142526 159200 142582 160000
rect 143814 159200 143870 160000
rect 145102 159200 145158 160000
rect 146390 159200 146446 160000
rect 147678 159200 147734 160000
rect 148966 159200 149022 160000
rect 150254 159200 150310 160000
rect 151542 159200 151598 160000
rect 152830 159200 152886 160000
rect 154118 159200 154174 160000
rect 155406 159200 155462 160000
rect 156694 159200 156750 160000
rect 157982 159200 158038 160000
rect 159270 159200 159326 160000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26514 0 26570 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31390 0 31446 800
rect 31666 0 31722 800
rect 32034 0 32090 800
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35254 0 35310 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36174 0 36230 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39118 0 39174 800
rect 39394 0 39450 800
rect 39762 0 39818 800
rect 40038 0 40094 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41326 0 41382 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42982 0 43038 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43902 0 43958 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44914 0 44970 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46846 0 46902 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 50986 0 51042 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54942 0 54998 800
rect 55218 0 55274 800
rect 55586 0 55642 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57150 0 57206 800
rect 57518 0 57574 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58806 0 58862 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59726 0 59782 800
rect 60094 0 60150 800
rect 60370 0 60426 800
rect 60738 0 60794 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61658 0 61714 800
rect 62026 0 62082 800
rect 62302 0 62358 800
rect 62670 0 62726 800
rect 62946 0 63002 800
rect 63314 0 63370 800
rect 63590 0 63646 800
rect 63958 0 64014 800
rect 64234 0 64290 800
rect 64602 0 64658 800
rect 64878 0 64934 800
rect 65246 0 65302 800
rect 65522 0 65578 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67454 0 67510 800
rect 67822 0 67878 800
rect 68098 0 68154 800
rect 68466 0 68522 800
rect 68742 0 68798 800
rect 69110 0 69166 800
rect 69386 0 69442 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70398 0 70454 800
rect 70674 0 70730 800
rect 71042 0 71098 800
rect 71318 0 71374 800
rect 71686 0 71742 800
rect 71962 0 72018 800
rect 72330 0 72386 800
rect 72606 0 72662 800
rect 72974 0 73030 800
rect 73250 0 73306 800
rect 73618 0 73674 800
rect 73894 0 73950 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75182 0 75238 800
rect 75550 0 75606 800
rect 75826 0 75882 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76838 0 76894 800
rect 77114 0 77170 800
rect 77482 0 77538 800
rect 77758 0 77814 800
rect 78126 0 78182 800
rect 78402 0 78458 800
rect 78770 0 78826 800
rect 79046 0 79102 800
rect 79414 0 79470 800
rect 79690 0 79746 800
rect 80058 0 80114 800
rect 80426 0 80482 800
rect 80702 0 80758 800
rect 81070 0 81126 800
rect 81346 0 81402 800
rect 81714 0 81770 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82634 0 82690 800
rect 83002 0 83058 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 83922 0 83978 800
rect 84290 0 84346 800
rect 84566 0 84622 800
rect 84934 0 84990 800
rect 85210 0 85266 800
rect 85578 0 85634 800
rect 85854 0 85910 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86866 0 86922 800
rect 87142 0 87198 800
rect 87510 0 87566 800
rect 87786 0 87842 800
rect 88154 0 88210 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89074 0 89130 800
rect 89442 0 89498 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90730 0 90786 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91650 0 91706 800
rect 92018 0 92074 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 92938 0 92994 800
rect 93306 0 93362 800
rect 93582 0 93638 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94594 0 94650 800
rect 94870 0 94926 800
rect 95238 0 95294 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96158 0 96214 800
rect 96526 0 96582 800
rect 96802 0 96858 800
rect 97170 0 97226 800
rect 97446 0 97502 800
rect 97814 0 97870 800
rect 98090 0 98146 800
rect 98458 0 98514 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99378 0 99434 800
rect 99746 0 99802 800
rect 100022 0 100078 800
rect 100390 0 100446 800
rect 100666 0 100722 800
rect 101034 0 101090 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 101954 0 102010 800
rect 102322 0 102378 800
rect 102598 0 102654 800
rect 102966 0 103022 800
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 103886 0 103942 800
rect 104254 0 104310 800
rect 104530 0 104586 800
rect 104898 0 104954 800
rect 105174 0 105230 800
rect 105542 0 105598 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109406 0 109462 800
rect 109774 0 109830 800
rect 110050 0 110106 800
rect 110418 0 110474 800
rect 110694 0 110750 800
rect 111062 0 111118 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112626 0 112682 800
rect 112994 0 113050 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 113914 0 113970 800
rect 114282 0 114338 800
rect 114558 0 114614 800
rect 114926 0 114982 800
rect 115202 0 115258 800
rect 115570 0 115626 800
rect 115846 0 115902 800
rect 116214 0 116270 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117134 0 117190 800
rect 117502 0 117558 800
rect 117778 0 117834 800
rect 118146 0 118202 800
rect 118422 0 118478 800
rect 118790 0 118846 800
rect 119066 0 119122 800
rect 119434 0 119490 800
rect 119710 0 119766 800
rect 120078 0 120134 800
rect 120354 0 120410 800
rect 120722 0 120778 800
rect 120998 0 121054 800
rect 121366 0 121422 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122286 0 122342 800
rect 122654 0 122710 800
rect 122930 0 122986 800
rect 123298 0 123354 800
rect 123574 0 123630 800
rect 123942 0 123998 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124862 0 124918 800
rect 125230 0 125286 800
rect 125506 0 125562 800
rect 125874 0 125930 800
rect 126150 0 126206 800
rect 126518 0 126574 800
rect 126794 0 126850 800
rect 127162 0 127218 800
rect 127438 0 127494 800
rect 127806 0 127862 800
rect 128082 0 128138 800
rect 128450 0 128506 800
rect 128726 0 128782 800
rect 129094 0 129150 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130014 0 130070 800
rect 130382 0 130438 800
rect 130658 0 130714 800
rect 131026 0 131082 800
rect 131302 0 131358 800
rect 131670 0 131726 800
rect 131946 0 132002 800
rect 132314 0 132370 800
rect 132590 0 132646 800
rect 132958 0 133014 800
rect 133234 0 133290 800
rect 133602 0 133658 800
rect 133970 0 134026 800
rect 134246 0 134302 800
rect 134614 0 134670 800
rect 134890 0 134946 800
rect 135258 0 135314 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136178 0 136234 800
rect 136546 0 136602 800
rect 136822 0 136878 800
rect 137190 0 137246 800
rect 137466 0 137522 800
rect 137834 0 137890 800
rect 138110 0 138166 800
rect 138478 0 138534 800
rect 138754 0 138810 800
rect 139122 0 139178 800
rect 139398 0 139454 800
rect 139766 0 139822 800
rect 140042 0 140098 800
rect 140410 0 140466 800
rect 140686 0 140742 800
rect 141054 0 141110 800
rect 141330 0 141386 800
rect 141698 0 141754 800
rect 141974 0 142030 800
rect 142342 0 142398 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143262 0 143318 800
rect 143630 0 143686 800
rect 143906 0 143962 800
rect 144274 0 144330 800
rect 144550 0 144606 800
rect 144918 0 144974 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145838 0 145894 800
rect 146206 0 146262 800
rect 146482 0 146538 800
rect 146850 0 146906 800
rect 147126 0 147182 800
rect 147494 0 147550 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148414 0 148470 800
rect 148782 0 148838 800
rect 149058 0 149114 800
rect 149426 0 149482 800
rect 149702 0 149758 800
rect 150070 0 150126 800
rect 150346 0 150402 800
rect 150714 0 150770 800
rect 150990 0 151046 800
rect 151358 0 151414 800
rect 151634 0 151690 800
rect 152002 0 152058 800
rect 152278 0 152334 800
rect 152646 0 152702 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153566 0 153622 800
rect 153934 0 153990 800
rect 154210 0 154266 800
rect 154578 0 154634 800
rect 154854 0 154910 800
rect 155222 0 155278 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156142 0 156198 800
rect 156510 0 156566 800
rect 156786 0 156842 800
rect 157154 0 157210 800
rect 157430 0 157486 800
rect 157798 0 157854 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158718 0 158774 800
rect 159086 0 159142 800
rect 159362 0 159418 800
rect 159730 0 159786 800
<< obsm2 >>
rect 110 159144 606 159202
rect 774 159144 1894 159202
rect 2062 159144 3182 159202
rect 3350 159144 4470 159202
rect 4638 159144 5758 159202
rect 5926 159144 7046 159202
rect 7214 159144 8334 159202
rect 8502 159144 9622 159202
rect 9790 159144 10910 159202
rect 11078 159144 12198 159202
rect 12366 159144 13486 159202
rect 13654 159144 14774 159202
rect 14942 159144 16062 159202
rect 16230 159144 17350 159202
rect 17518 159144 18638 159202
rect 18806 159144 19926 159202
rect 20094 159144 21214 159202
rect 21382 159144 22502 159202
rect 22670 159144 23790 159202
rect 23958 159144 25078 159202
rect 25246 159144 26366 159202
rect 26534 159144 27654 159202
rect 27822 159144 28942 159202
rect 29110 159144 30230 159202
rect 30398 159144 31518 159202
rect 31686 159144 32806 159202
rect 32974 159144 34094 159202
rect 34262 159144 35382 159202
rect 35550 159144 36670 159202
rect 36838 159144 37958 159202
rect 38126 159144 39246 159202
rect 39414 159144 40534 159202
rect 40702 159144 41822 159202
rect 41990 159144 43110 159202
rect 43278 159144 44398 159202
rect 44566 159144 45686 159202
rect 45854 159144 46974 159202
rect 47142 159144 48262 159202
rect 48430 159144 49550 159202
rect 49718 159144 50838 159202
rect 51006 159144 52126 159202
rect 52294 159144 53414 159202
rect 53582 159144 54794 159202
rect 54962 159144 56082 159202
rect 56250 159144 57370 159202
rect 57538 159144 58658 159202
rect 58826 159144 59946 159202
rect 60114 159144 61234 159202
rect 61402 159144 62522 159202
rect 62690 159144 63810 159202
rect 63978 159144 65098 159202
rect 65266 159144 66386 159202
rect 66554 159144 67674 159202
rect 67842 159144 68962 159202
rect 69130 159144 70250 159202
rect 70418 159144 71538 159202
rect 71706 159144 72826 159202
rect 72994 159144 74114 159202
rect 74282 159144 75402 159202
rect 75570 159144 76690 159202
rect 76858 159144 77978 159202
rect 78146 159144 79266 159202
rect 79434 159144 80554 159202
rect 80722 159144 81842 159202
rect 82010 159144 83130 159202
rect 83298 159144 84418 159202
rect 84586 159144 85706 159202
rect 85874 159144 86994 159202
rect 87162 159144 88282 159202
rect 88450 159144 89570 159202
rect 89738 159144 90858 159202
rect 91026 159144 92146 159202
rect 92314 159144 93434 159202
rect 93602 159144 94722 159202
rect 94890 159144 96010 159202
rect 96178 159144 97298 159202
rect 97466 159144 98586 159202
rect 98754 159144 99874 159202
rect 100042 159144 101162 159202
rect 101330 159144 102450 159202
rect 102618 159144 103738 159202
rect 103906 159144 105026 159202
rect 105194 159144 106314 159202
rect 106482 159144 107694 159202
rect 107862 159144 108982 159202
rect 109150 159144 110270 159202
rect 110438 159144 111558 159202
rect 111726 159144 112846 159202
rect 113014 159144 114134 159202
rect 114302 159144 115422 159202
rect 115590 159144 116710 159202
rect 116878 159144 117998 159202
rect 118166 159144 119286 159202
rect 119454 159144 120574 159202
rect 120742 159144 121862 159202
rect 122030 159144 123150 159202
rect 123318 159144 124438 159202
rect 124606 159144 125726 159202
rect 125894 159144 127014 159202
rect 127182 159144 128302 159202
rect 128470 159144 129590 159202
rect 129758 159144 130878 159202
rect 131046 159144 132166 159202
rect 132334 159144 133454 159202
rect 133622 159144 134742 159202
rect 134910 159144 136030 159202
rect 136198 159144 137318 159202
rect 137486 159144 138606 159202
rect 138774 159144 139894 159202
rect 140062 159144 141182 159202
rect 141350 159144 142470 159202
rect 142638 159144 143758 159202
rect 143926 159144 145046 159202
rect 145214 159144 146334 159202
rect 146502 159144 147622 159202
rect 147790 159144 148910 159202
rect 149078 159144 150198 159202
rect 150366 159144 151486 159202
rect 151654 159144 152774 159202
rect 152942 159144 154062 159202
rect 154230 159144 155350 159202
rect 155518 159144 156638 159202
rect 156806 159144 157926 159202
rect 158094 159144 158116 159202
rect 110 856 158116 159144
rect 222 800 330 856
rect 498 800 698 856
rect 866 800 974 856
rect 1142 800 1342 856
rect 1510 800 1618 856
rect 1786 800 1986 856
rect 2154 800 2262 856
rect 2430 800 2630 856
rect 2798 800 2906 856
rect 3074 800 3274 856
rect 3442 800 3550 856
rect 3718 800 3918 856
rect 4086 800 4194 856
rect 4362 800 4562 856
rect 4730 800 4838 856
rect 5006 800 5206 856
rect 5374 800 5482 856
rect 5650 800 5850 856
rect 6018 800 6126 856
rect 6294 800 6494 856
rect 6662 800 6770 856
rect 6938 800 7138 856
rect 7306 800 7414 856
rect 7582 800 7782 856
rect 7950 800 8058 856
rect 8226 800 8426 856
rect 8594 800 8702 856
rect 8870 800 9070 856
rect 9238 800 9346 856
rect 9514 800 9714 856
rect 9882 800 9990 856
rect 10158 800 10358 856
rect 10526 800 10634 856
rect 10802 800 11002 856
rect 11170 800 11278 856
rect 11446 800 11646 856
rect 11814 800 11922 856
rect 12090 800 12290 856
rect 12458 800 12566 856
rect 12734 800 12934 856
rect 13102 800 13210 856
rect 13378 800 13578 856
rect 13746 800 13854 856
rect 14022 800 14222 856
rect 14390 800 14498 856
rect 14666 800 14866 856
rect 15034 800 15142 856
rect 15310 800 15510 856
rect 15678 800 15786 856
rect 15954 800 16154 856
rect 16322 800 16430 856
rect 16598 800 16798 856
rect 16966 800 17074 856
rect 17242 800 17442 856
rect 17610 800 17718 856
rect 17886 800 18086 856
rect 18254 800 18362 856
rect 18530 800 18730 856
rect 18898 800 19006 856
rect 19174 800 19374 856
rect 19542 800 19650 856
rect 19818 800 20018 856
rect 20186 800 20294 856
rect 20462 800 20662 856
rect 20830 800 20938 856
rect 21106 800 21306 856
rect 21474 800 21582 856
rect 21750 800 21950 856
rect 22118 800 22226 856
rect 22394 800 22594 856
rect 22762 800 22870 856
rect 23038 800 23238 856
rect 23406 800 23514 856
rect 23682 800 23882 856
rect 24050 800 24158 856
rect 24326 800 24526 856
rect 24694 800 24802 856
rect 24970 800 25170 856
rect 25338 800 25446 856
rect 25614 800 25814 856
rect 25982 800 26090 856
rect 26258 800 26458 856
rect 26626 800 26826 856
rect 26994 800 27102 856
rect 27270 800 27470 856
rect 27638 800 27746 856
rect 27914 800 28114 856
rect 28282 800 28390 856
rect 28558 800 28758 856
rect 28926 800 29034 856
rect 29202 800 29402 856
rect 29570 800 29678 856
rect 29846 800 30046 856
rect 30214 800 30322 856
rect 30490 800 30690 856
rect 30858 800 30966 856
rect 31134 800 31334 856
rect 31502 800 31610 856
rect 31778 800 31978 856
rect 32146 800 32254 856
rect 32422 800 32622 856
rect 32790 800 32898 856
rect 33066 800 33266 856
rect 33434 800 33542 856
rect 33710 800 33910 856
rect 34078 800 34186 856
rect 34354 800 34554 856
rect 34722 800 34830 856
rect 34998 800 35198 856
rect 35366 800 35474 856
rect 35642 800 35842 856
rect 36010 800 36118 856
rect 36286 800 36486 856
rect 36654 800 36762 856
rect 36930 800 37130 856
rect 37298 800 37406 856
rect 37574 800 37774 856
rect 37942 800 38050 856
rect 38218 800 38418 856
rect 38586 800 38694 856
rect 38862 800 39062 856
rect 39230 800 39338 856
rect 39506 800 39706 856
rect 39874 800 39982 856
rect 40150 800 40350 856
rect 40518 800 40626 856
rect 40794 800 40994 856
rect 41162 800 41270 856
rect 41438 800 41638 856
rect 41806 800 41914 856
rect 42082 800 42282 856
rect 42450 800 42558 856
rect 42726 800 42926 856
rect 43094 800 43202 856
rect 43370 800 43570 856
rect 43738 800 43846 856
rect 44014 800 44214 856
rect 44382 800 44490 856
rect 44658 800 44858 856
rect 45026 800 45134 856
rect 45302 800 45502 856
rect 45670 800 45778 856
rect 45946 800 46146 856
rect 46314 800 46422 856
rect 46590 800 46790 856
rect 46958 800 47066 856
rect 47234 800 47434 856
rect 47602 800 47710 856
rect 47878 800 48078 856
rect 48246 800 48354 856
rect 48522 800 48722 856
rect 48890 800 48998 856
rect 49166 800 49366 856
rect 49534 800 49642 856
rect 49810 800 50010 856
rect 50178 800 50286 856
rect 50454 800 50654 856
rect 50822 800 50930 856
rect 51098 800 51298 856
rect 51466 800 51574 856
rect 51742 800 51942 856
rect 52110 800 52218 856
rect 52386 800 52586 856
rect 52754 800 52862 856
rect 53030 800 53230 856
rect 53398 800 53598 856
rect 53766 800 53874 856
rect 54042 800 54242 856
rect 54410 800 54518 856
rect 54686 800 54886 856
rect 55054 800 55162 856
rect 55330 800 55530 856
rect 55698 800 55806 856
rect 55974 800 56174 856
rect 56342 800 56450 856
rect 56618 800 56818 856
rect 56986 800 57094 856
rect 57262 800 57462 856
rect 57630 800 57738 856
rect 57906 800 58106 856
rect 58274 800 58382 856
rect 58550 800 58750 856
rect 58918 800 59026 856
rect 59194 800 59394 856
rect 59562 800 59670 856
rect 59838 800 60038 856
rect 60206 800 60314 856
rect 60482 800 60682 856
rect 60850 800 60958 856
rect 61126 800 61326 856
rect 61494 800 61602 856
rect 61770 800 61970 856
rect 62138 800 62246 856
rect 62414 800 62614 856
rect 62782 800 62890 856
rect 63058 800 63258 856
rect 63426 800 63534 856
rect 63702 800 63902 856
rect 64070 800 64178 856
rect 64346 800 64546 856
rect 64714 800 64822 856
rect 64990 800 65190 856
rect 65358 800 65466 856
rect 65634 800 65834 856
rect 66002 800 66110 856
rect 66278 800 66478 856
rect 66646 800 66754 856
rect 66922 800 67122 856
rect 67290 800 67398 856
rect 67566 800 67766 856
rect 67934 800 68042 856
rect 68210 800 68410 856
rect 68578 800 68686 856
rect 68854 800 69054 856
rect 69222 800 69330 856
rect 69498 800 69698 856
rect 69866 800 69974 856
rect 70142 800 70342 856
rect 70510 800 70618 856
rect 70786 800 70986 856
rect 71154 800 71262 856
rect 71430 800 71630 856
rect 71798 800 71906 856
rect 72074 800 72274 856
rect 72442 800 72550 856
rect 72718 800 72918 856
rect 73086 800 73194 856
rect 73362 800 73562 856
rect 73730 800 73838 856
rect 74006 800 74206 856
rect 74374 800 74482 856
rect 74650 800 74850 856
rect 75018 800 75126 856
rect 75294 800 75494 856
rect 75662 800 75770 856
rect 75938 800 76138 856
rect 76306 800 76414 856
rect 76582 800 76782 856
rect 76950 800 77058 856
rect 77226 800 77426 856
rect 77594 800 77702 856
rect 77870 800 78070 856
rect 78238 800 78346 856
rect 78514 800 78714 856
rect 78882 800 78990 856
rect 79158 800 79358 856
rect 79526 800 79634 856
rect 79802 800 80002 856
rect 80170 800 80370 856
rect 80538 800 80646 856
rect 80814 800 81014 856
rect 81182 800 81290 856
rect 81458 800 81658 856
rect 81826 800 81934 856
rect 82102 800 82302 856
rect 82470 800 82578 856
rect 82746 800 82946 856
rect 83114 800 83222 856
rect 83390 800 83590 856
rect 83758 800 83866 856
rect 84034 800 84234 856
rect 84402 800 84510 856
rect 84678 800 84878 856
rect 85046 800 85154 856
rect 85322 800 85522 856
rect 85690 800 85798 856
rect 85966 800 86166 856
rect 86334 800 86442 856
rect 86610 800 86810 856
rect 86978 800 87086 856
rect 87254 800 87454 856
rect 87622 800 87730 856
rect 87898 800 88098 856
rect 88266 800 88374 856
rect 88542 800 88742 856
rect 88910 800 89018 856
rect 89186 800 89386 856
rect 89554 800 89662 856
rect 89830 800 90030 856
rect 90198 800 90306 856
rect 90474 800 90674 856
rect 90842 800 90950 856
rect 91118 800 91318 856
rect 91486 800 91594 856
rect 91762 800 91962 856
rect 92130 800 92238 856
rect 92406 800 92606 856
rect 92774 800 92882 856
rect 93050 800 93250 856
rect 93418 800 93526 856
rect 93694 800 93894 856
rect 94062 800 94170 856
rect 94338 800 94538 856
rect 94706 800 94814 856
rect 94982 800 95182 856
rect 95350 800 95458 856
rect 95626 800 95826 856
rect 95994 800 96102 856
rect 96270 800 96470 856
rect 96638 800 96746 856
rect 96914 800 97114 856
rect 97282 800 97390 856
rect 97558 800 97758 856
rect 97926 800 98034 856
rect 98202 800 98402 856
rect 98570 800 98678 856
rect 98846 800 99046 856
rect 99214 800 99322 856
rect 99490 800 99690 856
rect 99858 800 99966 856
rect 100134 800 100334 856
rect 100502 800 100610 856
rect 100778 800 100978 856
rect 101146 800 101254 856
rect 101422 800 101622 856
rect 101790 800 101898 856
rect 102066 800 102266 856
rect 102434 800 102542 856
rect 102710 800 102910 856
rect 103078 800 103186 856
rect 103354 800 103554 856
rect 103722 800 103830 856
rect 103998 800 104198 856
rect 104366 800 104474 856
rect 104642 800 104842 856
rect 105010 800 105118 856
rect 105286 800 105486 856
rect 105654 800 105762 856
rect 105930 800 106130 856
rect 106298 800 106406 856
rect 106574 800 106774 856
rect 106942 800 107142 856
rect 107310 800 107418 856
rect 107586 800 107786 856
rect 107954 800 108062 856
rect 108230 800 108430 856
rect 108598 800 108706 856
rect 108874 800 109074 856
rect 109242 800 109350 856
rect 109518 800 109718 856
rect 109886 800 109994 856
rect 110162 800 110362 856
rect 110530 800 110638 856
rect 110806 800 111006 856
rect 111174 800 111282 856
rect 111450 800 111650 856
rect 111818 800 111926 856
rect 112094 800 112294 856
rect 112462 800 112570 856
rect 112738 800 112938 856
rect 113106 800 113214 856
rect 113382 800 113582 856
rect 113750 800 113858 856
rect 114026 800 114226 856
rect 114394 800 114502 856
rect 114670 800 114870 856
rect 115038 800 115146 856
rect 115314 800 115514 856
rect 115682 800 115790 856
rect 115958 800 116158 856
rect 116326 800 116434 856
rect 116602 800 116802 856
rect 116970 800 117078 856
rect 117246 800 117446 856
rect 117614 800 117722 856
rect 117890 800 118090 856
rect 118258 800 118366 856
rect 118534 800 118734 856
rect 118902 800 119010 856
rect 119178 800 119378 856
rect 119546 800 119654 856
rect 119822 800 120022 856
rect 120190 800 120298 856
rect 120466 800 120666 856
rect 120834 800 120942 856
rect 121110 800 121310 856
rect 121478 800 121586 856
rect 121754 800 121954 856
rect 122122 800 122230 856
rect 122398 800 122598 856
rect 122766 800 122874 856
rect 123042 800 123242 856
rect 123410 800 123518 856
rect 123686 800 123886 856
rect 124054 800 124162 856
rect 124330 800 124530 856
rect 124698 800 124806 856
rect 124974 800 125174 856
rect 125342 800 125450 856
rect 125618 800 125818 856
rect 125986 800 126094 856
rect 126262 800 126462 856
rect 126630 800 126738 856
rect 126906 800 127106 856
rect 127274 800 127382 856
rect 127550 800 127750 856
rect 127918 800 128026 856
rect 128194 800 128394 856
rect 128562 800 128670 856
rect 128838 800 129038 856
rect 129206 800 129314 856
rect 129482 800 129682 856
rect 129850 800 129958 856
rect 130126 800 130326 856
rect 130494 800 130602 856
rect 130770 800 130970 856
rect 131138 800 131246 856
rect 131414 800 131614 856
rect 131782 800 131890 856
rect 132058 800 132258 856
rect 132426 800 132534 856
rect 132702 800 132902 856
rect 133070 800 133178 856
rect 133346 800 133546 856
rect 133714 800 133914 856
rect 134082 800 134190 856
rect 134358 800 134558 856
rect 134726 800 134834 856
rect 135002 800 135202 856
rect 135370 800 135478 856
rect 135646 800 135846 856
rect 136014 800 136122 856
rect 136290 800 136490 856
rect 136658 800 136766 856
rect 136934 800 137134 856
rect 137302 800 137410 856
rect 137578 800 137778 856
rect 137946 800 138054 856
rect 138222 800 138422 856
rect 138590 800 138698 856
rect 138866 800 139066 856
rect 139234 800 139342 856
rect 139510 800 139710 856
rect 139878 800 139986 856
rect 140154 800 140354 856
rect 140522 800 140630 856
rect 140798 800 140998 856
rect 141166 800 141274 856
rect 141442 800 141642 856
rect 141810 800 141918 856
rect 142086 800 142286 856
rect 142454 800 142562 856
rect 142730 800 142930 856
rect 143098 800 143206 856
rect 143374 800 143574 856
rect 143742 800 143850 856
rect 144018 800 144218 856
rect 144386 800 144494 856
rect 144662 800 144862 856
rect 145030 800 145138 856
rect 145306 800 145506 856
rect 145674 800 145782 856
rect 145950 800 146150 856
rect 146318 800 146426 856
rect 146594 800 146794 856
rect 146962 800 147070 856
rect 147238 800 147438 856
rect 147606 800 147714 856
rect 147882 800 148082 856
rect 148250 800 148358 856
rect 148526 800 148726 856
rect 148894 800 149002 856
rect 149170 800 149370 856
rect 149538 800 149646 856
rect 149814 800 150014 856
rect 150182 800 150290 856
rect 150458 800 150658 856
rect 150826 800 150934 856
rect 151102 800 151302 856
rect 151470 800 151578 856
rect 151746 800 151946 856
rect 152114 800 152222 856
rect 152390 800 152590 856
rect 152758 800 152866 856
rect 153034 800 153234 856
rect 153402 800 153510 856
rect 153678 800 153878 856
rect 154046 800 154154 856
rect 154322 800 154522 856
rect 154690 800 154798 856
rect 154966 800 155166 856
rect 155334 800 155442 856
rect 155610 800 155810 856
rect 155978 800 156086 856
rect 156254 800 156454 856
rect 156622 800 156730 856
rect 156898 800 157098 856
rect 157266 800 157374 856
rect 157542 800 157742 856
rect 157910 800 158018 856
<< metal3 >>
rect 0 150968 800 151088
rect 159200 146616 160000 146736
rect 0 133152 800 133272
rect 159200 119960 160000 120080
rect 0 115472 800 115592
rect 0 97656 800 97776
rect 159200 93304 160000 93424
rect 0 79840 800 79960
rect 159200 66648 160000 66768
rect 0 62160 800 62280
rect 0 44344 800 44464
rect 159200 39992 160000 40112
rect 0 26528 800 26648
rect 159200 13336 160000 13456
rect 0 8848 800 8968
<< obsm3 >>
rect 105 151168 158128 157793
rect 880 150888 158128 151168
rect 105 133352 158128 150888
rect 880 133072 158128 133352
rect 105 115672 158128 133072
rect 880 115392 158128 115672
rect 105 97856 158128 115392
rect 880 97576 158128 97856
rect 105 80040 158128 97576
rect 880 79760 158128 80040
rect 105 62360 158128 79760
rect 880 62080 158128 62360
rect 105 44544 158128 62080
rect 880 44264 158128 44544
rect 105 26728 158128 44264
rect 880 26448 158128 26728
rect 105 9048 158128 26448
rect 880 8768 158128 9048
rect 105 851 158128 8768
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
<< obsm4 >>
rect 30235 2128 158128 157808
<< labels >>
rlabel metal3 s 0 8848 800 8968 6 analog_io[0]
port 1 nsew default bidirectional
rlabel metal3 s 159200 66648 160000 66768 6 analog_io[10]
port 2 nsew default bidirectional
rlabel metal2 s 150254 159200 150310 160000 6 analog_io[11]
port 3 nsew default bidirectional
rlabel metal2 s 151542 159200 151598 160000 6 analog_io[12]
port 4 nsew default bidirectional
rlabel metal3 s 159200 93304 160000 93424 6 analog_io[13]
port 5 nsew default bidirectional
rlabel metal2 s 158442 0 158498 800 6 analog_io[14]
port 6 nsew default bidirectional
rlabel metal2 s 152830 159200 152886 160000 6 analog_io[15]
port 7 nsew default bidirectional
rlabel metal2 s 158718 0 158774 800 6 analog_io[16]
port 8 nsew default bidirectional
rlabel metal2 s 159086 0 159142 800 6 analog_io[17]
port 9 nsew default bidirectional
rlabel metal2 s 159362 0 159418 800 6 analog_io[18]
port 10 nsew default bidirectional
rlabel metal3 s 159200 119960 160000 120080 6 analog_io[19]
port 11 nsew default bidirectional
rlabel metal3 s 0 26528 800 26648 6 analog_io[1]
port 12 nsew default bidirectional
rlabel metal2 s 154118 159200 154174 160000 6 analog_io[20]
port 13 nsew default bidirectional
rlabel metal3 s 0 97656 800 97776 6 analog_io[21]
port 14 nsew default bidirectional
rlabel metal3 s 0 115472 800 115592 6 analog_io[22]
port 15 nsew default bidirectional
rlabel metal3 s 159200 146616 160000 146736 6 analog_io[23]
port 16 nsew default bidirectional
rlabel metal3 s 0 133152 800 133272 6 analog_io[24]
port 17 nsew default bidirectional
rlabel metal2 s 155406 159200 155462 160000 6 analog_io[25]
port 18 nsew default bidirectional
rlabel metal2 s 156694 159200 156750 160000 6 analog_io[26]
port 19 nsew default bidirectional
rlabel metal2 s 157982 159200 158038 160000 6 analog_io[27]
port 20 nsew default bidirectional
rlabel metal3 s 0 150968 800 151088 6 analog_io[28]
port 21 nsew default bidirectional
rlabel metal2 s 159730 0 159786 800 6 analog_io[29]
port 22 nsew default bidirectional
rlabel metal3 s 0 44344 800 44464 6 analog_io[2]
port 23 nsew default bidirectional
rlabel metal2 s 159270 159200 159326 160000 6 analog_io[30]
port 24 nsew default bidirectional
rlabel metal3 s 0 62160 800 62280 6 analog_io[3]
port 25 nsew default bidirectional
rlabel metal3 s 159200 13336 160000 13456 6 analog_io[4]
port 26 nsew default bidirectional
rlabel metal3 s 159200 39992 160000 40112 6 analog_io[5]
port 27 nsew default bidirectional
rlabel metal2 s 147678 159200 147734 160000 6 analog_io[6]
port 28 nsew default bidirectional
rlabel metal2 s 148966 159200 149022 160000 6 analog_io[7]
port 29 nsew default bidirectional
rlabel metal3 s 0 79840 800 79960 6 analog_io[8]
port 30 nsew default bidirectional
rlabel metal2 s 158074 0 158130 800 6 analog_io[9]
port 31 nsew default bidirectional
rlabel metal2 s 662 159200 718 160000 6 io_in[0]
port 32 nsew default input
rlabel metal2 s 39302 159200 39358 160000 6 io_in[10]
port 33 nsew default input
rlabel metal2 s 43166 159200 43222 160000 6 io_in[11]
port 34 nsew default input
rlabel metal2 s 47030 159200 47086 160000 6 io_in[12]
port 35 nsew default input
rlabel metal2 s 50894 159200 50950 160000 6 io_in[13]
port 36 nsew default input
rlabel metal2 s 54850 159200 54906 160000 6 io_in[14]
port 37 nsew default input
rlabel metal2 s 58714 159200 58770 160000 6 io_in[15]
port 38 nsew default input
rlabel metal2 s 62578 159200 62634 160000 6 io_in[16]
port 39 nsew default input
rlabel metal2 s 66442 159200 66498 160000 6 io_in[17]
port 40 nsew default input
rlabel metal2 s 70306 159200 70362 160000 6 io_in[18]
port 41 nsew default input
rlabel metal2 s 74170 159200 74226 160000 6 io_in[19]
port 42 nsew default input
rlabel metal2 s 4526 159200 4582 160000 6 io_in[1]
port 43 nsew default input
rlabel metal2 s 78034 159200 78090 160000 6 io_in[20]
port 44 nsew default input
rlabel metal2 s 81898 159200 81954 160000 6 io_in[21]
port 45 nsew default input
rlabel metal2 s 85762 159200 85818 160000 6 io_in[22]
port 46 nsew default input
rlabel metal2 s 89626 159200 89682 160000 6 io_in[23]
port 47 nsew default input
rlabel metal2 s 93490 159200 93546 160000 6 io_in[24]
port 48 nsew default input
rlabel metal2 s 97354 159200 97410 160000 6 io_in[25]
port 49 nsew default input
rlabel metal2 s 101218 159200 101274 160000 6 io_in[26]
port 50 nsew default input
rlabel metal2 s 105082 159200 105138 160000 6 io_in[27]
port 51 nsew default input
rlabel metal2 s 109038 159200 109094 160000 6 io_in[28]
port 52 nsew default input
rlabel metal2 s 112902 159200 112958 160000 6 io_in[29]
port 53 nsew default input
rlabel metal2 s 8390 159200 8446 160000 6 io_in[2]
port 54 nsew default input
rlabel metal2 s 116766 159200 116822 160000 6 io_in[30]
port 55 nsew default input
rlabel metal2 s 120630 159200 120686 160000 6 io_in[31]
port 56 nsew default input
rlabel metal2 s 124494 159200 124550 160000 6 io_in[32]
port 57 nsew default input
rlabel metal2 s 128358 159200 128414 160000 6 io_in[33]
port 58 nsew default input
rlabel metal2 s 132222 159200 132278 160000 6 io_in[34]
port 59 nsew default input
rlabel metal2 s 136086 159200 136142 160000 6 io_in[35]
port 60 nsew default input
rlabel metal2 s 139950 159200 140006 160000 6 io_in[36]
port 61 nsew default input
rlabel metal2 s 143814 159200 143870 160000 6 io_in[37]
port 62 nsew default input
rlabel metal2 s 12254 159200 12310 160000 6 io_in[3]
port 63 nsew default input
rlabel metal2 s 16118 159200 16174 160000 6 io_in[4]
port 64 nsew default input
rlabel metal2 s 19982 159200 20038 160000 6 io_in[5]
port 65 nsew default input
rlabel metal2 s 23846 159200 23902 160000 6 io_in[6]
port 66 nsew default input
rlabel metal2 s 27710 159200 27766 160000 6 io_in[7]
port 67 nsew default input
rlabel metal2 s 31574 159200 31630 160000 6 io_in[8]
port 68 nsew default input
rlabel metal2 s 35438 159200 35494 160000 6 io_in[9]
port 69 nsew default input
rlabel metal2 s 1950 159200 2006 160000 6 io_oeb[0]
port 70 nsew default output
rlabel metal2 s 40590 159200 40646 160000 6 io_oeb[10]
port 71 nsew default output
rlabel metal2 s 44454 159200 44510 160000 6 io_oeb[11]
port 72 nsew default output
rlabel metal2 s 48318 159200 48374 160000 6 io_oeb[12]
port 73 nsew default output
rlabel metal2 s 52182 159200 52238 160000 6 io_oeb[13]
port 74 nsew default output
rlabel metal2 s 56138 159200 56194 160000 6 io_oeb[14]
port 75 nsew default output
rlabel metal2 s 60002 159200 60058 160000 6 io_oeb[15]
port 76 nsew default output
rlabel metal2 s 63866 159200 63922 160000 6 io_oeb[16]
port 77 nsew default output
rlabel metal2 s 67730 159200 67786 160000 6 io_oeb[17]
port 78 nsew default output
rlabel metal2 s 71594 159200 71650 160000 6 io_oeb[18]
port 79 nsew default output
rlabel metal2 s 75458 159200 75514 160000 6 io_oeb[19]
port 80 nsew default output
rlabel metal2 s 5814 159200 5870 160000 6 io_oeb[1]
port 81 nsew default output
rlabel metal2 s 79322 159200 79378 160000 6 io_oeb[20]
port 82 nsew default output
rlabel metal2 s 83186 159200 83242 160000 6 io_oeb[21]
port 83 nsew default output
rlabel metal2 s 87050 159200 87106 160000 6 io_oeb[22]
port 84 nsew default output
rlabel metal2 s 90914 159200 90970 160000 6 io_oeb[23]
port 85 nsew default output
rlabel metal2 s 94778 159200 94834 160000 6 io_oeb[24]
port 86 nsew default output
rlabel metal2 s 98642 159200 98698 160000 6 io_oeb[25]
port 87 nsew default output
rlabel metal2 s 102506 159200 102562 160000 6 io_oeb[26]
port 88 nsew default output
rlabel metal2 s 106370 159200 106426 160000 6 io_oeb[27]
port 89 nsew default output
rlabel metal2 s 110326 159200 110382 160000 6 io_oeb[28]
port 90 nsew default output
rlabel metal2 s 114190 159200 114246 160000 6 io_oeb[29]
port 91 nsew default output
rlabel metal2 s 9678 159200 9734 160000 6 io_oeb[2]
port 92 nsew default output
rlabel metal2 s 118054 159200 118110 160000 6 io_oeb[30]
port 93 nsew default output
rlabel metal2 s 121918 159200 121974 160000 6 io_oeb[31]
port 94 nsew default output
rlabel metal2 s 125782 159200 125838 160000 6 io_oeb[32]
port 95 nsew default output
rlabel metal2 s 129646 159200 129702 160000 6 io_oeb[33]
port 96 nsew default output
rlabel metal2 s 133510 159200 133566 160000 6 io_oeb[34]
port 97 nsew default output
rlabel metal2 s 137374 159200 137430 160000 6 io_oeb[35]
port 98 nsew default output
rlabel metal2 s 141238 159200 141294 160000 6 io_oeb[36]
port 99 nsew default output
rlabel metal2 s 145102 159200 145158 160000 6 io_oeb[37]
port 100 nsew default output
rlabel metal2 s 13542 159200 13598 160000 6 io_oeb[3]
port 101 nsew default output
rlabel metal2 s 17406 159200 17462 160000 6 io_oeb[4]
port 102 nsew default output
rlabel metal2 s 21270 159200 21326 160000 6 io_oeb[5]
port 103 nsew default output
rlabel metal2 s 25134 159200 25190 160000 6 io_oeb[6]
port 104 nsew default output
rlabel metal2 s 28998 159200 29054 160000 6 io_oeb[7]
port 105 nsew default output
rlabel metal2 s 32862 159200 32918 160000 6 io_oeb[8]
port 106 nsew default output
rlabel metal2 s 36726 159200 36782 160000 6 io_oeb[9]
port 107 nsew default output
rlabel metal2 s 3238 159200 3294 160000 6 io_out[0]
port 108 nsew default output
rlabel metal2 s 41878 159200 41934 160000 6 io_out[10]
port 109 nsew default output
rlabel metal2 s 45742 159200 45798 160000 6 io_out[11]
port 110 nsew default output
rlabel metal2 s 49606 159200 49662 160000 6 io_out[12]
port 111 nsew default output
rlabel metal2 s 53470 159200 53526 160000 6 io_out[13]
port 112 nsew default output
rlabel metal2 s 57426 159200 57482 160000 6 io_out[14]
port 113 nsew default output
rlabel metal2 s 61290 159200 61346 160000 6 io_out[15]
port 114 nsew default output
rlabel metal2 s 65154 159200 65210 160000 6 io_out[16]
port 115 nsew default output
rlabel metal2 s 69018 159200 69074 160000 6 io_out[17]
port 116 nsew default output
rlabel metal2 s 72882 159200 72938 160000 6 io_out[18]
port 117 nsew default output
rlabel metal2 s 76746 159200 76802 160000 6 io_out[19]
port 118 nsew default output
rlabel metal2 s 7102 159200 7158 160000 6 io_out[1]
port 119 nsew default output
rlabel metal2 s 80610 159200 80666 160000 6 io_out[20]
port 120 nsew default output
rlabel metal2 s 84474 159200 84530 160000 6 io_out[21]
port 121 nsew default output
rlabel metal2 s 88338 159200 88394 160000 6 io_out[22]
port 122 nsew default output
rlabel metal2 s 92202 159200 92258 160000 6 io_out[23]
port 123 nsew default output
rlabel metal2 s 96066 159200 96122 160000 6 io_out[24]
port 124 nsew default output
rlabel metal2 s 99930 159200 99986 160000 6 io_out[25]
port 125 nsew default output
rlabel metal2 s 103794 159200 103850 160000 6 io_out[26]
port 126 nsew default output
rlabel metal2 s 107750 159200 107806 160000 6 io_out[27]
port 127 nsew default output
rlabel metal2 s 111614 159200 111670 160000 6 io_out[28]
port 128 nsew default output
rlabel metal2 s 115478 159200 115534 160000 6 io_out[29]
port 129 nsew default output
rlabel metal2 s 10966 159200 11022 160000 6 io_out[2]
port 130 nsew default output
rlabel metal2 s 119342 159200 119398 160000 6 io_out[30]
port 131 nsew default output
rlabel metal2 s 123206 159200 123262 160000 6 io_out[31]
port 132 nsew default output
rlabel metal2 s 127070 159200 127126 160000 6 io_out[32]
port 133 nsew default output
rlabel metal2 s 130934 159200 130990 160000 6 io_out[33]
port 134 nsew default output
rlabel metal2 s 134798 159200 134854 160000 6 io_out[34]
port 135 nsew default output
rlabel metal2 s 138662 159200 138718 160000 6 io_out[35]
port 136 nsew default output
rlabel metal2 s 142526 159200 142582 160000 6 io_out[36]
port 137 nsew default output
rlabel metal2 s 146390 159200 146446 160000 6 io_out[37]
port 138 nsew default output
rlabel metal2 s 14830 159200 14886 160000 6 io_out[3]
port 139 nsew default output
rlabel metal2 s 18694 159200 18750 160000 6 io_out[4]
port 140 nsew default output
rlabel metal2 s 22558 159200 22614 160000 6 io_out[5]
port 141 nsew default output
rlabel metal2 s 26422 159200 26478 160000 6 io_out[6]
port 142 nsew default output
rlabel metal2 s 30286 159200 30342 160000 6 io_out[7]
port 143 nsew default output
rlabel metal2 s 34150 159200 34206 160000 6 io_out[8]
port 144 nsew default output
rlabel metal2 s 38014 159200 38070 160000 6 io_out[9]
port 145 nsew default output
rlabel metal2 s 34242 0 34298 800 6 la_data_in[0]
port 146 nsew default input
rlabel metal2 s 131026 0 131082 800 6 la_data_in[100]
port 147 nsew default input
rlabel metal2 s 131946 0 132002 800 6 la_data_in[101]
port 148 nsew default input
rlabel metal2 s 132958 0 133014 800 6 la_data_in[102]
port 149 nsew default input
rlabel metal2 s 133970 0 134026 800 6 la_data_in[103]
port 150 nsew default input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[104]
port 151 nsew default input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[105]
port 152 nsew default input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[106]
port 153 nsew default input
rlabel metal2 s 137834 0 137890 800 6 la_data_in[107]
port 154 nsew default input
rlabel metal2 s 138754 0 138810 800 6 la_data_in[108]
port 155 nsew default input
rlabel metal2 s 139766 0 139822 800 6 la_data_in[109]
port 156 nsew default input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[10]
port 157 nsew default input
rlabel metal2 s 140686 0 140742 800 6 la_data_in[110]
port 158 nsew default input
rlabel metal2 s 141698 0 141754 800 6 la_data_in[111]
port 159 nsew default input
rlabel metal2 s 142618 0 142674 800 6 la_data_in[112]
port 160 nsew default input
rlabel metal2 s 143630 0 143686 800 6 la_data_in[113]
port 161 nsew default input
rlabel metal2 s 144550 0 144606 800 6 la_data_in[114]
port 162 nsew default input
rlabel metal2 s 145562 0 145618 800 6 la_data_in[115]
port 163 nsew default input
rlabel metal2 s 146482 0 146538 800 6 la_data_in[116]
port 164 nsew default input
rlabel metal2 s 147494 0 147550 800 6 la_data_in[117]
port 165 nsew default input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[118]
port 166 nsew default input
rlabel metal2 s 149426 0 149482 800 6 la_data_in[119]
port 167 nsew default input
rlabel metal2 s 44914 0 44970 800 6 la_data_in[11]
port 168 nsew default input
rlabel metal2 s 150346 0 150402 800 6 la_data_in[120]
port 169 nsew default input
rlabel metal2 s 151358 0 151414 800 6 la_data_in[121]
port 170 nsew default input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[122]
port 171 nsew default input
rlabel metal2 s 153290 0 153346 800 6 la_data_in[123]
port 172 nsew default input
rlabel metal2 s 154210 0 154266 800 6 la_data_in[124]
port 173 nsew default input
rlabel metal2 s 155222 0 155278 800 6 la_data_in[125]
port 174 nsew default input
rlabel metal2 s 156142 0 156198 800 6 la_data_in[126]
port 175 nsew default input
rlabel metal2 s 157154 0 157210 800 6 la_data_in[127]
port 176 nsew default input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[12]
port 177 nsew default input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[13]
port 178 nsew default input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[14]
port 179 nsew default input
rlabel metal2 s 48778 0 48834 800 6 la_data_in[15]
port 180 nsew default input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[16]
port 181 nsew default input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[17]
port 182 nsew default input
rlabel metal2 s 51630 0 51686 800 6 la_data_in[18]
port 183 nsew default input
rlabel metal2 s 52642 0 52698 800 6 la_data_in[19]
port 184 nsew default input
rlabel metal2 s 35254 0 35310 800 6 la_data_in[1]
port 185 nsew default input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[20]
port 186 nsew default input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[21]
port 187 nsew default input
rlabel metal2 s 55586 0 55642 800 6 la_data_in[22]
port 188 nsew default input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[23]
port 189 nsew default input
rlabel metal2 s 57518 0 57574 800 6 la_data_in[24]
port 190 nsew default input
rlabel metal2 s 58438 0 58494 800 6 la_data_in[25]
port 191 nsew default input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[26]
port 192 nsew default input
rlabel metal2 s 60370 0 60426 800 6 la_data_in[27]
port 193 nsew default input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[28]
port 194 nsew default input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[29]
port 195 nsew default input
rlabel metal2 s 36174 0 36230 800 6 la_data_in[2]
port 196 nsew default input
rlabel metal2 s 63314 0 63370 800 6 la_data_in[30]
port 197 nsew default input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[31]
port 198 nsew default input
rlabel metal2 s 65246 0 65302 800 6 la_data_in[32]
port 199 nsew default input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[33]
port 200 nsew default input
rlabel metal2 s 67178 0 67234 800 6 la_data_in[34]
port 201 nsew default input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[35]
port 202 nsew default input
rlabel metal2 s 69110 0 69166 800 6 la_data_in[36]
port 203 nsew default input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[37]
port 204 nsew default input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[38]
port 205 nsew default input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[39]
port 206 nsew default input
rlabel metal2 s 37186 0 37242 800 6 la_data_in[3]
port 207 nsew default input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[40]
port 208 nsew default input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[41]
port 209 nsew default input
rlabel metal2 s 74906 0 74962 800 6 la_data_in[42]
port 210 nsew default input
rlabel metal2 s 75826 0 75882 800 6 la_data_in[43]
port 211 nsew default input
rlabel metal2 s 76838 0 76894 800 6 la_data_in[44]
port 212 nsew default input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[45]
port 213 nsew default input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[46]
port 214 nsew default input
rlabel metal2 s 79690 0 79746 800 6 la_data_in[47]
port 215 nsew default input
rlabel metal2 s 80702 0 80758 800 6 la_data_in[48]
port 216 nsew default input
rlabel metal2 s 81714 0 81770 800 6 la_data_in[49]
port 217 nsew default input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[4]
port 218 nsew default input
rlabel metal2 s 82634 0 82690 800 6 la_data_in[50]
port 219 nsew default input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[51]
port 220 nsew default input
rlabel metal2 s 84566 0 84622 800 6 la_data_in[52]
port 221 nsew default input
rlabel metal2 s 85578 0 85634 800 6 la_data_in[53]
port 222 nsew default input
rlabel metal2 s 86498 0 86554 800 6 la_data_in[54]
port 223 nsew default input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[55]
port 224 nsew default input
rlabel metal2 s 88430 0 88486 800 6 la_data_in[56]
port 225 nsew default input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[57]
port 226 nsew default input
rlabel metal2 s 90362 0 90418 800 6 la_data_in[58]
port 227 nsew default input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[59]
port 228 nsew default input
rlabel metal2 s 39118 0 39174 800 6 la_data_in[5]
port 229 nsew default input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[60]
port 230 nsew default input
rlabel metal2 s 93306 0 93362 800 6 la_data_in[61]
port 231 nsew default input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[62]
port 232 nsew default input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[63]
port 233 nsew default input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[64]
port 234 nsew default input
rlabel metal2 s 97170 0 97226 800 6 la_data_in[65]
port 235 nsew default input
rlabel metal2 s 98090 0 98146 800 6 la_data_in[66]
port 236 nsew default input
rlabel metal2 s 99102 0 99158 800 6 la_data_in[67]
port 237 nsew default input
rlabel metal2 s 100022 0 100078 800 6 la_data_in[68]
port 238 nsew default input
rlabel metal2 s 101034 0 101090 800 6 la_data_in[69]
port 239 nsew default input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[6]
port 240 nsew default input
rlabel metal2 s 101954 0 102010 800 6 la_data_in[70]
port 241 nsew default input
rlabel metal2 s 102966 0 103022 800 6 la_data_in[71]
port 242 nsew default input
rlabel metal2 s 103886 0 103942 800 6 la_data_in[72]
port 243 nsew default input
rlabel metal2 s 104898 0 104954 800 6 la_data_in[73]
port 244 nsew default input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[74]
port 245 nsew default input
rlabel metal2 s 106830 0 106886 800 6 la_data_in[75]
port 246 nsew default input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[76]
port 247 nsew default input
rlabel metal2 s 108762 0 108818 800 6 la_data_in[77]
port 248 nsew default input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[78]
port 249 nsew default input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[79]
port 250 nsew default input
rlabel metal2 s 41050 0 41106 800 6 la_data_in[7]
port 251 nsew default input
rlabel metal2 s 111706 0 111762 800 6 la_data_in[80]
port 252 nsew default input
rlabel metal2 s 112626 0 112682 800 6 la_data_in[81]
port 253 nsew default input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[82]
port 254 nsew default input
rlabel metal2 s 114558 0 114614 800 6 la_data_in[83]
port 255 nsew default input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[84]
port 256 nsew default input
rlabel metal2 s 116490 0 116546 800 6 la_data_in[85]
port 257 nsew default input
rlabel metal2 s 117502 0 117558 800 6 la_data_in[86]
port 258 nsew default input
rlabel metal2 s 118422 0 118478 800 6 la_data_in[87]
port 259 nsew default input
rlabel metal2 s 119434 0 119490 800 6 la_data_in[88]
port 260 nsew default input
rlabel metal2 s 120354 0 120410 800 6 la_data_in[89]
port 261 nsew default input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[8]
port 262 nsew default input
rlabel metal2 s 121366 0 121422 800 6 la_data_in[90]
port 263 nsew default input
rlabel metal2 s 122286 0 122342 800 6 la_data_in[91]
port 264 nsew default input
rlabel metal2 s 123298 0 123354 800 6 la_data_in[92]
port 265 nsew default input
rlabel metal2 s 124218 0 124274 800 6 la_data_in[93]
port 266 nsew default input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[94]
port 267 nsew default input
rlabel metal2 s 126150 0 126206 800 6 la_data_in[95]
port 268 nsew default input
rlabel metal2 s 127162 0 127218 800 6 la_data_in[96]
port 269 nsew default input
rlabel metal2 s 128082 0 128138 800 6 la_data_in[97]
port 270 nsew default input
rlabel metal2 s 129094 0 129150 800 6 la_data_in[98]
port 271 nsew default input
rlabel metal2 s 130014 0 130070 800 6 la_data_in[99]
port 272 nsew default input
rlabel metal2 s 42982 0 43038 800 6 la_data_in[9]
port 273 nsew default input
rlabel metal2 s 34610 0 34666 800 6 la_data_out[0]
port 274 nsew default output
rlabel metal2 s 131302 0 131358 800 6 la_data_out[100]
port 275 nsew default output
rlabel metal2 s 132314 0 132370 800 6 la_data_out[101]
port 276 nsew default output
rlabel metal2 s 133234 0 133290 800 6 la_data_out[102]
port 277 nsew default output
rlabel metal2 s 134246 0 134302 800 6 la_data_out[103]
port 278 nsew default output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[104]
port 279 nsew default output
rlabel metal2 s 136178 0 136234 800 6 la_data_out[105]
port 280 nsew default output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[106]
port 281 nsew default output
rlabel metal2 s 138110 0 138166 800 6 la_data_out[107]
port 282 nsew default output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[108]
port 283 nsew default output
rlabel metal2 s 140042 0 140098 800 6 la_data_out[109]
port 284 nsew default output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[10]
port 285 nsew default output
rlabel metal2 s 141054 0 141110 800 6 la_data_out[110]
port 286 nsew default output
rlabel metal2 s 141974 0 142030 800 6 la_data_out[111]
port 287 nsew default output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[112]
port 288 nsew default output
rlabel metal2 s 143906 0 143962 800 6 la_data_out[113]
port 289 nsew default output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[114]
port 290 nsew default output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[115]
port 291 nsew default output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[116]
port 292 nsew default output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[117]
port 293 nsew default output
rlabel metal2 s 148782 0 148838 800 6 la_data_out[118]
port 294 nsew default output
rlabel metal2 s 149702 0 149758 800 6 la_data_out[119]
port 295 nsew default output
rlabel metal2 s 45190 0 45246 800 6 la_data_out[11]
port 296 nsew default output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[120]
port 297 nsew default output
rlabel metal2 s 151634 0 151690 800 6 la_data_out[121]
port 298 nsew default output
rlabel metal2 s 152646 0 152702 800 6 la_data_out[122]
port 299 nsew default output
rlabel metal2 s 153566 0 153622 800 6 la_data_out[123]
port 300 nsew default output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[124]
port 301 nsew default output
rlabel metal2 s 155498 0 155554 800 6 la_data_out[125]
port 302 nsew default output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[126]
port 303 nsew default output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[127]
port 304 nsew default output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[12]
port 305 nsew default output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[13]
port 306 nsew default output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[14]
port 307 nsew default output
rlabel metal2 s 49054 0 49110 800 6 la_data_out[15]
port 308 nsew default output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[16]
port 309 nsew default output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[17]
port 310 nsew default output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[18]
port 311 nsew default output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[19]
port 312 nsew default output
rlabel metal2 s 35530 0 35586 800 6 la_data_out[1]
port 313 nsew default output
rlabel metal2 s 53930 0 53986 800 6 la_data_out[20]
port 314 nsew default output
rlabel metal2 s 54942 0 54998 800 6 la_data_out[21]
port 315 nsew default output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[22]
port 316 nsew default output
rlabel metal2 s 56874 0 56930 800 6 la_data_out[23]
port 317 nsew default output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[24]
port 318 nsew default output
rlabel metal2 s 58806 0 58862 800 6 la_data_out[25]
port 319 nsew default output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[26]
port 320 nsew default output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[27]
port 321 nsew default output
rlabel metal2 s 61658 0 61714 800 6 la_data_out[28]
port 322 nsew default output
rlabel metal2 s 62670 0 62726 800 6 la_data_out[29]
port 323 nsew default output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[2]
port 324 nsew default output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[30]
port 325 nsew default output
rlabel metal2 s 64602 0 64658 800 6 la_data_out[31]
port 326 nsew default output
rlabel metal2 s 65522 0 65578 800 6 la_data_out[32]
port 327 nsew default output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[33]
port 328 nsew default output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[34]
port 329 nsew default output
rlabel metal2 s 68466 0 68522 800 6 la_data_out[35]
port 330 nsew default output
rlabel metal2 s 69386 0 69442 800 6 la_data_out[36]
port 331 nsew default output
rlabel metal2 s 70398 0 70454 800 6 la_data_out[37]
port 332 nsew default output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[38]
port 333 nsew default output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[39]
port 334 nsew default output
rlabel metal2 s 37462 0 37518 800 6 la_data_out[3]
port 335 nsew default output
rlabel metal2 s 73250 0 73306 800 6 la_data_out[40]
port 336 nsew default output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[41]
port 337 nsew default output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[42]
port 338 nsew default output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[43]
port 339 nsew default output
rlabel metal2 s 77114 0 77170 800 6 la_data_out[44]
port 340 nsew default output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[45]
port 341 nsew default output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[46]
port 342 nsew default output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[47]
port 343 nsew default output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[48]
port 344 nsew default output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[49]
port 345 nsew default output
rlabel metal2 s 38474 0 38530 800 6 la_data_out[4]
port 346 nsew default output
rlabel metal2 s 83002 0 83058 800 6 la_data_out[50]
port 347 nsew default output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[51]
port 348 nsew default output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[52]
port 349 nsew default output
rlabel metal2 s 85854 0 85910 800 6 la_data_out[53]
port 350 nsew default output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[54]
port 351 nsew default output
rlabel metal2 s 87786 0 87842 800 6 la_data_out[55]
port 352 nsew default output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[56]
port 353 nsew default output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[57]
port 354 nsew default output
rlabel metal2 s 90730 0 90786 800 6 la_data_out[58]
port 355 nsew default output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[59]
port 356 nsew default output
rlabel metal2 s 39394 0 39450 800 6 la_data_out[5]
port 357 nsew default output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[60]
port 358 nsew default output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[61]
port 359 nsew default output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[62]
port 360 nsew default output
rlabel metal2 s 95514 0 95570 800 6 la_data_out[63]
port 361 nsew default output
rlabel metal2 s 96526 0 96582 800 6 la_data_out[64]
port 362 nsew default output
rlabel metal2 s 97446 0 97502 800 6 la_data_out[65]
port 363 nsew default output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[66]
port 364 nsew default output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[67]
port 365 nsew default output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[68]
port 366 nsew default output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[69]
port 367 nsew default output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[6]
port 368 nsew default output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[70]
port 369 nsew default output
rlabel metal2 s 103242 0 103298 800 6 la_data_out[71]
port 370 nsew default output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[72]
port 371 nsew default output
rlabel metal2 s 105174 0 105230 800 6 la_data_out[73]
port 372 nsew default output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[74]
port 373 nsew default output
rlabel metal2 s 107198 0 107254 800 6 la_data_out[75]
port 374 nsew default output
rlabel metal2 s 108118 0 108174 800 6 la_data_out[76]
port 375 nsew default output
rlabel metal2 s 109130 0 109186 800 6 la_data_out[77]
port 376 nsew default output
rlabel metal2 s 110050 0 110106 800 6 la_data_out[78]
port 377 nsew default output
rlabel metal2 s 111062 0 111118 800 6 la_data_out[79]
port 378 nsew default output
rlabel metal2 s 41326 0 41382 800 6 la_data_out[7]
port 379 nsew default output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[80]
port 380 nsew default output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[81]
port 381 nsew default output
rlabel metal2 s 113914 0 113970 800 6 la_data_out[82]
port 382 nsew default output
rlabel metal2 s 114926 0 114982 800 6 la_data_out[83]
port 383 nsew default output
rlabel metal2 s 115846 0 115902 800 6 la_data_out[84]
port 384 nsew default output
rlabel metal2 s 116858 0 116914 800 6 la_data_out[85]
port 385 nsew default output
rlabel metal2 s 117778 0 117834 800 6 la_data_out[86]
port 386 nsew default output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[87]
port 387 nsew default output
rlabel metal2 s 119710 0 119766 800 6 la_data_out[88]
port 388 nsew default output
rlabel metal2 s 120722 0 120778 800 6 la_data_out[89]
port 389 nsew default output
rlabel metal2 s 42338 0 42394 800 6 la_data_out[8]
port 390 nsew default output
rlabel metal2 s 121642 0 121698 800 6 la_data_out[90]
port 391 nsew default output
rlabel metal2 s 122654 0 122710 800 6 la_data_out[91]
port 392 nsew default output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[92]
port 393 nsew default output
rlabel metal2 s 124586 0 124642 800 6 la_data_out[93]
port 394 nsew default output
rlabel metal2 s 125506 0 125562 800 6 la_data_out[94]
port 395 nsew default output
rlabel metal2 s 126518 0 126574 800 6 la_data_out[95]
port 396 nsew default output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[96]
port 397 nsew default output
rlabel metal2 s 128450 0 128506 800 6 la_data_out[97]
port 398 nsew default output
rlabel metal2 s 129370 0 129426 800 6 la_data_out[98]
port 399 nsew default output
rlabel metal2 s 130382 0 130438 800 6 la_data_out[99]
port 400 nsew default output
rlabel metal2 s 43258 0 43314 800 6 la_data_out[9]
port 401 nsew default output
rlabel metal2 s 34886 0 34942 800 6 la_oen[0]
port 402 nsew default input
rlabel metal2 s 131670 0 131726 800 6 la_oen[100]
port 403 nsew default input
rlabel metal2 s 132590 0 132646 800 6 la_oen[101]
port 404 nsew default input
rlabel metal2 s 133602 0 133658 800 6 la_oen[102]
port 405 nsew default input
rlabel metal2 s 134614 0 134670 800 6 la_oen[103]
port 406 nsew default input
rlabel metal2 s 135534 0 135590 800 6 la_oen[104]
port 407 nsew default input
rlabel metal2 s 136546 0 136602 800 6 la_oen[105]
port 408 nsew default input
rlabel metal2 s 137466 0 137522 800 6 la_oen[106]
port 409 nsew default input
rlabel metal2 s 138478 0 138534 800 6 la_oen[107]
port 410 nsew default input
rlabel metal2 s 139398 0 139454 800 6 la_oen[108]
port 411 nsew default input
rlabel metal2 s 140410 0 140466 800 6 la_oen[109]
port 412 nsew default input
rlabel metal2 s 44546 0 44602 800 6 la_oen[10]
port 413 nsew default input
rlabel metal2 s 141330 0 141386 800 6 la_oen[110]
port 414 nsew default input
rlabel metal2 s 142342 0 142398 800 6 la_oen[111]
port 415 nsew default input
rlabel metal2 s 143262 0 143318 800 6 la_oen[112]
port 416 nsew default input
rlabel metal2 s 144274 0 144330 800 6 la_oen[113]
port 417 nsew default input
rlabel metal2 s 145194 0 145250 800 6 la_oen[114]
port 418 nsew default input
rlabel metal2 s 146206 0 146262 800 6 la_oen[115]
port 419 nsew default input
rlabel metal2 s 147126 0 147182 800 6 la_oen[116]
port 420 nsew default input
rlabel metal2 s 148138 0 148194 800 6 la_oen[117]
port 421 nsew default input
rlabel metal2 s 149058 0 149114 800 6 la_oen[118]
port 422 nsew default input
rlabel metal2 s 150070 0 150126 800 6 la_oen[119]
port 423 nsew default input
rlabel metal2 s 45558 0 45614 800 6 la_oen[11]
port 424 nsew default input
rlabel metal2 s 150990 0 151046 800 6 la_oen[120]
port 425 nsew default input
rlabel metal2 s 152002 0 152058 800 6 la_oen[121]
port 426 nsew default input
rlabel metal2 s 152922 0 152978 800 6 la_oen[122]
port 427 nsew default input
rlabel metal2 s 153934 0 153990 800 6 la_oen[123]
port 428 nsew default input
rlabel metal2 s 154854 0 154910 800 6 la_oen[124]
port 429 nsew default input
rlabel metal2 s 155866 0 155922 800 6 la_oen[125]
port 430 nsew default input
rlabel metal2 s 156786 0 156842 800 6 la_oen[126]
port 431 nsew default input
rlabel metal2 s 157798 0 157854 800 6 la_oen[127]
port 432 nsew default input
rlabel metal2 s 46478 0 46534 800 6 la_oen[12]
port 433 nsew default input
rlabel metal2 s 47490 0 47546 800 6 la_oen[13]
port 434 nsew default input
rlabel metal2 s 48410 0 48466 800 6 la_oen[14]
port 435 nsew default input
rlabel metal2 s 49422 0 49478 800 6 la_oen[15]
port 436 nsew default input
rlabel metal2 s 50342 0 50398 800 6 la_oen[16]
port 437 nsew default input
rlabel metal2 s 51354 0 51410 800 6 la_oen[17]
port 438 nsew default input
rlabel metal2 s 52274 0 52330 800 6 la_oen[18]
port 439 nsew default input
rlabel metal2 s 53286 0 53342 800 6 la_oen[19]
port 440 nsew default input
rlabel metal2 s 35898 0 35954 800 6 la_oen[1]
port 441 nsew default input
rlabel metal2 s 54298 0 54354 800 6 la_oen[20]
port 442 nsew default input
rlabel metal2 s 55218 0 55274 800 6 la_oen[21]
port 443 nsew default input
rlabel metal2 s 56230 0 56286 800 6 la_oen[22]
port 444 nsew default input
rlabel metal2 s 57150 0 57206 800 6 la_oen[23]
port 445 nsew default input
rlabel metal2 s 58162 0 58218 800 6 la_oen[24]
port 446 nsew default input
rlabel metal2 s 59082 0 59138 800 6 la_oen[25]
port 447 nsew default input
rlabel metal2 s 60094 0 60150 800 6 la_oen[26]
port 448 nsew default input
rlabel metal2 s 61014 0 61070 800 6 la_oen[27]
port 449 nsew default input
rlabel metal2 s 62026 0 62082 800 6 la_oen[28]
port 450 nsew default input
rlabel metal2 s 62946 0 63002 800 6 la_oen[29]
port 451 nsew default input
rlabel metal2 s 36818 0 36874 800 6 la_oen[2]
port 452 nsew default input
rlabel metal2 s 63958 0 64014 800 6 la_oen[30]
port 453 nsew default input
rlabel metal2 s 64878 0 64934 800 6 la_oen[31]
port 454 nsew default input
rlabel metal2 s 65890 0 65946 800 6 la_oen[32]
port 455 nsew default input
rlabel metal2 s 66810 0 66866 800 6 la_oen[33]
port 456 nsew default input
rlabel metal2 s 67822 0 67878 800 6 la_oen[34]
port 457 nsew default input
rlabel metal2 s 68742 0 68798 800 6 la_oen[35]
port 458 nsew default input
rlabel metal2 s 69754 0 69810 800 6 la_oen[36]
port 459 nsew default input
rlabel metal2 s 70674 0 70730 800 6 la_oen[37]
port 460 nsew default input
rlabel metal2 s 71686 0 71742 800 6 la_oen[38]
port 461 nsew default input
rlabel metal2 s 72606 0 72662 800 6 la_oen[39]
port 462 nsew default input
rlabel metal2 s 37830 0 37886 800 6 la_oen[3]
port 463 nsew default input
rlabel metal2 s 73618 0 73674 800 6 la_oen[40]
port 464 nsew default input
rlabel metal2 s 74538 0 74594 800 6 la_oen[41]
port 465 nsew default input
rlabel metal2 s 75550 0 75606 800 6 la_oen[42]
port 466 nsew default input
rlabel metal2 s 76470 0 76526 800 6 la_oen[43]
port 467 nsew default input
rlabel metal2 s 77482 0 77538 800 6 la_oen[44]
port 468 nsew default input
rlabel metal2 s 78402 0 78458 800 6 la_oen[45]
port 469 nsew default input
rlabel metal2 s 79414 0 79470 800 6 la_oen[46]
port 470 nsew default input
rlabel metal2 s 80426 0 80482 800 6 la_oen[47]
port 471 nsew default input
rlabel metal2 s 81346 0 81402 800 6 la_oen[48]
port 472 nsew default input
rlabel metal2 s 82358 0 82414 800 6 la_oen[49]
port 473 nsew default input
rlabel metal2 s 38750 0 38806 800 6 la_oen[4]
port 474 nsew default input
rlabel metal2 s 83278 0 83334 800 6 la_oen[50]
port 475 nsew default input
rlabel metal2 s 84290 0 84346 800 6 la_oen[51]
port 476 nsew default input
rlabel metal2 s 85210 0 85266 800 6 la_oen[52]
port 477 nsew default input
rlabel metal2 s 86222 0 86278 800 6 la_oen[53]
port 478 nsew default input
rlabel metal2 s 87142 0 87198 800 6 la_oen[54]
port 479 nsew default input
rlabel metal2 s 88154 0 88210 800 6 la_oen[55]
port 480 nsew default input
rlabel metal2 s 89074 0 89130 800 6 la_oen[56]
port 481 nsew default input
rlabel metal2 s 90086 0 90142 800 6 la_oen[57]
port 482 nsew default input
rlabel metal2 s 91006 0 91062 800 6 la_oen[58]
port 483 nsew default input
rlabel metal2 s 92018 0 92074 800 6 la_oen[59]
port 484 nsew default input
rlabel metal2 s 39762 0 39818 800 6 la_oen[5]
port 485 nsew default input
rlabel metal2 s 92938 0 92994 800 6 la_oen[60]
port 486 nsew default input
rlabel metal2 s 93950 0 94006 800 6 la_oen[61]
port 487 nsew default input
rlabel metal2 s 94870 0 94926 800 6 la_oen[62]
port 488 nsew default input
rlabel metal2 s 95882 0 95938 800 6 la_oen[63]
port 489 nsew default input
rlabel metal2 s 96802 0 96858 800 6 la_oen[64]
port 490 nsew default input
rlabel metal2 s 97814 0 97870 800 6 la_oen[65]
port 491 nsew default input
rlabel metal2 s 98734 0 98790 800 6 la_oen[66]
port 492 nsew default input
rlabel metal2 s 99746 0 99802 800 6 la_oen[67]
port 493 nsew default input
rlabel metal2 s 100666 0 100722 800 6 la_oen[68]
port 494 nsew default input
rlabel metal2 s 101678 0 101734 800 6 la_oen[69]
port 495 nsew default input
rlabel metal2 s 40682 0 40738 800 6 la_oen[6]
port 496 nsew default input
rlabel metal2 s 102598 0 102654 800 6 la_oen[70]
port 497 nsew default input
rlabel metal2 s 103610 0 103666 800 6 la_oen[71]
port 498 nsew default input
rlabel metal2 s 104530 0 104586 800 6 la_oen[72]
port 499 nsew default input
rlabel metal2 s 105542 0 105598 800 6 la_oen[73]
port 500 nsew default input
rlabel metal2 s 106462 0 106518 800 6 la_oen[74]
port 501 nsew default input
rlabel metal2 s 107474 0 107530 800 6 la_oen[75]
port 502 nsew default input
rlabel metal2 s 108486 0 108542 800 6 la_oen[76]
port 503 nsew default input
rlabel metal2 s 109406 0 109462 800 6 la_oen[77]
port 504 nsew default input
rlabel metal2 s 110418 0 110474 800 6 la_oen[78]
port 505 nsew default input
rlabel metal2 s 111338 0 111394 800 6 la_oen[79]
port 506 nsew default input
rlabel metal2 s 41694 0 41750 800 6 la_oen[7]
port 507 nsew default input
rlabel metal2 s 112350 0 112406 800 6 la_oen[80]
port 508 nsew default input
rlabel metal2 s 113270 0 113326 800 6 la_oen[81]
port 509 nsew default input
rlabel metal2 s 114282 0 114338 800 6 la_oen[82]
port 510 nsew default input
rlabel metal2 s 115202 0 115258 800 6 la_oen[83]
port 511 nsew default input
rlabel metal2 s 116214 0 116270 800 6 la_oen[84]
port 512 nsew default input
rlabel metal2 s 117134 0 117190 800 6 la_oen[85]
port 513 nsew default input
rlabel metal2 s 118146 0 118202 800 6 la_oen[86]
port 514 nsew default input
rlabel metal2 s 119066 0 119122 800 6 la_oen[87]
port 515 nsew default input
rlabel metal2 s 120078 0 120134 800 6 la_oen[88]
port 516 nsew default input
rlabel metal2 s 120998 0 121054 800 6 la_oen[89]
port 517 nsew default input
rlabel metal2 s 42614 0 42670 800 6 la_oen[8]
port 518 nsew default input
rlabel metal2 s 122010 0 122066 800 6 la_oen[90]
port 519 nsew default input
rlabel metal2 s 122930 0 122986 800 6 la_oen[91]
port 520 nsew default input
rlabel metal2 s 123942 0 123998 800 6 la_oen[92]
port 521 nsew default input
rlabel metal2 s 124862 0 124918 800 6 la_oen[93]
port 522 nsew default input
rlabel metal2 s 125874 0 125930 800 6 la_oen[94]
port 523 nsew default input
rlabel metal2 s 126794 0 126850 800 6 la_oen[95]
port 524 nsew default input
rlabel metal2 s 127806 0 127862 800 6 la_oen[96]
port 525 nsew default input
rlabel metal2 s 128726 0 128782 800 6 la_oen[97]
port 526 nsew default input
rlabel metal2 s 129738 0 129794 800 6 la_oen[98]
port 527 nsew default input
rlabel metal2 s 130658 0 130714 800 6 la_oen[99]
port 528 nsew default input
rlabel metal2 s 43626 0 43682 800 6 la_oen[9]
port 529 nsew default input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 530 nsew default input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 531 nsew default input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 532 nsew default output
rlabel metal2 s 2042 0 2098 800 6 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 13910 0 13966 800 6 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 20718 0 20774 800 6 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 21638 0 21694 800 6 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 22650 0 22706 800 6 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 26514 0 26570 800 6 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 28446 0 28502 800 6 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 29458 0 29514 800 6 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 4618 0 4674 800 6 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 33322 0 33378 800 6 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 11058 0 11114 800 6 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 1030 0 1086 800 6 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_o[0]
port 598 nsew default output
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_o[10]
port 599 nsew default output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[11]
port 600 nsew default output
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_o[12]
port 601 nsew default output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[13]
port 602 nsew default output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[14]
port 603 nsew default output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[15]
port 604 nsew default output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[16]
port 605 nsew default output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[17]
port 606 nsew default output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[18]
port 607 nsew default output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[19]
port 608 nsew default output
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_o[1]
port 609 nsew default output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[20]
port 610 nsew default output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[21]
port 611 nsew default output
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_o[22]
port 612 nsew default output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[23]
port 613 nsew default output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[24]
port 614 nsew default output
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[25]
port 615 nsew default output
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[26]
port 616 nsew default output
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_o[27]
port 617 nsew default output
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_o[28]
port 618 nsew default output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[29]
port 619 nsew default output
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_o[2]
port 620 nsew default output
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_o[30]
port 621 nsew default output
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_o[31]
port 622 nsew default output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[3]
port 623 nsew default output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[4]
port 624 nsew default output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[5]
port 625 nsew default output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[6]
port 626 nsew default output
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_o[7]
port 627 nsew default output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[8]
port 628 nsew default output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[9]
port 629 nsew default output
rlabel metal2 s 2962 0 3018 800 6 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 4250 0 4306 800 6 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 5538 0 5594 800 6 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 6826 0 6882 800 6 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 1398 0 1454 800 6 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 1674 0 1730 800 6 wbs_we_i
port 635 nsew default input
rlabel metal4 s 4208 2128 4528 157808 6 VPWR
port 636 nsew power input
rlabel metal4 s 19568 2128 19888 157808 6 VGND
port 637 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 160000 160000
string LEFview TRUE
<< end >>
