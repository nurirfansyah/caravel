magic
tech sky130A
magscale 1 2
timestamp 1608359845
<< obsli1 >>
rect 1104 2159 278852 237745
<< obsm1 >>
rect 290 1096 279666 237776
<< metal2 >>
rect 1122 239200 1178 240000
rect 3330 239200 3386 240000
rect 5538 239200 5594 240000
rect 7838 239200 7894 240000
rect 10046 239200 10102 240000
rect 12254 239200 12310 240000
rect 14554 239200 14610 240000
rect 16762 239200 16818 240000
rect 18970 239200 19026 240000
rect 21270 239200 21326 240000
rect 23478 239200 23534 240000
rect 25686 239200 25742 240000
rect 27986 239200 28042 240000
rect 30194 239200 30250 240000
rect 32402 239200 32458 240000
rect 34702 239200 34758 240000
rect 36910 239200 36966 240000
rect 39118 239200 39174 240000
rect 41418 239200 41474 240000
rect 43626 239200 43682 240000
rect 45834 239200 45890 240000
rect 48134 239200 48190 240000
rect 50342 239200 50398 240000
rect 52550 239200 52606 240000
rect 54850 239200 54906 240000
rect 57058 239200 57114 240000
rect 59266 239200 59322 240000
rect 61566 239200 61622 240000
rect 63774 239200 63830 240000
rect 65982 239200 66038 240000
rect 68282 239200 68338 240000
rect 70490 239200 70546 240000
rect 72790 239200 72846 240000
rect 74998 239200 75054 240000
rect 77206 239200 77262 240000
rect 79506 239200 79562 240000
rect 81714 239200 81770 240000
rect 83922 239200 83978 240000
rect 86222 239200 86278 240000
rect 88430 239200 88486 240000
rect 90638 239200 90694 240000
rect 92938 239200 92994 240000
rect 95146 239200 95202 240000
rect 97354 239200 97410 240000
rect 99654 239200 99710 240000
rect 101862 239200 101918 240000
rect 104070 239200 104126 240000
rect 106370 239200 106426 240000
rect 108578 239200 108634 240000
rect 110786 239200 110842 240000
rect 113086 239200 113142 240000
rect 115294 239200 115350 240000
rect 117502 239200 117558 240000
rect 119802 239200 119858 240000
rect 122010 239200 122066 240000
rect 124218 239200 124274 240000
rect 126518 239200 126574 240000
rect 128726 239200 128782 240000
rect 130934 239200 130990 240000
rect 133234 239200 133290 240000
rect 135442 239200 135498 240000
rect 137650 239200 137706 240000
rect 139950 239200 140006 240000
rect 142158 239200 142214 240000
rect 144458 239200 144514 240000
rect 146666 239200 146722 240000
rect 148874 239200 148930 240000
rect 151174 239200 151230 240000
rect 153382 239200 153438 240000
rect 155590 239200 155646 240000
rect 157890 239200 157946 240000
rect 160098 239200 160154 240000
rect 162306 239200 162362 240000
rect 164606 239200 164662 240000
rect 166814 239200 166870 240000
rect 169022 239200 169078 240000
rect 171322 239200 171378 240000
rect 173530 239200 173586 240000
rect 175738 239200 175794 240000
rect 178038 239200 178094 240000
rect 180246 239200 180302 240000
rect 182454 239200 182510 240000
rect 184754 239200 184810 240000
rect 186962 239200 187018 240000
rect 189170 239200 189226 240000
rect 191470 239200 191526 240000
rect 193678 239200 193734 240000
rect 195886 239200 195942 240000
rect 198186 239200 198242 240000
rect 200394 239200 200450 240000
rect 202602 239200 202658 240000
rect 204902 239200 204958 240000
rect 207110 239200 207166 240000
rect 209318 239200 209374 240000
rect 211618 239200 211674 240000
rect 213826 239200 213882 240000
rect 216126 239200 216182 240000
rect 218334 239200 218390 240000
rect 220542 239200 220598 240000
rect 222842 239200 222898 240000
rect 225050 239200 225106 240000
rect 227258 239200 227314 240000
rect 229558 239200 229614 240000
rect 231766 239200 231822 240000
rect 233974 239200 234030 240000
rect 236274 239200 236330 240000
rect 238482 239200 238538 240000
rect 240690 239200 240746 240000
rect 242990 239200 243046 240000
rect 245198 239200 245254 240000
rect 247406 239200 247462 240000
rect 249706 239200 249762 240000
rect 251914 239200 251970 240000
rect 254122 239200 254178 240000
rect 256422 239200 256478 240000
rect 258630 239200 258686 240000
rect 260838 239200 260894 240000
rect 263138 239200 263194 240000
rect 265346 239200 265402 240000
rect 267554 239200 267610 240000
rect 269854 239200 269910 240000
rect 272062 239200 272118 240000
rect 274270 239200 274326 240000
rect 276570 239200 276626 240000
rect 278778 239200 278834 240000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9862 0 9918 800
rect 10414 0 10470 800
rect 10966 0 11022 800
rect 11518 0 11574 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13726 0 13782 800
rect 14370 0 14426 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 16026 0 16082 800
rect 16578 0 16634 800
rect 17130 0 17186 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18878 0 18934 800
rect 19430 0 19486 800
rect 19982 0 20038 800
rect 20534 0 20590 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22190 0 22246 800
rect 22742 0 22798 800
rect 23386 0 23442 800
rect 23938 0 23994 800
rect 24490 0 24546 800
rect 25042 0 25098 800
rect 25594 0 25650 800
rect 26146 0 26202 800
rect 26698 0 26754 800
rect 27250 0 27306 800
rect 27894 0 27950 800
rect 28446 0 28502 800
rect 28998 0 29054 800
rect 29550 0 29606 800
rect 30102 0 30158 800
rect 30654 0 30710 800
rect 31206 0 31262 800
rect 31758 0 31814 800
rect 32310 0 32366 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34058 0 34114 800
rect 34610 0 34666 800
rect 35162 0 35218 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37462 0 37518 800
rect 38014 0 38070 800
rect 38566 0 38622 800
rect 39118 0 39174 800
rect 39670 0 39726 800
rect 40222 0 40278 800
rect 40774 0 40830 800
rect 41326 0 41382 800
rect 41970 0 42026 800
rect 42522 0 42578 800
rect 43074 0 43130 800
rect 43626 0 43682 800
rect 44178 0 44234 800
rect 44730 0 44786 800
rect 45282 0 45338 800
rect 45834 0 45890 800
rect 46478 0 46534 800
rect 47030 0 47086 800
rect 47582 0 47638 800
rect 48134 0 48190 800
rect 48686 0 48742 800
rect 49238 0 49294 800
rect 49790 0 49846 800
rect 50342 0 50398 800
rect 50986 0 51042 800
rect 51538 0 51594 800
rect 52090 0 52146 800
rect 52642 0 52698 800
rect 53194 0 53250 800
rect 53746 0 53802 800
rect 54298 0 54354 800
rect 54850 0 54906 800
rect 55494 0 55550 800
rect 56046 0 56102 800
rect 56598 0 56654 800
rect 57150 0 57206 800
rect 57702 0 57758 800
rect 58254 0 58310 800
rect 58806 0 58862 800
rect 59358 0 59414 800
rect 60002 0 60058 800
rect 60554 0 60610 800
rect 61106 0 61162 800
rect 61658 0 61714 800
rect 62210 0 62266 800
rect 62762 0 62818 800
rect 63314 0 63370 800
rect 63866 0 63922 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65614 0 65670 800
rect 66166 0 66222 800
rect 66718 0 66774 800
rect 67270 0 67326 800
rect 67822 0 67878 800
rect 68374 0 68430 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70122 0 70178 800
rect 70674 0 70730 800
rect 71226 0 71282 800
rect 71778 0 71834 800
rect 72330 0 72386 800
rect 72882 0 72938 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74630 0 74686 800
rect 75182 0 75238 800
rect 75734 0 75790 800
rect 76286 0 76342 800
rect 76838 0 76894 800
rect 77390 0 77446 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79138 0 79194 800
rect 79690 0 79746 800
rect 80242 0 80298 800
rect 80794 0 80850 800
rect 81346 0 81402 800
rect 81898 0 81954 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 83646 0 83702 800
rect 84198 0 84254 800
rect 84750 0 84806 800
rect 85302 0 85358 800
rect 85854 0 85910 800
rect 86406 0 86462 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88154 0 88210 800
rect 88706 0 88762 800
rect 89258 0 89314 800
rect 89810 0 89866 800
rect 90362 0 90418 800
rect 90914 0 90970 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 92662 0 92718 800
rect 93214 0 93270 800
rect 93766 0 93822 800
rect 94318 0 94374 800
rect 94870 0 94926 800
rect 95422 0 95478 800
rect 95974 0 96030 800
rect 96526 0 96582 800
rect 97170 0 97226 800
rect 97722 0 97778 800
rect 98274 0 98330 800
rect 98826 0 98882 800
rect 99378 0 99434 800
rect 99930 0 99986 800
rect 100482 0 100538 800
rect 101034 0 101090 800
rect 101678 0 101734 800
rect 102230 0 102286 800
rect 102782 0 102838 800
rect 103334 0 103390 800
rect 103886 0 103942 800
rect 104438 0 104494 800
rect 104990 0 105046 800
rect 105542 0 105598 800
rect 106186 0 106242 800
rect 106738 0 106794 800
rect 107290 0 107346 800
rect 107842 0 107898 800
rect 108394 0 108450 800
rect 108946 0 109002 800
rect 109498 0 109554 800
rect 110050 0 110106 800
rect 110694 0 110750 800
rect 111246 0 111302 800
rect 111798 0 111854 800
rect 112350 0 112406 800
rect 112902 0 112958 800
rect 113454 0 113510 800
rect 114006 0 114062 800
rect 114558 0 114614 800
rect 115202 0 115258 800
rect 115754 0 115810 800
rect 116306 0 116362 800
rect 116858 0 116914 800
rect 117410 0 117466 800
rect 117962 0 118018 800
rect 118514 0 118570 800
rect 119066 0 119122 800
rect 119710 0 119766 800
rect 120262 0 120318 800
rect 120814 0 120870 800
rect 121366 0 121422 800
rect 121918 0 121974 800
rect 122470 0 122526 800
rect 123022 0 123078 800
rect 123574 0 123630 800
rect 124218 0 124274 800
rect 124770 0 124826 800
rect 125322 0 125378 800
rect 125874 0 125930 800
rect 126426 0 126482 800
rect 126978 0 127034 800
rect 127530 0 127586 800
rect 128082 0 128138 800
rect 128634 0 128690 800
rect 129278 0 129334 800
rect 129830 0 129886 800
rect 130382 0 130438 800
rect 130934 0 130990 800
rect 131486 0 131542 800
rect 132038 0 132094 800
rect 132590 0 132646 800
rect 133142 0 133198 800
rect 133786 0 133842 800
rect 134338 0 134394 800
rect 134890 0 134946 800
rect 135442 0 135498 800
rect 135994 0 136050 800
rect 136546 0 136602 800
rect 137098 0 137154 800
rect 137650 0 137706 800
rect 138294 0 138350 800
rect 138846 0 138902 800
rect 139398 0 139454 800
rect 139950 0 140006 800
rect 140502 0 140558 800
rect 141054 0 141110 800
rect 141606 0 141662 800
rect 142158 0 142214 800
rect 142802 0 142858 800
rect 143354 0 143410 800
rect 143906 0 143962 800
rect 144458 0 144514 800
rect 145010 0 145066 800
rect 145562 0 145618 800
rect 146114 0 146170 800
rect 146666 0 146722 800
rect 147310 0 147366 800
rect 147862 0 147918 800
rect 148414 0 148470 800
rect 148966 0 149022 800
rect 149518 0 149574 800
rect 150070 0 150126 800
rect 150622 0 150678 800
rect 151174 0 151230 800
rect 151818 0 151874 800
rect 152370 0 152426 800
rect 152922 0 152978 800
rect 153474 0 153530 800
rect 154026 0 154082 800
rect 154578 0 154634 800
rect 155130 0 155186 800
rect 155682 0 155738 800
rect 156234 0 156290 800
rect 156878 0 156934 800
rect 157430 0 157486 800
rect 157982 0 158038 800
rect 158534 0 158590 800
rect 159086 0 159142 800
rect 159638 0 159694 800
rect 160190 0 160246 800
rect 160742 0 160798 800
rect 161386 0 161442 800
rect 161938 0 161994 800
rect 162490 0 162546 800
rect 163042 0 163098 800
rect 163594 0 163650 800
rect 164146 0 164202 800
rect 164698 0 164754 800
rect 165250 0 165306 800
rect 165894 0 165950 800
rect 166446 0 166502 800
rect 166998 0 167054 800
rect 167550 0 167606 800
rect 168102 0 168158 800
rect 168654 0 168710 800
rect 169206 0 169262 800
rect 169758 0 169814 800
rect 170402 0 170458 800
rect 170954 0 171010 800
rect 171506 0 171562 800
rect 172058 0 172114 800
rect 172610 0 172666 800
rect 173162 0 173218 800
rect 173714 0 173770 800
rect 174266 0 174322 800
rect 174910 0 174966 800
rect 175462 0 175518 800
rect 176014 0 176070 800
rect 176566 0 176622 800
rect 177118 0 177174 800
rect 177670 0 177726 800
rect 178222 0 178278 800
rect 178774 0 178830 800
rect 179418 0 179474 800
rect 179970 0 180026 800
rect 180522 0 180578 800
rect 181074 0 181130 800
rect 181626 0 181682 800
rect 182178 0 182234 800
rect 182730 0 182786 800
rect 183282 0 183338 800
rect 183926 0 183982 800
rect 184478 0 184534 800
rect 185030 0 185086 800
rect 185582 0 185638 800
rect 186134 0 186190 800
rect 186686 0 186742 800
rect 187238 0 187294 800
rect 187790 0 187846 800
rect 188342 0 188398 800
rect 188986 0 189042 800
rect 189538 0 189594 800
rect 190090 0 190146 800
rect 190642 0 190698 800
rect 191194 0 191250 800
rect 191746 0 191802 800
rect 192298 0 192354 800
rect 192850 0 192906 800
rect 193494 0 193550 800
rect 194046 0 194102 800
rect 194598 0 194654 800
rect 195150 0 195206 800
rect 195702 0 195758 800
rect 196254 0 196310 800
rect 196806 0 196862 800
rect 197358 0 197414 800
rect 198002 0 198058 800
rect 198554 0 198610 800
rect 199106 0 199162 800
rect 199658 0 199714 800
rect 200210 0 200266 800
rect 200762 0 200818 800
rect 201314 0 201370 800
rect 201866 0 201922 800
rect 202510 0 202566 800
rect 203062 0 203118 800
rect 203614 0 203670 800
rect 204166 0 204222 800
rect 204718 0 204774 800
rect 205270 0 205326 800
rect 205822 0 205878 800
rect 206374 0 206430 800
rect 207018 0 207074 800
rect 207570 0 207626 800
rect 208122 0 208178 800
rect 208674 0 208730 800
rect 209226 0 209282 800
rect 209778 0 209834 800
rect 210330 0 210386 800
rect 210882 0 210938 800
rect 211526 0 211582 800
rect 212078 0 212134 800
rect 212630 0 212686 800
rect 213182 0 213238 800
rect 213734 0 213790 800
rect 214286 0 214342 800
rect 214838 0 214894 800
rect 215390 0 215446 800
rect 216034 0 216090 800
rect 216586 0 216642 800
rect 217138 0 217194 800
rect 217690 0 217746 800
rect 218242 0 218298 800
rect 218794 0 218850 800
rect 219346 0 219402 800
rect 219898 0 219954 800
rect 220450 0 220506 800
rect 221094 0 221150 800
rect 221646 0 221702 800
rect 222198 0 222254 800
rect 222750 0 222806 800
rect 223302 0 223358 800
rect 223854 0 223910 800
rect 224406 0 224462 800
rect 224958 0 225014 800
rect 225602 0 225658 800
rect 226154 0 226210 800
rect 226706 0 226762 800
rect 227258 0 227314 800
rect 227810 0 227866 800
rect 228362 0 228418 800
rect 228914 0 228970 800
rect 229466 0 229522 800
rect 230110 0 230166 800
rect 230662 0 230718 800
rect 231214 0 231270 800
rect 231766 0 231822 800
rect 232318 0 232374 800
rect 232870 0 232926 800
rect 233422 0 233478 800
rect 233974 0 234030 800
rect 234618 0 234674 800
rect 235170 0 235226 800
rect 235722 0 235778 800
rect 236274 0 236330 800
rect 236826 0 236882 800
rect 237378 0 237434 800
rect 237930 0 237986 800
rect 238482 0 238538 800
rect 239126 0 239182 800
rect 239678 0 239734 800
rect 240230 0 240286 800
rect 240782 0 240838 800
rect 241334 0 241390 800
rect 241886 0 241942 800
rect 242438 0 242494 800
rect 242990 0 243046 800
rect 243634 0 243690 800
rect 244186 0 244242 800
rect 244738 0 244794 800
rect 245290 0 245346 800
rect 245842 0 245898 800
rect 246394 0 246450 800
rect 246946 0 247002 800
rect 247498 0 247554 800
rect 248142 0 248198 800
rect 248694 0 248750 800
rect 249246 0 249302 800
rect 249798 0 249854 800
rect 250350 0 250406 800
rect 250902 0 250958 800
rect 251454 0 251510 800
rect 252006 0 252062 800
rect 252558 0 252614 800
rect 253202 0 253258 800
rect 253754 0 253810 800
rect 254306 0 254362 800
rect 254858 0 254914 800
rect 255410 0 255466 800
rect 255962 0 256018 800
rect 256514 0 256570 800
rect 257066 0 257122 800
rect 257710 0 257766 800
rect 258262 0 258318 800
rect 258814 0 258870 800
rect 259366 0 259422 800
rect 259918 0 259974 800
rect 260470 0 260526 800
rect 261022 0 261078 800
rect 261574 0 261630 800
rect 262218 0 262274 800
rect 262770 0 262826 800
rect 263322 0 263378 800
rect 263874 0 263930 800
rect 264426 0 264482 800
rect 264978 0 265034 800
rect 265530 0 265586 800
rect 266082 0 266138 800
rect 266726 0 266782 800
rect 267278 0 267334 800
rect 267830 0 267886 800
rect 268382 0 268438 800
rect 268934 0 268990 800
rect 269486 0 269542 800
rect 270038 0 270094 800
rect 270590 0 270646 800
rect 271234 0 271290 800
rect 271786 0 271842 800
rect 272338 0 272394 800
rect 272890 0 272946 800
rect 273442 0 273498 800
rect 273994 0 274050 800
rect 274546 0 274602 800
rect 275098 0 275154 800
rect 275742 0 275798 800
rect 276294 0 276350 800
rect 276846 0 276902 800
rect 277398 0 277454 800
rect 277950 0 278006 800
rect 278502 0 278558 800
rect 279054 0 279110 800
rect 279606 0 279662 800
<< obsm2 >>
rect 296 239144 1066 239200
rect 1234 239144 3274 239200
rect 3442 239144 5482 239200
rect 5650 239144 7782 239200
rect 7950 239144 9990 239200
rect 10158 239144 12198 239200
rect 12366 239144 14498 239200
rect 14666 239144 16706 239200
rect 16874 239144 18914 239200
rect 19082 239144 21214 239200
rect 21382 239144 23422 239200
rect 23590 239144 25630 239200
rect 25798 239144 27930 239200
rect 28098 239144 30138 239200
rect 30306 239144 32346 239200
rect 32514 239144 34646 239200
rect 34814 239144 36854 239200
rect 37022 239144 39062 239200
rect 39230 239144 41362 239200
rect 41530 239144 43570 239200
rect 43738 239144 45778 239200
rect 45946 239144 48078 239200
rect 48246 239144 50286 239200
rect 50454 239144 52494 239200
rect 52662 239144 54794 239200
rect 54962 239144 57002 239200
rect 57170 239144 59210 239200
rect 59378 239144 61510 239200
rect 61678 239144 63718 239200
rect 63886 239144 65926 239200
rect 66094 239144 68226 239200
rect 68394 239144 70434 239200
rect 70602 239144 72734 239200
rect 72902 239144 74942 239200
rect 75110 239144 77150 239200
rect 77318 239144 79450 239200
rect 79618 239144 81658 239200
rect 81826 239144 83866 239200
rect 84034 239144 86166 239200
rect 86334 239144 88374 239200
rect 88542 239144 90582 239200
rect 90750 239144 92882 239200
rect 93050 239144 95090 239200
rect 95258 239144 97298 239200
rect 97466 239144 99598 239200
rect 99766 239144 101806 239200
rect 101974 239144 104014 239200
rect 104182 239144 106314 239200
rect 106482 239144 108522 239200
rect 108690 239144 110730 239200
rect 110898 239144 113030 239200
rect 113198 239144 115238 239200
rect 115406 239144 117446 239200
rect 117614 239144 119746 239200
rect 119914 239144 121954 239200
rect 122122 239144 124162 239200
rect 124330 239144 126462 239200
rect 126630 239144 128670 239200
rect 128838 239144 130878 239200
rect 131046 239144 133178 239200
rect 133346 239144 135386 239200
rect 135554 239144 137594 239200
rect 137762 239144 139894 239200
rect 140062 239144 142102 239200
rect 142270 239144 144402 239200
rect 144570 239144 146610 239200
rect 146778 239144 148818 239200
rect 148986 239144 151118 239200
rect 151286 239144 153326 239200
rect 153494 239144 155534 239200
rect 155702 239144 157834 239200
rect 158002 239144 160042 239200
rect 160210 239144 162250 239200
rect 162418 239144 164550 239200
rect 164718 239144 166758 239200
rect 166926 239144 168966 239200
rect 169134 239144 171266 239200
rect 171434 239144 173474 239200
rect 173642 239144 175682 239200
rect 175850 239144 177982 239200
rect 178150 239144 180190 239200
rect 180358 239144 182398 239200
rect 182566 239144 184698 239200
rect 184866 239144 186906 239200
rect 187074 239144 189114 239200
rect 189282 239144 191414 239200
rect 191582 239144 193622 239200
rect 193790 239144 195830 239200
rect 195998 239144 198130 239200
rect 198298 239144 200338 239200
rect 200506 239144 202546 239200
rect 202714 239144 204846 239200
rect 205014 239144 207054 239200
rect 207222 239144 209262 239200
rect 209430 239144 211562 239200
rect 211730 239144 213770 239200
rect 213938 239144 216070 239200
rect 216238 239144 218278 239200
rect 218446 239144 220486 239200
rect 220654 239144 222786 239200
rect 222954 239144 224994 239200
rect 225162 239144 227202 239200
rect 227370 239144 229502 239200
rect 229670 239144 231710 239200
rect 231878 239144 233918 239200
rect 234086 239144 236218 239200
rect 236386 239144 238426 239200
rect 238594 239144 240634 239200
rect 240802 239144 242934 239200
rect 243102 239144 245142 239200
rect 245310 239144 247350 239200
rect 247518 239144 249650 239200
rect 249818 239144 251858 239200
rect 252026 239144 254066 239200
rect 254234 239144 256366 239200
rect 256534 239144 258574 239200
rect 258742 239144 260782 239200
rect 260950 239144 263082 239200
rect 263250 239144 265290 239200
rect 265458 239144 267498 239200
rect 267666 239144 269798 239200
rect 269966 239144 272006 239200
rect 272174 239144 274214 239200
rect 274382 239144 276514 239200
rect 276682 239144 278722 239200
rect 278890 239144 279660 239200
rect 296 856 279660 239144
rect 406 800 790 856
rect 958 800 1342 856
rect 1510 800 1894 856
rect 2062 800 2446 856
rect 2614 800 2998 856
rect 3166 800 3550 856
rect 3718 800 4102 856
rect 4270 800 4654 856
rect 4822 800 5298 856
rect 5466 800 5850 856
rect 6018 800 6402 856
rect 6570 800 6954 856
rect 7122 800 7506 856
rect 7674 800 8058 856
rect 8226 800 8610 856
rect 8778 800 9162 856
rect 9330 800 9806 856
rect 9974 800 10358 856
rect 10526 800 10910 856
rect 11078 800 11462 856
rect 11630 800 12014 856
rect 12182 800 12566 856
rect 12734 800 13118 856
rect 13286 800 13670 856
rect 13838 800 14314 856
rect 14482 800 14866 856
rect 15034 800 15418 856
rect 15586 800 15970 856
rect 16138 800 16522 856
rect 16690 800 17074 856
rect 17242 800 17626 856
rect 17794 800 18178 856
rect 18346 800 18822 856
rect 18990 800 19374 856
rect 19542 800 19926 856
rect 20094 800 20478 856
rect 20646 800 21030 856
rect 21198 800 21582 856
rect 21750 800 22134 856
rect 22302 800 22686 856
rect 22854 800 23330 856
rect 23498 800 23882 856
rect 24050 800 24434 856
rect 24602 800 24986 856
rect 25154 800 25538 856
rect 25706 800 26090 856
rect 26258 800 26642 856
rect 26810 800 27194 856
rect 27362 800 27838 856
rect 28006 800 28390 856
rect 28558 800 28942 856
rect 29110 800 29494 856
rect 29662 800 30046 856
rect 30214 800 30598 856
rect 30766 800 31150 856
rect 31318 800 31702 856
rect 31870 800 32254 856
rect 32422 800 32898 856
rect 33066 800 33450 856
rect 33618 800 34002 856
rect 34170 800 34554 856
rect 34722 800 35106 856
rect 35274 800 35658 856
rect 35826 800 36210 856
rect 36378 800 36762 856
rect 36930 800 37406 856
rect 37574 800 37958 856
rect 38126 800 38510 856
rect 38678 800 39062 856
rect 39230 800 39614 856
rect 39782 800 40166 856
rect 40334 800 40718 856
rect 40886 800 41270 856
rect 41438 800 41914 856
rect 42082 800 42466 856
rect 42634 800 43018 856
rect 43186 800 43570 856
rect 43738 800 44122 856
rect 44290 800 44674 856
rect 44842 800 45226 856
rect 45394 800 45778 856
rect 45946 800 46422 856
rect 46590 800 46974 856
rect 47142 800 47526 856
rect 47694 800 48078 856
rect 48246 800 48630 856
rect 48798 800 49182 856
rect 49350 800 49734 856
rect 49902 800 50286 856
rect 50454 800 50930 856
rect 51098 800 51482 856
rect 51650 800 52034 856
rect 52202 800 52586 856
rect 52754 800 53138 856
rect 53306 800 53690 856
rect 53858 800 54242 856
rect 54410 800 54794 856
rect 54962 800 55438 856
rect 55606 800 55990 856
rect 56158 800 56542 856
rect 56710 800 57094 856
rect 57262 800 57646 856
rect 57814 800 58198 856
rect 58366 800 58750 856
rect 58918 800 59302 856
rect 59470 800 59946 856
rect 60114 800 60498 856
rect 60666 800 61050 856
rect 61218 800 61602 856
rect 61770 800 62154 856
rect 62322 800 62706 856
rect 62874 800 63258 856
rect 63426 800 63810 856
rect 63978 800 64362 856
rect 64530 800 65006 856
rect 65174 800 65558 856
rect 65726 800 66110 856
rect 66278 800 66662 856
rect 66830 800 67214 856
rect 67382 800 67766 856
rect 67934 800 68318 856
rect 68486 800 68870 856
rect 69038 800 69514 856
rect 69682 800 70066 856
rect 70234 800 70618 856
rect 70786 800 71170 856
rect 71338 800 71722 856
rect 71890 800 72274 856
rect 72442 800 72826 856
rect 72994 800 73378 856
rect 73546 800 74022 856
rect 74190 800 74574 856
rect 74742 800 75126 856
rect 75294 800 75678 856
rect 75846 800 76230 856
rect 76398 800 76782 856
rect 76950 800 77334 856
rect 77502 800 77886 856
rect 78054 800 78530 856
rect 78698 800 79082 856
rect 79250 800 79634 856
rect 79802 800 80186 856
rect 80354 800 80738 856
rect 80906 800 81290 856
rect 81458 800 81842 856
rect 82010 800 82394 856
rect 82562 800 83038 856
rect 83206 800 83590 856
rect 83758 800 84142 856
rect 84310 800 84694 856
rect 84862 800 85246 856
rect 85414 800 85798 856
rect 85966 800 86350 856
rect 86518 800 86902 856
rect 87070 800 87546 856
rect 87714 800 88098 856
rect 88266 800 88650 856
rect 88818 800 89202 856
rect 89370 800 89754 856
rect 89922 800 90306 856
rect 90474 800 90858 856
rect 91026 800 91410 856
rect 91578 800 92054 856
rect 92222 800 92606 856
rect 92774 800 93158 856
rect 93326 800 93710 856
rect 93878 800 94262 856
rect 94430 800 94814 856
rect 94982 800 95366 856
rect 95534 800 95918 856
rect 96086 800 96470 856
rect 96638 800 97114 856
rect 97282 800 97666 856
rect 97834 800 98218 856
rect 98386 800 98770 856
rect 98938 800 99322 856
rect 99490 800 99874 856
rect 100042 800 100426 856
rect 100594 800 100978 856
rect 101146 800 101622 856
rect 101790 800 102174 856
rect 102342 800 102726 856
rect 102894 800 103278 856
rect 103446 800 103830 856
rect 103998 800 104382 856
rect 104550 800 104934 856
rect 105102 800 105486 856
rect 105654 800 106130 856
rect 106298 800 106682 856
rect 106850 800 107234 856
rect 107402 800 107786 856
rect 107954 800 108338 856
rect 108506 800 108890 856
rect 109058 800 109442 856
rect 109610 800 109994 856
rect 110162 800 110638 856
rect 110806 800 111190 856
rect 111358 800 111742 856
rect 111910 800 112294 856
rect 112462 800 112846 856
rect 113014 800 113398 856
rect 113566 800 113950 856
rect 114118 800 114502 856
rect 114670 800 115146 856
rect 115314 800 115698 856
rect 115866 800 116250 856
rect 116418 800 116802 856
rect 116970 800 117354 856
rect 117522 800 117906 856
rect 118074 800 118458 856
rect 118626 800 119010 856
rect 119178 800 119654 856
rect 119822 800 120206 856
rect 120374 800 120758 856
rect 120926 800 121310 856
rect 121478 800 121862 856
rect 122030 800 122414 856
rect 122582 800 122966 856
rect 123134 800 123518 856
rect 123686 800 124162 856
rect 124330 800 124714 856
rect 124882 800 125266 856
rect 125434 800 125818 856
rect 125986 800 126370 856
rect 126538 800 126922 856
rect 127090 800 127474 856
rect 127642 800 128026 856
rect 128194 800 128578 856
rect 128746 800 129222 856
rect 129390 800 129774 856
rect 129942 800 130326 856
rect 130494 800 130878 856
rect 131046 800 131430 856
rect 131598 800 131982 856
rect 132150 800 132534 856
rect 132702 800 133086 856
rect 133254 800 133730 856
rect 133898 800 134282 856
rect 134450 800 134834 856
rect 135002 800 135386 856
rect 135554 800 135938 856
rect 136106 800 136490 856
rect 136658 800 137042 856
rect 137210 800 137594 856
rect 137762 800 138238 856
rect 138406 800 138790 856
rect 138958 800 139342 856
rect 139510 800 139894 856
rect 140062 800 140446 856
rect 140614 800 140998 856
rect 141166 800 141550 856
rect 141718 800 142102 856
rect 142270 800 142746 856
rect 142914 800 143298 856
rect 143466 800 143850 856
rect 144018 800 144402 856
rect 144570 800 144954 856
rect 145122 800 145506 856
rect 145674 800 146058 856
rect 146226 800 146610 856
rect 146778 800 147254 856
rect 147422 800 147806 856
rect 147974 800 148358 856
rect 148526 800 148910 856
rect 149078 800 149462 856
rect 149630 800 150014 856
rect 150182 800 150566 856
rect 150734 800 151118 856
rect 151286 800 151762 856
rect 151930 800 152314 856
rect 152482 800 152866 856
rect 153034 800 153418 856
rect 153586 800 153970 856
rect 154138 800 154522 856
rect 154690 800 155074 856
rect 155242 800 155626 856
rect 155794 800 156178 856
rect 156346 800 156822 856
rect 156990 800 157374 856
rect 157542 800 157926 856
rect 158094 800 158478 856
rect 158646 800 159030 856
rect 159198 800 159582 856
rect 159750 800 160134 856
rect 160302 800 160686 856
rect 160854 800 161330 856
rect 161498 800 161882 856
rect 162050 800 162434 856
rect 162602 800 162986 856
rect 163154 800 163538 856
rect 163706 800 164090 856
rect 164258 800 164642 856
rect 164810 800 165194 856
rect 165362 800 165838 856
rect 166006 800 166390 856
rect 166558 800 166942 856
rect 167110 800 167494 856
rect 167662 800 168046 856
rect 168214 800 168598 856
rect 168766 800 169150 856
rect 169318 800 169702 856
rect 169870 800 170346 856
rect 170514 800 170898 856
rect 171066 800 171450 856
rect 171618 800 172002 856
rect 172170 800 172554 856
rect 172722 800 173106 856
rect 173274 800 173658 856
rect 173826 800 174210 856
rect 174378 800 174854 856
rect 175022 800 175406 856
rect 175574 800 175958 856
rect 176126 800 176510 856
rect 176678 800 177062 856
rect 177230 800 177614 856
rect 177782 800 178166 856
rect 178334 800 178718 856
rect 178886 800 179362 856
rect 179530 800 179914 856
rect 180082 800 180466 856
rect 180634 800 181018 856
rect 181186 800 181570 856
rect 181738 800 182122 856
rect 182290 800 182674 856
rect 182842 800 183226 856
rect 183394 800 183870 856
rect 184038 800 184422 856
rect 184590 800 184974 856
rect 185142 800 185526 856
rect 185694 800 186078 856
rect 186246 800 186630 856
rect 186798 800 187182 856
rect 187350 800 187734 856
rect 187902 800 188286 856
rect 188454 800 188930 856
rect 189098 800 189482 856
rect 189650 800 190034 856
rect 190202 800 190586 856
rect 190754 800 191138 856
rect 191306 800 191690 856
rect 191858 800 192242 856
rect 192410 800 192794 856
rect 192962 800 193438 856
rect 193606 800 193990 856
rect 194158 800 194542 856
rect 194710 800 195094 856
rect 195262 800 195646 856
rect 195814 800 196198 856
rect 196366 800 196750 856
rect 196918 800 197302 856
rect 197470 800 197946 856
rect 198114 800 198498 856
rect 198666 800 199050 856
rect 199218 800 199602 856
rect 199770 800 200154 856
rect 200322 800 200706 856
rect 200874 800 201258 856
rect 201426 800 201810 856
rect 201978 800 202454 856
rect 202622 800 203006 856
rect 203174 800 203558 856
rect 203726 800 204110 856
rect 204278 800 204662 856
rect 204830 800 205214 856
rect 205382 800 205766 856
rect 205934 800 206318 856
rect 206486 800 206962 856
rect 207130 800 207514 856
rect 207682 800 208066 856
rect 208234 800 208618 856
rect 208786 800 209170 856
rect 209338 800 209722 856
rect 209890 800 210274 856
rect 210442 800 210826 856
rect 210994 800 211470 856
rect 211638 800 212022 856
rect 212190 800 212574 856
rect 212742 800 213126 856
rect 213294 800 213678 856
rect 213846 800 214230 856
rect 214398 800 214782 856
rect 214950 800 215334 856
rect 215502 800 215978 856
rect 216146 800 216530 856
rect 216698 800 217082 856
rect 217250 800 217634 856
rect 217802 800 218186 856
rect 218354 800 218738 856
rect 218906 800 219290 856
rect 219458 800 219842 856
rect 220010 800 220394 856
rect 220562 800 221038 856
rect 221206 800 221590 856
rect 221758 800 222142 856
rect 222310 800 222694 856
rect 222862 800 223246 856
rect 223414 800 223798 856
rect 223966 800 224350 856
rect 224518 800 224902 856
rect 225070 800 225546 856
rect 225714 800 226098 856
rect 226266 800 226650 856
rect 226818 800 227202 856
rect 227370 800 227754 856
rect 227922 800 228306 856
rect 228474 800 228858 856
rect 229026 800 229410 856
rect 229578 800 230054 856
rect 230222 800 230606 856
rect 230774 800 231158 856
rect 231326 800 231710 856
rect 231878 800 232262 856
rect 232430 800 232814 856
rect 232982 800 233366 856
rect 233534 800 233918 856
rect 234086 800 234562 856
rect 234730 800 235114 856
rect 235282 800 235666 856
rect 235834 800 236218 856
rect 236386 800 236770 856
rect 236938 800 237322 856
rect 237490 800 237874 856
rect 238042 800 238426 856
rect 238594 800 239070 856
rect 239238 800 239622 856
rect 239790 800 240174 856
rect 240342 800 240726 856
rect 240894 800 241278 856
rect 241446 800 241830 856
rect 241998 800 242382 856
rect 242550 800 242934 856
rect 243102 800 243578 856
rect 243746 800 244130 856
rect 244298 800 244682 856
rect 244850 800 245234 856
rect 245402 800 245786 856
rect 245954 800 246338 856
rect 246506 800 246890 856
rect 247058 800 247442 856
rect 247610 800 248086 856
rect 248254 800 248638 856
rect 248806 800 249190 856
rect 249358 800 249742 856
rect 249910 800 250294 856
rect 250462 800 250846 856
rect 251014 800 251398 856
rect 251566 800 251950 856
rect 252118 800 252502 856
rect 252670 800 253146 856
rect 253314 800 253698 856
rect 253866 800 254250 856
rect 254418 800 254802 856
rect 254970 800 255354 856
rect 255522 800 255906 856
rect 256074 800 256458 856
rect 256626 800 257010 856
rect 257178 800 257654 856
rect 257822 800 258206 856
rect 258374 800 258758 856
rect 258926 800 259310 856
rect 259478 800 259862 856
rect 260030 800 260414 856
rect 260582 800 260966 856
rect 261134 800 261518 856
rect 261686 800 262162 856
rect 262330 800 262714 856
rect 262882 800 263266 856
rect 263434 800 263818 856
rect 263986 800 264370 856
rect 264538 800 264922 856
rect 265090 800 265474 856
rect 265642 800 266026 856
rect 266194 800 266670 856
rect 266838 800 267222 856
rect 267390 800 267774 856
rect 267942 800 268326 856
rect 268494 800 268878 856
rect 269046 800 269430 856
rect 269598 800 269982 856
rect 270150 800 270534 856
rect 270702 800 271178 856
rect 271346 800 271730 856
rect 271898 800 272282 856
rect 272450 800 272834 856
rect 273002 800 273386 856
rect 273554 800 273938 856
rect 274106 800 274490 856
rect 274658 800 275042 856
rect 275210 800 275686 856
rect 275854 800 276238 856
rect 276406 800 276790 856
rect 276958 800 277342 856
rect 277510 800 277894 856
rect 278062 800 278446 856
rect 278614 800 278998 856
rect 279166 800 279550 856
<< metal3 >>
rect 0 224952 800 225072
rect 0 194896 800 195016
rect 0 164976 800 165096
rect 0 134920 800 135040
rect 0 104864 800 104984
rect 0 74944 800 75064
rect 0 44888 800 45008
rect 0 14968 800 15088
rect 279200 215976 280000 216096
rect 279200 167968 280000 168088
rect 279200 119960 280000 120080
rect 279200 71952 280000 72072
rect 279200 23944 280000 24064
<< obsm3 >>
rect 4208 2143 273871 237761
<< metal4 >>
rect 4208 2128 4528 237776
rect 4868 2176 5188 237728
rect 5528 2176 5848 237728
rect 6188 2176 6508 237728
rect 19568 2128 19888 237776
rect 20228 2176 20548 237728
rect 20888 2176 21208 237728
rect 21548 2176 21868 237728
rect 34928 2128 35248 237776
rect 35588 2176 35908 237728
rect 36248 2176 36568 237728
rect 36908 2176 37228 237728
rect 50288 2128 50608 237776
rect 50948 2176 51268 237728
rect 51608 2176 51928 237728
rect 52268 2176 52588 237728
rect 65648 2128 65968 237776
rect 66308 2176 66628 237728
rect 66968 2176 67288 237728
rect 67628 2176 67948 237728
rect 81008 2128 81328 237776
rect 81668 2176 81988 237728
rect 82328 2176 82648 237728
rect 82988 2176 83308 237728
rect 96368 2128 96688 237776
rect 97028 2176 97348 237728
rect 97688 2176 98008 237728
rect 98348 2176 98668 237728
rect 111728 2128 112048 237776
rect 112388 2176 112708 237728
rect 113048 2176 113368 237728
rect 113708 2176 114028 237728
rect 127088 2128 127408 237776
rect 127748 2176 128068 237728
rect 128408 2176 128728 237728
rect 129068 2176 129388 237728
rect 142448 2128 142768 237776
rect 143108 2176 143428 237728
rect 143768 2176 144088 237728
rect 144428 2176 144748 237728
rect 157808 2128 158128 237776
rect 158468 2176 158788 237728
rect 159128 2176 159448 237728
rect 159788 2176 160108 237728
rect 173168 2128 173488 237776
rect 173828 2176 174148 237728
rect 174488 2176 174808 237728
rect 175148 2176 175468 237728
rect 188528 2128 188848 237776
rect 189188 2176 189508 237728
rect 189848 2176 190168 237728
rect 190508 2176 190828 237728
rect 203888 2128 204208 237776
rect 204548 2176 204868 237728
rect 205208 2176 205528 237728
rect 205868 2176 206188 237728
rect 219248 2128 219568 237776
rect 219908 2176 220228 237728
rect 220568 2176 220888 237728
rect 221228 2176 221548 237728
rect 234608 2128 234928 237776
rect 235268 2176 235588 237728
rect 235928 2176 236248 237728
rect 236588 2176 236908 237728
rect 249968 2128 250288 237776
rect 250628 2176 250948 237728
rect 251288 2176 251608 237728
rect 251948 2176 252268 237728
rect 265328 2128 265648 237776
rect 265988 2176 266308 237728
rect 266648 2176 266968 237728
rect 267308 2176 267628 237728
<< obsm4 >>
rect 46979 5339 50208 211037
rect 50688 5339 50868 211037
rect 51348 5339 51528 211037
rect 52008 5339 52188 211037
rect 52668 5339 65568 211037
rect 66048 5339 66228 211037
rect 66708 5339 66888 211037
rect 67368 5339 67548 211037
rect 68028 5339 80928 211037
rect 81408 5339 81588 211037
rect 82068 5339 82248 211037
rect 82728 5339 82908 211037
rect 83388 5339 96288 211037
rect 96768 5339 96948 211037
rect 97428 5339 97608 211037
rect 98088 5339 98268 211037
rect 98748 5339 111648 211037
rect 112128 5339 112308 211037
rect 112788 5339 112968 211037
rect 113448 5339 113628 211037
rect 114108 5339 127008 211037
rect 127488 5339 127668 211037
rect 128148 5339 128328 211037
rect 128808 5339 128988 211037
rect 129468 5339 142368 211037
rect 142848 5339 143028 211037
rect 143508 5339 143688 211037
rect 144168 5339 144348 211037
rect 144828 5339 157728 211037
rect 158208 5339 158388 211037
rect 158868 5339 159048 211037
rect 159528 5339 159708 211037
rect 160188 5339 173088 211037
rect 173568 5339 173748 211037
rect 174228 5339 174408 211037
rect 174888 5339 175068 211037
rect 175548 5339 186517 211037
<< obsm5 >>
rect 116588 136180 134572 144660
<< labels >>
rlabel metal2 s 276294 0 276350 800 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 263138 239200 263194 240000 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 279200 71952 280000 72072 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 0 104864 800 104984 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 277950 0 278006 800 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 265346 239200 265402 240000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 279200 119960 280000 120080 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal3 s 0 134920 800 135040 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 278502 0 278558 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 267554 239200 267610 240000 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 279054 0 279110 800 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 256422 239200 256478 240000 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 279200 167968 280000 168088 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 269854 239200 269910 240000 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 279200 215976 280000 216096 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 272062 239200 272118 240000 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 274270 239200 274326 240000 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 279606 0 279662 800 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 164976 800 165096 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 194896 800 195016 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 276570 239200 276626 240000 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 0 224952 800 225072 6 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal2 s 276846 0 276902 800 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 278778 239200 278834 240000 6 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal3 s 279200 23944 280000 24064 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 0 14968 800 15088 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal2 s 258630 239200 258686 240000 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal2 s 260838 239200 260894 240000 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal2 s 277398 0 277454 800 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal3 s 0 44888 800 45008 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal3 s 0 74944 800 75064 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 1122 239200 1178 240000 6 io_in[0]
port 32 nsew signal input
rlabel metal2 s 68282 239200 68338 240000 6 io_in[10]
port 33 nsew signal input
rlabel metal2 s 74998 239200 75054 240000 6 io_in[11]
port 34 nsew signal input
rlabel metal2 s 81714 239200 81770 240000 6 io_in[12]
port 35 nsew signal input
rlabel metal2 s 88430 239200 88486 240000 6 io_in[13]
port 36 nsew signal input
rlabel metal2 s 95146 239200 95202 240000 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 101862 239200 101918 240000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 108578 239200 108634 240000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 115294 239200 115350 240000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 122010 239200 122066 240000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 128726 239200 128782 240000 6 io_in[19]
port 42 nsew signal input
rlabel metal2 s 7838 239200 7894 240000 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 135442 239200 135498 240000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 142158 239200 142214 240000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 148874 239200 148930 240000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 155590 239200 155646 240000 6 io_in[23]
port 47 nsew signal input
rlabel metal2 s 162306 239200 162362 240000 6 io_in[24]
port 48 nsew signal input
rlabel metal2 s 169022 239200 169078 240000 6 io_in[25]
port 49 nsew signal input
rlabel metal2 s 175738 239200 175794 240000 6 io_in[26]
port 50 nsew signal input
rlabel metal2 s 182454 239200 182510 240000 6 io_in[27]
port 51 nsew signal input
rlabel metal2 s 189170 239200 189226 240000 6 io_in[28]
port 52 nsew signal input
rlabel metal2 s 195886 239200 195942 240000 6 io_in[29]
port 53 nsew signal input
rlabel metal2 s 14554 239200 14610 240000 6 io_in[2]
port 54 nsew signal input
rlabel metal2 s 202602 239200 202658 240000 6 io_in[30]
port 55 nsew signal input
rlabel metal2 s 209318 239200 209374 240000 6 io_in[31]
port 56 nsew signal input
rlabel metal2 s 216126 239200 216182 240000 6 io_in[32]
port 57 nsew signal input
rlabel metal2 s 222842 239200 222898 240000 6 io_in[33]
port 58 nsew signal input
rlabel metal2 s 229558 239200 229614 240000 6 io_in[34]
port 59 nsew signal input
rlabel metal2 s 236274 239200 236330 240000 6 io_in[35]
port 60 nsew signal input
rlabel metal2 s 242990 239200 243046 240000 6 io_in[36]
port 61 nsew signal input
rlabel metal2 s 249706 239200 249762 240000 6 io_in[37]
port 62 nsew signal input
rlabel metal2 s 21270 239200 21326 240000 6 io_in[3]
port 63 nsew signal input
rlabel metal2 s 27986 239200 28042 240000 6 io_in[4]
port 64 nsew signal input
rlabel metal2 s 34702 239200 34758 240000 6 io_in[5]
port 65 nsew signal input
rlabel metal2 s 41418 239200 41474 240000 6 io_in[6]
port 66 nsew signal input
rlabel metal2 s 48134 239200 48190 240000 6 io_in[7]
port 67 nsew signal input
rlabel metal2 s 54850 239200 54906 240000 6 io_in[8]
port 68 nsew signal input
rlabel metal2 s 61566 239200 61622 240000 6 io_in[9]
port 69 nsew signal input
rlabel metal2 s 3330 239200 3386 240000 6 io_oeb[0]
port 70 nsew signal output
rlabel metal2 s 70490 239200 70546 240000 6 io_oeb[10]
port 71 nsew signal output
rlabel metal2 s 77206 239200 77262 240000 6 io_oeb[11]
port 72 nsew signal output
rlabel metal2 s 83922 239200 83978 240000 6 io_oeb[12]
port 73 nsew signal output
rlabel metal2 s 90638 239200 90694 240000 6 io_oeb[13]
port 74 nsew signal output
rlabel metal2 s 97354 239200 97410 240000 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 104070 239200 104126 240000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 110786 239200 110842 240000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 117502 239200 117558 240000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 124218 239200 124274 240000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 130934 239200 130990 240000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal2 s 10046 239200 10102 240000 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 137650 239200 137706 240000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 144458 239200 144514 240000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 151174 239200 151230 240000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 157890 239200 157946 240000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal2 s 164606 239200 164662 240000 6 io_oeb[24]
port 86 nsew signal output
rlabel metal2 s 171322 239200 171378 240000 6 io_oeb[25]
port 87 nsew signal output
rlabel metal2 s 178038 239200 178094 240000 6 io_oeb[26]
port 88 nsew signal output
rlabel metal2 s 184754 239200 184810 240000 6 io_oeb[27]
port 89 nsew signal output
rlabel metal2 s 191470 239200 191526 240000 6 io_oeb[28]
port 90 nsew signal output
rlabel metal2 s 198186 239200 198242 240000 6 io_oeb[29]
port 91 nsew signal output
rlabel metal2 s 16762 239200 16818 240000 6 io_oeb[2]
port 92 nsew signal output
rlabel metal2 s 204902 239200 204958 240000 6 io_oeb[30]
port 93 nsew signal output
rlabel metal2 s 211618 239200 211674 240000 6 io_oeb[31]
port 94 nsew signal output
rlabel metal2 s 218334 239200 218390 240000 6 io_oeb[32]
port 95 nsew signal output
rlabel metal2 s 225050 239200 225106 240000 6 io_oeb[33]
port 96 nsew signal output
rlabel metal2 s 231766 239200 231822 240000 6 io_oeb[34]
port 97 nsew signal output
rlabel metal2 s 238482 239200 238538 240000 6 io_oeb[35]
port 98 nsew signal output
rlabel metal2 s 245198 239200 245254 240000 6 io_oeb[36]
port 99 nsew signal output
rlabel metal2 s 251914 239200 251970 240000 6 io_oeb[37]
port 100 nsew signal output
rlabel metal2 s 23478 239200 23534 240000 6 io_oeb[3]
port 101 nsew signal output
rlabel metal2 s 30194 239200 30250 240000 6 io_oeb[4]
port 102 nsew signal output
rlabel metal2 s 36910 239200 36966 240000 6 io_oeb[5]
port 103 nsew signal output
rlabel metal2 s 43626 239200 43682 240000 6 io_oeb[6]
port 104 nsew signal output
rlabel metal2 s 50342 239200 50398 240000 6 io_oeb[7]
port 105 nsew signal output
rlabel metal2 s 57058 239200 57114 240000 6 io_oeb[8]
port 106 nsew signal output
rlabel metal2 s 63774 239200 63830 240000 6 io_oeb[9]
port 107 nsew signal output
rlabel metal2 s 5538 239200 5594 240000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 72790 239200 72846 240000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 79506 239200 79562 240000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 86222 239200 86278 240000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 92938 239200 92994 240000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 99654 239200 99710 240000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 106370 239200 106426 240000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 113086 239200 113142 240000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 119802 239200 119858 240000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 126518 239200 126574 240000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 133234 239200 133290 240000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 12254 239200 12310 240000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 139950 239200 140006 240000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 146666 239200 146722 240000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 153382 239200 153438 240000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 160098 239200 160154 240000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 166814 239200 166870 240000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 173530 239200 173586 240000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 180246 239200 180302 240000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 186962 239200 187018 240000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 193678 239200 193734 240000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 200394 239200 200450 240000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 18970 239200 19026 240000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 207110 239200 207166 240000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 213826 239200 213882 240000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 220542 239200 220598 240000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 227258 239200 227314 240000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 233974 239200 234030 240000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 240690 239200 240746 240000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 247406 239200 247462 240000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 254122 239200 254178 240000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 25686 239200 25742 240000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 32402 239200 32458 240000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 39118 239200 39174 240000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 45834 239200 45890 240000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 52550 239200 52606 240000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 59266 239200 59322 240000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 65982 239200 66038 240000 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 228914 0 228970 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 230662 0 230718 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 232318 0 232374 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 233974 0 234030 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 237378 0 237434 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 239126 0 239182 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 240782 0 240838 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 242438 0 242494 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 244186 0 244242 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 245842 0 245898 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 247498 0 247554 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 249246 0 249302 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 250902 0 250958 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 252558 0 252614 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 254306 0 254362 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 257710 0 257766 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 259366 0 259422 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 261022 0 261078 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 262770 0 262826 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 264426 0 264482 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 266082 0 266138 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 267830 0 267886 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 269486 0 269542 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 271234 0 271290 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 272890 0 272946 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 274546 0 274602 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 174910 0 174966 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 176566 0 176622 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 179970 0 180026 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 181626 0 181682 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 185030 0 185086 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 190090 0 190146 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 191746 0 191802 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 195150 0 195206 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 196806 0 196862 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 200210 0 200266 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 201866 0 201922 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 205270 0 205326 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 212078 0 212134 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 213734 0 213790 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 217138 0 217194 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 218794 0 218850 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 223854 0 223910 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 225602 0 225658 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 229466 0 229522 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 231214 0 231270 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 232870 0 232926 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 234618 0 234674 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 236274 0 236330 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 237930 0 237986 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 239678 0 239734 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 241334 0 241390 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 242990 0 243046 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 244738 0 244794 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 246394 0 246450 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 248142 0 248198 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 249798 0 249854 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 251454 0 251510 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 253202 0 253258 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 254858 0 254914 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 256514 0 256570 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 258262 0 258318 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 259918 0 259974 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 261574 0 261630 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 263322 0 263378 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 264978 0 265034 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 266726 0 266782 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 268382 0 268438 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 270038 0 270094 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 271786 0 271842 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 273442 0 273498 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 275098 0 275154 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 123022 0 123078 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 134890 0 134946 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 141606 0 141662 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 145010 0 145066 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 156878 0 156934 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 158534 0 158590 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 160190 0 160246 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 165250 0 165306 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 166998 0 167054 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 168654 0 168710 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 170402 0 170458 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 173714 0 173770 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 175462 0 175518 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 177118 0 177174 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 178774 0 178830 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 180522 0 180578 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 182178 0 182234 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 183926 0 183982 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 185582 0 185638 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 187238 0 187294 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 188986 0 189042 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 190642 0 190698 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 192298 0 192354 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 194046 0 194102 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 195702 0 195758 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 197358 0 197414 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 199106 0 199162 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 200762 0 200818 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 202510 0 202566 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 205822 0 205878 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 207570 0 207626 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 209226 0 209282 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 212630 0 212686 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 214286 0 214342 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 216034 0 216090 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 217690 0 217746 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 219346 0 219402 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 221094 0 221150 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 222750 0 222806 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 224406 0 224462 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 226154 0 226210 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 227810 0 227866 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 230110 0 230166 800 6 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 231766 0 231822 800 6 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 233422 0 233478 800 6 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 235170 0 235226 800 6 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 236826 0 236882 800 6 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 238482 0 238538 800 6 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 241886 0 241942 800 6 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 243634 0 243690 800 6 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 245290 0 245346 800 6 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 246946 0 247002 800 6 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 248694 0 248750 800 6 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 250350 0 250406 800 6 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 252006 0 252062 800 6 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 253754 0 253810 800 6 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 255410 0 255466 800 6 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 257066 0 257122 800 6 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 258814 0 258870 800 6 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 260470 0 260526 800 6 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 262218 0 262274 800 6 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 263874 0 263930 800 6 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 265530 0 265586 800 6 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 267278 0 267334 800 6 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 268934 0 268990 800 6 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 270590 0 270646 800 6 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 272338 0 272394 800 6 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 273994 0 274050 800 6 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 275742 0 275798 800 6 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 152370 0 152426 800 6 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 169206 0 169262 800 6 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 176014 0 176070 800 6 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 181074 0 181130 800 6 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 182730 0 182786 800 6 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 192850 0 192906 800 6 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 194598 0 194654 800 6 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 196254 0 196310 800 6 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 201314 0 201370 800 6 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 206374 0 206430 800 6 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 208122 0 208178 800 6 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 211526 0 211582 800 6 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 214838 0 214894 800 6 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 216586 0 216642 800 6 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 221646 0 221702 800 6 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 223302 0 223358 800 6 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 224958 0 225014 800 6 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 226706 0 226762 800 6 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 228362 0 228418 800 6 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 530 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 531 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 532 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 wbs_adr_i[0]
port 533 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[10]
port 534 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[11]
port 535 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_adr_i[12]
port 536 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[13]
port 537 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[14]
port 538 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[15]
port 539 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[16]
port 540 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[17]
port 541 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[18]
port 542 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_adr_i[19]
port 543 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[1]
port 544 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_adr_i[20]
port 545 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_adr_i[21]
port 546 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 wbs_adr_i[22]
port 547 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 wbs_adr_i[23]
port 548 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[24]
port 549 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 wbs_adr_i[25]
port 550 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 wbs_adr_i[26]
port 551 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 wbs_adr_i[27]
port 552 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_adr_i[28]
port 553 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 wbs_adr_i[29]
port 554 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[2]
port 555 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 wbs_adr_i[30]
port 556 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 wbs_adr_i[31]
port 557 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[3]
port 558 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[4]
port 559 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_adr_i[5]
port 560 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[6]
port 561 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[7]
port 562 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[8]
port 563 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[9]
port 564 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_cyc_i
port 565 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_i[0]
port 566 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_i[10]
port 567 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[11]
port 568 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[12]
port 569 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_i[13]
port 570 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[14]
port 571 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[15]
port 572 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[16]
port 573 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_i[17]
port 574 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[18]
port 575 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_i[19]
port 576 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[1]
port 577 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[20]
port 578 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_dat_i[21]
port 579 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_i[22]
port 580 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_i[23]
port 581 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_i[24]
port 582 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_dat_i[25]
port 583 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_dat_i[26]
port 584 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 wbs_dat_i[27]
port 585 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_i[28]
port 586 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_dat_i[29]
port 587 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_i[2]
port 588 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 wbs_dat_i[30]
port 589 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 wbs_dat_i[31]
port 590 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[3]
port 591 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[4]
port 592 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[5]
port 593 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_i[6]
port 594 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[7]
port 595 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[8]
port 596 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[9]
port 597 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_o[0]
port 598 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[10]
port 599 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_o[11]
port 600 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_o[12]
port 601 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_o[13]
port 602 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_o[14]
port 603 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[15]
port 604 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[16]
port 605 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[17]
port 606 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[18]
port 607 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_o[19]
port 608 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_o[1]
port 609 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 wbs_dat_o[20]
port 610 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_o[21]
port 611 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_o[22]
port 612 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_o[23]
port 613 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[24]
port 614 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_o[25]
port 615 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_o[26]
port 616 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_o[27]
port 617 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_o[28]
port 618 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_o[29]
port 619 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[2]
port 620 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 wbs_dat_o[30]
port 621 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 wbs_dat_o[31]
port 622 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_o[3]
port 623 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[4]
port 624 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[5]
port 625 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[6]
port 626 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[7]
port 627 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[8]
port 628 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[9]
port 629 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 wbs_sel_i[0]
port 630 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_sel_i[1]
port 631 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_sel_i[2]
port 632 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_sel_i[3]
port 633 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_stb_i
port 634 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_we_i
port 635 nsew signal input
rlabel metal4 s 249968 2128 250288 237776 6 vccd1
port 636 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 237776 6 vccd1
port 637 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 237776 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 237776 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 237776 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 237776 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 237776 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 237776 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 237776 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 265328 2128 265648 237776 6 vssd1
port 645 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 237776 6 vssd1
port 646 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 237776 6 vssd1
port 647 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 237776 6 vssd1
port 648 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 237776 6 vssd1
port 649 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 237776 6 vssd1
port 650 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 237776 6 vssd1
port 651 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 237776 6 vssd1
port 652 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 237776 6 vssd1
port 653 nsew ground bidirectional
rlabel metal4 s 250628 2176 250948 237728 6 vccd2
port 654 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 237728 6 vccd2
port 655 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 237728 6 vccd2
port 656 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 237728 6 vccd2
port 657 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 237728 6 vccd2
port 658 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 237728 6 vccd2
port 659 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 237728 6 vccd2
port 660 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 237728 6 vccd2
port 661 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 237728 6 vccd2
port 662 nsew power bidirectional
rlabel metal4 s 265988 2176 266308 237728 6 vssd2
port 663 nsew ground bidirectional
rlabel metal4 s 235268 2176 235588 237728 6 vssd2
port 664 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 237728 6 vssd2
port 665 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 237728 6 vssd2
port 666 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 237728 6 vssd2
port 667 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 237728 6 vssd2
port 668 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 237728 6 vssd2
port 669 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 237728 6 vssd2
port 670 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 237728 6 vssd2
port 671 nsew ground bidirectional
rlabel metal4 s 251288 2176 251608 237728 6 vdda1
port 672 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 237728 6 vdda1
port 673 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 237728 6 vdda1
port 674 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 237728 6 vdda1
port 675 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 237728 6 vdda1
port 676 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 237728 6 vdda1
port 677 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 237728 6 vdda1
port 678 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 237728 6 vdda1
port 679 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 237728 6 vdda1
port 680 nsew power bidirectional
rlabel metal4 s 266648 2176 266968 237728 6 vssa1
port 681 nsew ground bidirectional
rlabel metal4 s 235928 2176 236248 237728 6 vssa1
port 682 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 237728 6 vssa1
port 683 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 237728 6 vssa1
port 684 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 237728 6 vssa1
port 685 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 237728 6 vssa1
port 686 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 237728 6 vssa1
port 687 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 237728 6 vssa1
port 688 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 237728 6 vssa1
port 689 nsew ground bidirectional
rlabel metal4 s 251948 2176 252268 237728 6 vdda2
port 690 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 237728 6 vdda2
port 691 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 237728 6 vdda2
port 692 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 237728 6 vdda2
port 693 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 237728 6 vdda2
port 694 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 237728 6 vdda2
port 695 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 237728 6 vdda2
port 696 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 237728 6 vdda2
port 697 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 237728 6 vdda2
port 698 nsew power bidirectional
rlabel metal4 s 267308 2176 267628 237728 6 vssa2
port 699 nsew ground bidirectional
rlabel metal4 s 236588 2176 236908 237728 6 vssa2
port 700 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 237728 6 vssa2
port 701 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 237728 6 vssa2
port 702 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 237728 6 vssa2
port 703 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 237728 6 vssa2
port 704 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 237728 6 vssa2
port 705 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 237728 6 vssa2
port 706 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 237728 6 vssa2
port 707 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 280000 240000
string LEFview TRUE
<< end >>
