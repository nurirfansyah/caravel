VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1906.770 2512.160 1907.090 2512.220 ;
        RECT 2570.090 2512.160 2570.410 2512.220 ;
        RECT 1906.770 2512.020 2570.410 2512.160 ;
        RECT 1906.770 2511.960 1907.090 2512.020 ;
        RECT 2570.090 2511.960 2570.410 2512.020 ;
        RECT 2570.090 34.240 2570.410 34.300 ;
        RECT 2900.830 34.240 2901.150 34.300 ;
        RECT 2570.090 34.100 2901.150 34.240 ;
        RECT 2570.090 34.040 2570.410 34.100 ;
        RECT 2900.830 34.040 2901.150 34.100 ;
      LAYER via ;
        RECT 1906.800 2511.960 1907.060 2512.220 ;
        RECT 2570.120 2511.960 2570.380 2512.220 ;
        RECT 2570.120 34.040 2570.380 34.300 ;
        RECT 2900.860 34.040 2901.120 34.300 ;
      LAYER met2 ;
        RECT 1906.800 2511.930 1907.060 2512.250 ;
        RECT 2570.120 2511.930 2570.380 2512.250 ;
        RECT 1906.860 2500.000 1907.000 2511.930 ;
        RECT 1906.790 2496.000 1907.070 2500.000 ;
        RECT 2570.180 34.330 2570.320 2511.930 ;
        RECT 2570.120 34.010 2570.380 34.330 ;
        RECT 2900.860 34.010 2901.120 34.330 ;
        RECT 2900.920 29.765 2901.060 34.010 ;
        RECT 2900.850 29.395 2901.130 29.765 ;
      LAYER via2 ;
        RECT 2900.850 29.440 2901.130 29.720 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 28.980 2924.800 30.180 ;
=======
        RECT 2900.825 29.730 2901.155 29.745 ;
        RECT 2917.600 29.730 2924.800 30.180 ;
        RECT 2900.825 29.430 2924.800 29.730 ;
        RECT 2900.825 29.415 2901.155 29.430 ;
        RECT 2917.600 28.980 2924.800 29.430 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1940.810 1697.180 1941.130 1697.240 ;
        RECT 2901.750 1697.180 2902.070 1697.240 ;
        RECT 1940.810 1697.040 2902.070 1697.180 ;
        RECT 1940.810 1696.980 1941.130 1697.040 ;
        RECT 2901.750 1696.980 2902.070 1697.040 ;
      LAYER via ;
        RECT 1940.840 1696.980 1941.100 1697.240 ;
        RECT 2901.780 1696.980 2902.040 1697.240 ;
      LAYER met2 ;
        RECT 2901.770 2375.395 2902.050 2375.765 ;
        RECT 1940.830 1700.000 1941.110 1704.000 ;
        RECT 1940.900 1697.270 1941.040 1700.000 ;
        RECT 2901.840 1697.270 2901.980 2375.395 ;
        RECT 1940.840 1696.950 1941.100 1697.270 ;
        RECT 2901.780 1696.950 2902.040 1697.270 ;
      LAYER via2 ;
        RECT 2901.770 2375.440 2902.050 2375.720 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2374.980 2924.800 2376.180 ;
=======
        RECT 2901.745 2375.730 2902.075 2375.745 ;
        RECT 2917.600 2375.730 2924.800 2376.180 ;
        RECT 2901.745 2375.430 2924.800 2375.730 ;
        RECT 2901.745 2375.415 2902.075 2375.430 ;
        RECT 2917.600 2374.980 2924.800 2375.430 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2064.625 2608.225 2065.715 2608.395 ;
        RECT 2147.425 2608.225 2148.515 2608.395 ;
        RECT 2713.225 2608.225 2714.315 2608.395 ;
      LAYER mcon ;
        RECT 2065.545 2608.225 2065.715 2608.395 ;
        RECT 2148.345 2608.225 2148.515 2608.395 ;
        RECT 2714.145 2608.225 2714.315 2608.395 ;
      LAYER met1 ;
        RECT 1963.350 2608.380 1963.670 2608.440 ;
        RECT 2064.565 2608.380 2064.855 2608.425 ;
        RECT 1963.350 2608.240 2064.855 2608.380 ;
        RECT 1963.350 2608.180 1963.670 2608.240 ;
        RECT 2064.565 2608.195 2064.855 2608.240 ;
        RECT 2065.485 2608.380 2065.775 2608.425 ;
        RECT 2147.365 2608.380 2147.655 2608.425 ;
        RECT 2065.485 2608.240 2147.655 2608.380 ;
        RECT 2065.485 2608.195 2065.775 2608.240 ;
        RECT 2147.365 2608.195 2147.655 2608.240 ;
        RECT 2148.285 2608.380 2148.575 2608.425 ;
        RECT 2713.165 2608.380 2713.455 2608.425 ;
        RECT 2148.285 2608.240 2713.455 2608.380 ;
        RECT 2148.285 2608.195 2148.575 2608.240 ;
        RECT 2713.165 2608.195 2713.455 2608.240 ;
        RECT 2714.085 2608.380 2714.375 2608.425 ;
        RECT 2900.830 2608.380 2901.150 2608.440 ;
        RECT 2714.085 2608.240 2901.150 2608.380 ;
        RECT 2714.085 2608.195 2714.375 2608.240 ;
        RECT 2900.830 2608.180 2901.150 2608.240 ;
      LAYER via ;
        RECT 1963.380 2608.180 1963.640 2608.440 ;
        RECT 2900.860 2608.180 2901.120 2608.440 ;
      LAYER met2 ;
        RECT 2900.850 2609.995 2901.130 2610.365 ;
        RECT 2900.920 2608.470 2901.060 2609.995 ;
        RECT 1963.380 2608.150 1963.640 2608.470 ;
        RECT 2900.860 2608.150 2901.120 2608.470 ;
        RECT 1963.440 1900.445 1963.580 2608.150 ;
        RECT 1963.370 1900.075 1963.650 1900.445 ;
      LAYER via2 ;
        RECT 2900.850 2610.040 2901.130 2610.320 ;
        RECT 1963.370 1900.120 1963.650 1900.400 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2609.580 2924.800 2610.780 ;
=======
        RECT 2900.825 2610.330 2901.155 2610.345 ;
        RECT 2917.600 2610.330 2924.800 2610.780 ;
        RECT 2900.825 2610.030 2924.800 2610.330 ;
        RECT 2900.825 2610.015 2901.155 2610.030 ;
        RECT 2917.600 2609.580 2924.800 2610.030 ;
        RECT 1946.000 1900.410 1950.000 1900.560 ;
        RECT 1963.345 1900.410 1963.675 1900.425 ;
        RECT 1946.000 1900.110 1963.675 1900.410 ;
        RECT 1946.000 1899.960 1950.000 1900.110 ;
        RECT 1963.345 1900.095 1963.675 1900.110 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1931.610 2842.980 1931.930 2843.040 ;
        RECT 2900.830 2842.980 2901.150 2843.040 ;
        RECT 1931.610 2842.840 2901.150 2842.980 ;
        RECT 1931.610 2842.780 1931.930 2842.840 ;
        RECT 2900.830 2842.780 2901.150 2842.840 ;
        RECT 1926.550 2514.540 1926.870 2514.600 ;
        RECT 1931.610 2514.540 1931.930 2514.600 ;
        RECT 1926.550 2514.400 1931.930 2514.540 ;
        RECT 1926.550 2514.340 1926.870 2514.400 ;
        RECT 1931.610 2514.340 1931.930 2514.400 ;
      LAYER via ;
        RECT 1931.640 2842.780 1931.900 2843.040 ;
        RECT 2900.860 2842.780 2901.120 2843.040 ;
        RECT 1926.580 2514.340 1926.840 2514.600 ;
        RECT 1931.640 2514.340 1931.900 2514.600 ;
      LAYER met2 ;
        RECT 2900.850 2844.595 2901.130 2844.965 ;
        RECT 2900.920 2843.070 2901.060 2844.595 ;
        RECT 1931.640 2842.750 1931.900 2843.070 ;
        RECT 2900.860 2842.750 2901.120 2843.070 ;
        RECT 1931.700 2514.630 1931.840 2842.750 ;
        RECT 1926.580 2514.310 1926.840 2514.630 ;
        RECT 1931.640 2514.310 1931.900 2514.630 ;
        RECT 1926.640 2500.000 1926.780 2514.310 ;
        RECT 1926.570 2496.000 1926.850 2500.000 ;
      LAYER via2 ;
        RECT 2900.850 2844.640 2901.130 2844.920 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2844.180 2924.800 2845.380 ;
=======
        RECT 2900.825 2844.930 2901.155 2844.945 ;
        RECT 2917.600 2844.930 2924.800 2845.380 ;
        RECT 2900.825 2844.630 2924.800 2844.930 ;
        RECT 2900.825 2844.615 2901.155 2844.630 ;
        RECT 2917.600 2844.180 2924.800 2844.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2028.670 3079.280 2028.990 3079.340 ;
        RECT 2042.930 3079.280 2043.250 3079.340 ;
        RECT 2028.670 3079.140 2043.250 3079.280 ;
        RECT 2028.670 3079.080 2028.990 3079.140 ;
        RECT 2042.930 3079.080 2043.250 3079.140 ;
        RECT 2669.910 3079.280 2670.230 3079.340 ;
        RECT 2704.410 3079.280 2704.730 3079.340 ;
        RECT 2669.910 3079.140 2704.730 3079.280 ;
        RECT 2669.910 3079.080 2670.230 3079.140 ;
        RECT 2704.410 3079.080 2704.730 3079.140 ;
      LAYER via ;
        RECT 2028.700 3079.080 2028.960 3079.340 ;
        RECT 2042.960 3079.080 2043.220 3079.340 ;
        RECT 2669.940 3079.080 2670.200 3079.340 ;
        RECT 2704.440 3079.080 2704.700 3079.340 ;
      LAYER met2 ;
        RECT 2028.690 3079.195 2028.970 3079.565 ;
        RECT 2028.700 3079.050 2028.960 3079.195 ;
        RECT 2042.960 3079.050 2043.220 3079.370 ;
        RECT 2207.630 3079.195 2207.910 3079.565 ;
        RECT 2669.930 3079.195 2670.210 3079.565 ;
        RECT 2704.430 3079.195 2704.710 3079.565 ;
        RECT 2787.230 3079.195 2787.510 3079.565 ;
        RECT 2043.020 3078.205 2043.160 3079.050 ;
        RECT 2090.330 3078.515 2090.610 3078.885 ;
        RECT 2042.950 3077.835 2043.230 3078.205 ;
        RECT 2090.400 3078.090 2090.540 3078.515 ;
        RECT 2090.790 3078.090 2091.070 3078.205 ;
        RECT 2090.400 3077.950 2091.070 3078.090 ;
        RECT 2090.790 3077.835 2091.070 3077.950 ;
        RECT 2207.700 3077.525 2207.840 3079.195 ;
        RECT 2669.940 3079.050 2670.200 3079.195 ;
        RECT 2704.440 3079.050 2704.700 3079.195 ;
        RECT 2787.300 3077.525 2787.440 3079.195 ;
        RECT 2207.630 3077.155 2207.910 3077.525 ;
        RECT 2787.230 3077.155 2787.510 3077.525 ;
        RECT 1942.210 1703.130 1942.490 1704.000 ;
        RECT 1943.130 1703.130 1943.410 1703.245 ;
        RECT 1942.210 1702.990 1943.410 1703.130 ;
        RECT 1942.210 1700.000 1942.490 1702.990 ;
        RECT 1943.130 1702.875 1943.410 1702.990 ;
      LAYER via2 ;
        RECT 2028.690 3079.240 2028.970 3079.520 ;
        RECT 2207.630 3079.240 2207.910 3079.520 ;
        RECT 2669.930 3079.240 2670.210 3079.520 ;
        RECT 2704.430 3079.240 2704.710 3079.520 ;
        RECT 2787.230 3079.240 2787.510 3079.520 ;
        RECT 2090.330 3078.560 2090.610 3078.840 ;
        RECT 2042.950 3077.880 2043.230 3078.160 ;
        RECT 2090.790 3077.880 2091.070 3078.160 ;
        RECT 2207.630 3077.200 2207.910 3077.480 ;
        RECT 2787.230 3077.200 2787.510 3077.480 ;
        RECT 1943.130 1702.920 1943.410 1703.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3078.780 2924.800 3079.980 ;
=======
        RECT 1943.310 3079.530 1943.690 3079.540 ;
        RECT 2028.665 3079.530 2028.995 3079.545 ;
        RECT 1943.310 3079.230 1966.650 3079.530 ;
        RECT 1943.310 3079.220 1943.690 3079.230 ;
        RECT 1966.350 3078.850 1966.650 3079.230 ;
        RECT 2015.110 3079.230 2028.995 3079.530 ;
        RECT 1966.350 3078.550 2014.490 3078.850 ;
        RECT 2014.190 3078.170 2014.490 3078.550 ;
        RECT 2015.110 3078.170 2015.410 3079.230 ;
        RECT 2028.665 3079.215 2028.995 3079.230 ;
        RECT 2207.605 3079.530 2207.935 3079.545 ;
        RECT 2669.905 3079.530 2670.235 3079.545 ;
        RECT 2207.605 3079.230 2256.450 3079.530 ;
        RECT 2207.605 3079.215 2207.935 3079.230 ;
        RECT 2090.305 3078.850 2090.635 3078.865 ;
        RECT 2173.310 3078.850 2173.690 3078.860 ;
        RECT 2076.750 3078.550 2090.635 3078.850 ;
        RECT 2014.190 3077.870 2015.410 3078.170 ;
        RECT 2042.925 3078.170 2043.255 3078.185 ;
        RECT 2076.750 3078.170 2077.050 3078.550 ;
        RECT 2090.305 3078.535 2090.635 3078.550 ;
        RECT 2139.310 3078.550 2173.690 3078.850 ;
        RECT 2256.150 3078.850 2256.450 3079.230 ;
        RECT 2304.910 3079.230 2353.050 3079.530 ;
        RECT 2256.150 3078.550 2304.290 3078.850 ;
        RECT 2042.925 3077.870 2077.050 3078.170 ;
        RECT 2090.765 3078.170 2091.095 3078.185 ;
        RECT 2139.310 3078.170 2139.610 3078.550 ;
        RECT 2173.310 3078.540 2173.690 3078.550 ;
        RECT 2090.765 3077.870 2139.610 3078.170 ;
        RECT 2303.990 3078.170 2304.290 3078.550 ;
        RECT 2304.910 3078.170 2305.210 3079.230 ;
        RECT 2352.750 3078.850 2353.050 3079.230 ;
        RECT 2401.510 3079.230 2449.650 3079.530 ;
        RECT 2352.750 3078.550 2400.890 3078.850 ;
        RECT 2303.990 3077.870 2305.210 3078.170 ;
        RECT 2400.590 3078.170 2400.890 3078.550 ;
        RECT 2401.510 3078.170 2401.810 3079.230 ;
        RECT 2449.350 3078.850 2449.650 3079.230 ;
        RECT 2498.110 3079.230 2546.250 3079.530 ;
        RECT 2449.350 3078.550 2497.490 3078.850 ;
        RECT 2400.590 3077.870 2401.810 3078.170 ;
        RECT 2497.190 3078.170 2497.490 3078.550 ;
        RECT 2498.110 3078.170 2498.410 3079.230 ;
        RECT 2545.950 3078.850 2546.250 3079.230 ;
        RECT 2594.710 3079.230 2670.235 3079.530 ;
        RECT 2545.950 3078.550 2594.090 3078.850 ;
        RECT 2497.190 3077.870 2498.410 3078.170 ;
        RECT 2593.790 3078.170 2594.090 3078.550 ;
        RECT 2594.710 3078.170 2595.010 3079.230 ;
        RECT 2669.905 3079.215 2670.235 3079.230 ;
        RECT 2704.405 3079.530 2704.735 3079.545 ;
        RECT 2787.205 3079.530 2787.535 3079.545 ;
        RECT 2917.600 3079.530 2924.800 3079.980 ;
        RECT 2704.405 3079.230 2718.290 3079.530 ;
        RECT 2704.405 3079.215 2704.735 3079.230 ;
        RECT 2593.790 3077.870 2595.010 3078.170 ;
        RECT 2717.990 3078.170 2718.290 3079.230 ;
        RECT 2787.205 3079.230 2836.050 3079.530 ;
        RECT 2787.205 3079.215 2787.535 3079.230 ;
        RECT 2752.910 3078.850 2753.290 3078.860 ;
        RECT 2718.910 3078.550 2753.290 3078.850 ;
        RECT 2835.750 3078.850 2836.050 3079.230 ;
        RECT 2916.710 3079.230 2924.800 3079.530 ;
        RECT 2916.710 3078.850 2917.010 3079.230 ;
        RECT 2835.750 3078.550 2883.890 3078.850 ;
        RECT 2718.910 3078.170 2719.210 3078.550 ;
        RECT 2752.910 3078.540 2753.290 3078.550 ;
        RECT 2717.990 3077.870 2719.210 3078.170 ;
        RECT 2883.590 3078.170 2883.890 3078.550 ;
        RECT 2884.510 3078.550 2917.010 3078.850 ;
        RECT 2917.600 3078.780 2924.800 3079.230 ;
        RECT 2884.510 3078.170 2884.810 3078.550 ;
        RECT 2883.590 3077.870 2884.810 3078.170 ;
        RECT 2042.925 3077.855 2043.255 3077.870 ;
        RECT 2090.765 3077.855 2091.095 3077.870 ;
        RECT 2173.310 3077.490 2173.690 3077.500 ;
        RECT 2207.605 3077.490 2207.935 3077.505 ;
        RECT 2173.310 3077.190 2207.935 3077.490 ;
        RECT 2173.310 3077.180 2173.690 3077.190 ;
        RECT 2207.605 3077.175 2207.935 3077.190 ;
        RECT 2752.910 3077.490 2753.290 3077.500 ;
        RECT 2787.205 3077.490 2787.535 3077.505 ;
        RECT 2752.910 3077.190 2787.535 3077.490 ;
        RECT 2752.910 3077.180 2753.290 3077.190 ;
        RECT 2787.205 3077.175 2787.535 3077.190 ;
        RECT 1943.105 1703.220 1943.435 1703.225 ;
        RECT 1943.105 1703.210 1943.690 1703.220 ;
        RECT 1942.880 1702.910 1943.690 1703.210 ;
        RECT 1943.105 1702.900 1943.690 1702.910 ;
        RECT 1943.105 1702.895 1943.435 1702.900 ;
      LAYER via3 ;
        RECT 1943.340 3079.220 1943.660 3079.540 ;
        RECT 2173.340 3078.540 2173.660 3078.860 ;
        RECT 2752.940 3078.540 2753.260 3078.860 ;
        RECT 2173.340 3077.180 2173.660 3077.500 ;
        RECT 2752.940 3077.180 2753.260 3077.500 ;
        RECT 1943.340 1702.900 1943.660 1703.220 ;
      LAYER met4 ;
        RECT 1943.335 3079.215 1943.665 3079.545 ;
        RECT 1943.350 1703.225 1943.650 3079.215 ;
        RECT 2173.335 3078.535 2173.665 3078.865 ;
        RECT 2752.935 3078.535 2753.265 3078.865 ;
        RECT 2173.350 3077.505 2173.650 3078.535 ;
        RECT 2752.950 3077.505 2753.250 3078.535 ;
        RECT 2173.335 3077.175 2173.665 3077.505 ;
        RECT 2752.935 3077.175 2753.265 3077.505 ;
        RECT 1943.335 1702.895 1943.665 1703.225 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1962.890 3312.180 1963.210 3312.240 ;
        RECT 2900.830 3312.180 2901.150 3312.240 ;
        RECT 1962.890 3312.040 2901.150 3312.180 ;
        RECT 1962.890 3311.980 1963.210 3312.040 ;
        RECT 2900.830 3311.980 2901.150 3312.040 ;
      LAYER via ;
        RECT 1962.920 3311.980 1963.180 3312.240 ;
        RECT 2900.860 3311.980 2901.120 3312.240 ;
      LAYER met2 ;
        RECT 2900.850 3313.795 2901.130 3314.165 ;
        RECT 2900.920 3312.270 2901.060 3313.795 ;
        RECT 1962.920 3311.950 1963.180 3312.270 ;
        RECT 2900.860 3311.950 2901.120 3312.270 ;
        RECT 1962.980 2033.725 1963.120 3311.950 ;
        RECT 1962.910 2033.355 1963.190 2033.725 ;
      LAYER via2 ;
        RECT 2900.850 3313.840 2901.130 3314.120 ;
        RECT 1962.910 2033.400 1963.190 2033.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3313.380 2924.800 3314.580 ;
=======
        RECT 2900.825 3314.130 2901.155 3314.145 ;
        RECT 2917.600 3314.130 2924.800 3314.580 ;
        RECT 2900.825 3313.830 2924.800 3314.130 ;
        RECT 2900.825 3313.815 2901.155 3313.830 ;
        RECT 2917.600 3313.380 2924.800 3313.830 ;
        RECT 1946.000 2033.690 1950.000 2033.840 ;
        RECT 1962.885 2033.690 1963.215 2033.705 ;
        RECT 1946.000 2033.390 1963.215 2033.690 ;
        RECT 1946.000 2033.240 1950.000 2033.390 ;
        RECT 1962.885 2033.375 1963.215 2033.390 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2879.090 3519.700 2879.650 3524.800 ;
=======
        RECT 2879.090 3517.600 2879.650 3524.800 ;
        RECT 2879.300 3501.845 2879.440 3517.600 ;
        RECT 2879.230 3501.475 2879.510 3501.845 ;
        RECT 1944.050 1703.130 1944.330 1704.000 ;
        RECT 1944.510 1703.130 1944.790 1703.245 ;
        RECT 1944.050 1702.990 1944.790 1703.130 ;
        RECT 1944.050 1700.000 1944.330 1702.990 ;
        RECT 1944.510 1702.875 1944.790 1702.990 ;
      LAYER via2 ;
        RECT 2879.230 3501.520 2879.510 3501.800 ;
        RECT 1944.510 1702.920 1944.790 1703.200 ;
      LAYER met3 ;
        RECT 1944.230 3501.810 1944.610 3501.820 ;
        RECT 2879.205 3501.810 2879.535 3501.825 ;
        RECT 1944.230 3501.510 2879.535 3501.810 ;
        RECT 1944.230 3501.500 1944.610 3501.510 ;
        RECT 2879.205 3501.495 2879.535 3501.510 ;
        RECT 1944.485 1703.220 1944.815 1703.225 ;
        RECT 1944.230 1703.210 1944.815 1703.220 ;
        RECT 1944.230 1702.910 1945.040 1703.210 ;
        RECT 1944.230 1702.900 1944.815 1702.910 ;
        RECT 1944.485 1702.895 1944.815 1702.900 ;
      LAYER via3 ;
        RECT 1944.260 3501.500 1944.580 3501.820 ;
        RECT 1944.260 1702.900 1944.580 1703.220 ;
      LAYER met4 ;
        RECT 1944.255 3501.495 1944.585 3501.825 ;
        RECT 1944.270 1703.225 1944.570 3501.495 ;
        RECT 1944.255 1702.895 1944.585 1703.225 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1938.510 3501.560 1938.830 3501.620 ;
        RECT 2554.910 3501.560 2555.230 3501.620 ;
        RECT 1938.510 3501.420 2555.230 3501.560 ;
        RECT 1938.510 3501.360 1938.830 3501.420 ;
        RECT 2554.910 3501.360 2555.230 3501.420 ;
        RECT 1932.990 2516.240 1933.310 2516.300 ;
        RECT 1938.510 2516.240 1938.830 2516.300 ;
        RECT 1932.990 2516.100 1938.830 2516.240 ;
        RECT 1932.990 2516.040 1933.310 2516.100 ;
        RECT 1938.510 2516.040 1938.830 2516.100 ;
      LAYER via ;
        RECT 1938.540 3501.360 1938.800 3501.620 ;
        RECT 2554.940 3501.360 2555.200 3501.620 ;
        RECT 1933.020 2516.040 1933.280 2516.300 ;
        RECT 1938.540 2516.040 1938.800 2516.300 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2554.790 3519.700 2555.350 3524.800 ;
=======
        RECT 2554.790 3517.600 2555.350 3524.800 ;
        RECT 2555.000 3501.650 2555.140 3517.600 ;
        RECT 1938.540 3501.330 1938.800 3501.650 ;
        RECT 2554.940 3501.330 2555.200 3501.650 ;
        RECT 1938.600 2516.330 1938.740 3501.330 ;
        RECT 1933.020 2516.010 1933.280 2516.330 ;
        RECT 1938.540 2516.010 1938.800 2516.330 ;
        RECT 1933.080 2500.000 1933.220 2516.010 ;
        RECT 1933.010 2496.000 1933.290 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2230.490 3519.700 2231.050 3524.800 ;
=======
        RECT 2230.490 3517.600 2231.050 3524.800 ;
        RECT 2230.700 3502.525 2230.840 3517.600 ;
        RECT 2230.630 3502.155 2230.910 3502.525 ;
        RECT 1944.970 1702.450 1945.250 1702.565 ;
        RECT 1945.430 1702.450 1945.710 1704.000 ;
        RECT 1944.970 1702.310 1945.710 1702.450 ;
        RECT 1944.970 1702.195 1945.250 1702.310 ;
        RECT 1945.430 1700.000 1945.710 1702.310 ;
      LAYER via2 ;
        RECT 2230.630 3502.200 2230.910 3502.480 ;
        RECT 1944.970 1702.240 1945.250 1702.520 ;
      LAYER met3 ;
        RECT 1945.150 3502.490 1945.530 3502.500 ;
        RECT 2230.605 3502.490 2230.935 3502.505 ;
        RECT 1945.150 3502.190 2230.935 3502.490 ;
        RECT 1945.150 3502.180 1945.530 3502.190 ;
        RECT 2230.605 3502.175 2230.935 3502.190 ;
        RECT 1944.945 1702.540 1945.275 1702.545 ;
        RECT 1944.945 1702.530 1945.530 1702.540 ;
        RECT 1944.720 1702.230 1945.530 1702.530 ;
        RECT 1944.945 1702.220 1945.530 1702.230 ;
        RECT 1944.945 1702.215 1945.275 1702.220 ;
      LAYER via3 ;
        RECT 1945.180 3502.180 1945.500 3502.500 ;
        RECT 1945.180 1702.220 1945.500 1702.540 ;
      LAYER met4 ;
        RECT 1945.175 3502.175 1945.505 3502.505 ;
        RECT 1945.190 1702.545 1945.490 3502.175 ;
        RECT 1945.175 1702.215 1945.505 1702.545 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1905.850 3502.240 1906.170 3502.300 ;
        RECT 1946.790 3502.240 1947.110 3502.300 ;
        RECT 1905.850 3502.100 1947.110 3502.240 ;
        RECT 1905.850 3502.040 1906.170 3502.100 ;
        RECT 1946.790 3502.040 1947.110 3502.100 ;
      LAYER via ;
        RECT 1905.880 3502.040 1906.140 3502.300 ;
        RECT 1946.820 3502.040 1947.080 3502.300 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1905.730 3519.700 1906.290 3524.800 ;
=======
        RECT 1905.730 3517.600 1906.290 3524.800 ;
        RECT 1905.940 3502.330 1906.080 3517.600 ;
        RECT 1905.880 3502.010 1906.140 3502.330 ;
        RECT 1946.820 3502.010 1947.080 3502.330 ;
        RECT 1946.880 1703.810 1947.020 3502.010 ;
        RECT 1947.270 1703.810 1947.550 1704.000 ;
        RECT 1946.880 1703.670 1947.550 1703.810 ;
        RECT 1947.270 1700.000 1947.550 1703.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1582.085 3422.525 1582.255 3429.835 ;
        RECT 1581.625 2946.525 1581.795 2994.635 ;
        RECT 1580.705 2656.505 1580.875 2704.615 ;
        RECT 1581.165 2559.945 1581.335 2596.155 ;
        RECT 1255.945 2496.025 1256.115 2496.875 ;
        RECT 1294.125 2496.195 1294.295 2496.875 ;
        RECT 1292.745 2496.025 1294.295 2496.195 ;
      LAYER mcon ;
        RECT 1582.085 3429.665 1582.255 3429.835 ;
        RECT 1581.625 2994.465 1581.795 2994.635 ;
        RECT 1580.705 2704.445 1580.875 2704.615 ;
        RECT 1581.165 2595.985 1581.335 2596.155 ;
        RECT 1255.945 2496.705 1256.115 2496.875 ;
        RECT 1294.125 2496.705 1294.295 2496.875 ;
      LAYER met1 ;
        RECT 1582.010 3429.820 1582.330 3429.880 ;
        RECT 1581.815 3429.680 1582.330 3429.820 ;
        RECT 1582.010 3429.620 1582.330 3429.680 ;
        RECT 1582.010 3422.680 1582.330 3422.740 ;
        RECT 1581.815 3422.540 1582.330 3422.680 ;
        RECT 1582.010 3422.480 1582.330 3422.540 ;
        RECT 1581.550 3326.120 1581.870 3326.180 ;
        RECT 1582.010 3326.120 1582.330 3326.180 ;
        RECT 1581.550 3325.980 1582.330 3326.120 ;
        RECT 1581.550 3325.920 1581.870 3325.980 ;
        RECT 1582.010 3325.920 1582.330 3325.980 ;
        RECT 1581.550 3298.580 1581.870 3298.640 ;
        RECT 1581.180 3298.440 1581.870 3298.580 ;
        RECT 1581.180 3298.300 1581.320 3298.440 ;
        RECT 1581.550 3298.380 1581.870 3298.440 ;
        RECT 1581.090 3298.040 1581.410 3298.300 ;
        RECT 1580.630 3153.400 1580.950 3153.460 ;
        RECT 1581.550 3153.400 1581.870 3153.460 ;
        RECT 1580.630 3153.260 1581.870 3153.400 ;
        RECT 1580.630 3153.200 1580.950 3153.260 ;
        RECT 1581.550 3153.200 1581.870 3153.260 ;
        RECT 1580.630 3056.840 1580.950 3056.900 ;
        RECT 1581.550 3056.840 1581.870 3056.900 ;
        RECT 1580.630 3056.700 1581.870 3056.840 ;
        RECT 1580.630 3056.640 1580.950 3056.700 ;
        RECT 1581.550 3056.640 1581.870 3056.700 ;
        RECT 1581.090 3008.700 1581.410 3008.960 ;
        RECT 1581.180 3008.560 1581.320 3008.700 ;
        RECT 1581.550 3008.560 1581.870 3008.620 ;
        RECT 1581.180 3008.420 1581.870 3008.560 ;
        RECT 1581.550 3008.360 1581.870 3008.420 ;
        RECT 1581.550 2994.620 1581.870 2994.680 ;
        RECT 1581.355 2994.480 1581.870 2994.620 ;
        RECT 1581.550 2994.420 1581.870 2994.480 ;
        RECT 1581.565 2946.680 1581.855 2946.725 ;
        RECT 1582.010 2946.680 1582.330 2946.740 ;
        RECT 1581.565 2946.540 1582.330 2946.680 ;
        RECT 1581.565 2946.495 1581.855 2946.540 ;
        RECT 1582.010 2946.480 1582.330 2946.540 ;
        RECT 1582.010 2912.340 1582.330 2912.400 ;
        RECT 1581.640 2912.200 1582.330 2912.340 ;
        RECT 1581.640 2911.720 1581.780 2912.200 ;
        RECT 1582.010 2912.140 1582.330 2912.200 ;
        RECT 1581.550 2911.460 1581.870 2911.720 ;
        RECT 1580.630 2863.720 1580.950 2863.780 ;
        RECT 1581.550 2863.720 1581.870 2863.780 ;
        RECT 1580.630 2863.580 1581.870 2863.720 ;
        RECT 1580.630 2863.520 1580.950 2863.580 ;
        RECT 1581.550 2863.520 1581.870 2863.580 ;
        RECT 1581.090 2753.220 1581.410 2753.280 ;
        RECT 1581.550 2753.220 1581.870 2753.280 ;
        RECT 1581.090 2753.080 1581.870 2753.220 ;
        RECT 1581.090 2753.020 1581.410 2753.080 ;
        RECT 1581.550 2753.020 1581.870 2753.080 ;
        RECT 1581.090 2719.220 1581.410 2719.280 ;
        RECT 1580.720 2719.080 1581.410 2719.220 ;
        RECT 1580.720 2718.600 1580.860 2719.080 ;
        RECT 1581.090 2719.020 1581.410 2719.080 ;
        RECT 1580.630 2718.340 1580.950 2718.600 ;
        RECT 1580.630 2704.600 1580.950 2704.660 ;
        RECT 1580.435 2704.460 1580.950 2704.600 ;
        RECT 1580.630 2704.400 1580.950 2704.460 ;
        RECT 1580.645 2656.660 1580.935 2656.705 ;
        RECT 1581.090 2656.660 1581.410 2656.720 ;
        RECT 1580.645 2656.520 1581.410 2656.660 ;
        RECT 1580.645 2656.475 1580.935 2656.520 ;
        RECT 1581.090 2656.460 1581.410 2656.520 ;
        RECT 1581.090 2622.460 1581.410 2622.720 ;
        RECT 1581.180 2621.700 1581.320 2622.460 ;
        RECT 1581.090 2621.440 1581.410 2621.700 ;
        RECT 1581.090 2596.140 1581.410 2596.200 ;
        RECT 1580.895 2596.000 1581.410 2596.140 ;
        RECT 1581.090 2595.940 1581.410 2596.000 ;
        RECT 1581.105 2560.100 1581.395 2560.145 ;
        RECT 1582.010 2560.100 1582.330 2560.160 ;
        RECT 1581.105 2559.960 1582.330 2560.100 ;
        RECT 1581.105 2559.915 1581.395 2559.960 ;
        RECT 1582.010 2559.900 1582.330 2559.960 ;
        RECT 1582.010 2526.100 1582.330 2526.160 ;
        RECT 1581.180 2525.960 1582.330 2526.100 ;
        RECT 1581.180 2525.480 1581.320 2525.960 ;
        RECT 1582.010 2525.900 1582.330 2525.960 ;
        RECT 1581.090 2525.220 1581.410 2525.480 ;
        RECT 1138.110 2496.860 1138.430 2496.920 ;
        RECT 1255.885 2496.860 1256.175 2496.905 ;
        RECT 1138.110 2496.720 1256.175 2496.860 ;
        RECT 1138.110 2496.660 1138.430 2496.720 ;
        RECT 1255.885 2496.675 1256.175 2496.720 ;
        RECT 1294.065 2496.860 1294.355 2496.905 ;
        RECT 1581.090 2496.860 1581.410 2496.920 ;
        RECT 1294.065 2496.720 1581.410 2496.860 ;
        RECT 1294.065 2496.675 1294.355 2496.720 ;
        RECT 1581.090 2496.660 1581.410 2496.720 ;
        RECT 1255.885 2496.180 1256.175 2496.225 ;
        RECT 1292.685 2496.180 1292.975 2496.225 ;
        RECT 1255.885 2496.040 1292.975 2496.180 ;
        RECT 1255.885 2495.995 1256.175 2496.040 ;
        RECT 1292.685 2495.995 1292.975 2496.040 ;
      LAYER via ;
        RECT 1582.040 3429.620 1582.300 3429.880 ;
        RECT 1582.040 3422.480 1582.300 3422.740 ;
        RECT 1581.580 3325.920 1581.840 3326.180 ;
        RECT 1582.040 3325.920 1582.300 3326.180 ;
        RECT 1581.580 3298.380 1581.840 3298.640 ;
        RECT 1581.120 3298.040 1581.380 3298.300 ;
        RECT 1580.660 3153.200 1580.920 3153.460 ;
        RECT 1581.580 3153.200 1581.840 3153.460 ;
        RECT 1580.660 3056.640 1580.920 3056.900 ;
        RECT 1581.580 3056.640 1581.840 3056.900 ;
        RECT 1581.120 3008.700 1581.380 3008.960 ;
        RECT 1581.580 3008.360 1581.840 3008.620 ;
        RECT 1581.580 2994.420 1581.840 2994.680 ;
        RECT 1582.040 2946.480 1582.300 2946.740 ;
        RECT 1582.040 2912.140 1582.300 2912.400 ;
        RECT 1581.580 2911.460 1581.840 2911.720 ;
        RECT 1580.660 2863.520 1580.920 2863.780 ;
        RECT 1581.580 2863.520 1581.840 2863.780 ;
        RECT 1581.120 2753.020 1581.380 2753.280 ;
        RECT 1581.580 2753.020 1581.840 2753.280 ;
        RECT 1581.120 2719.020 1581.380 2719.280 ;
        RECT 1580.660 2718.340 1580.920 2718.600 ;
        RECT 1580.660 2704.400 1580.920 2704.660 ;
        RECT 1581.120 2656.460 1581.380 2656.720 ;
        RECT 1581.120 2622.460 1581.380 2622.720 ;
        RECT 1581.120 2621.440 1581.380 2621.700 ;
        RECT 1581.120 2595.940 1581.380 2596.200 ;
        RECT 1582.040 2559.900 1582.300 2560.160 ;
        RECT 1582.040 2525.900 1582.300 2526.160 ;
        RECT 1581.120 2525.220 1581.380 2525.480 ;
        RECT 1138.140 2496.660 1138.400 2496.920 ;
        RECT 1581.120 2496.660 1581.380 2496.920 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1581.430 3519.700 1581.990 3524.800 ;
=======
        RECT 1581.430 3517.600 1581.990 3524.800 ;
        RECT 1581.640 3477.930 1581.780 3517.600 ;
        RECT 1581.640 3477.790 1582.240 3477.930 ;
        RECT 1582.100 3429.910 1582.240 3477.790 ;
        RECT 1582.040 3429.590 1582.300 3429.910 ;
        RECT 1582.040 3422.450 1582.300 3422.770 ;
        RECT 1582.100 3326.210 1582.240 3422.450 ;
        RECT 1581.580 3325.890 1581.840 3326.210 ;
        RECT 1582.040 3325.890 1582.300 3326.210 ;
        RECT 1581.640 3298.670 1581.780 3325.890 ;
        RECT 1581.580 3298.350 1581.840 3298.670 ;
        RECT 1581.120 3298.010 1581.380 3298.330 ;
        RECT 1581.180 3250.130 1581.320 3298.010 ;
        RECT 1581.180 3249.990 1581.780 3250.130 ;
        RECT 1581.640 3153.490 1581.780 3249.990 ;
        RECT 1580.660 3153.170 1580.920 3153.490 ;
        RECT 1581.580 3153.170 1581.840 3153.490 ;
        RECT 1580.720 3152.890 1580.860 3153.170 ;
        RECT 1580.720 3152.750 1581.320 3152.890 ;
        RECT 1581.180 3105.290 1581.320 3152.750 ;
        RECT 1581.180 3105.150 1581.780 3105.290 ;
        RECT 1581.640 3056.930 1581.780 3105.150 ;
        RECT 1580.660 3056.610 1580.920 3056.930 ;
        RECT 1581.580 3056.610 1581.840 3056.930 ;
        RECT 1580.720 3056.330 1580.860 3056.610 ;
        RECT 1580.720 3056.190 1581.320 3056.330 ;
        RECT 1581.180 3008.990 1581.320 3056.190 ;
        RECT 1581.120 3008.670 1581.380 3008.990 ;
        RECT 1581.580 3008.330 1581.840 3008.650 ;
        RECT 1581.640 2994.710 1581.780 3008.330 ;
        RECT 1581.580 2994.390 1581.840 2994.710 ;
        RECT 1582.040 2946.450 1582.300 2946.770 ;
        RECT 1582.100 2912.430 1582.240 2946.450 ;
        RECT 1582.040 2912.110 1582.300 2912.430 ;
        RECT 1581.580 2911.430 1581.840 2911.750 ;
        RECT 1581.640 2863.810 1581.780 2911.430 ;
        RECT 1580.660 2863.490 1580.920 2863.810 ;
        RECT 1581.580 2863.490 1581.840 2863.810 ;
        RECT 1580.720 2863.210 1580.860 2863.490 ;
        RECT 1580.720 2863.070 1581.320 2863.210 ;
        RECT 1581.180 2815.610 1581.320 2863.070 ;
        RECT 1581.180 2815.470 1581.780 2815.610 ;
        RECT 1581.640 2753.310 1581.780 2815.470 ;
        RECT 1581.120 2752.990 1581.380 2753.310 ;
        RECT 1581.580 2752.990 1581.840 2753.310 ;
        RECT 1581.180 2719.310 1581.320 2752.990 ;
        RECT 1581.120 2718.990 1581.380 2719.310 ;
        RECT 1580.660 2718.310 1580.920 2718.630 ;
        RECT 1580.720 2704.690 1580.860 2718.310 ;
        RECT 1580.660 2704.370 1580.920 2704.690 ;
        RECT 1581.120 2656.430 1581.380 2656.750 ;
        RECT 1581.180 2622.750 1581.320 2656.430 ;
        RECT 1581.120 2622.430 1581.380 2622.750 ;
        RECT 1581.120 2621.410 1581.380 2621.730 ;
        RECT 1581.180 2596.230 1581.320 2621.410 ;
        RECT 1581.120 2595.910 1581.380 2596.230 ;
        RECT 1582.040 2559.870 1582.300 2560.190 ;
        RECT 1582.100 2526.190 1582.240 2559.870 ;
        RECT 1582.040 2525.870 1582.300 2526.190 ;
        RECT 1581.120 2525.190 1581.380 2525.510 ;
        RECT 1581.180 2496.950 1581.320 2525.190 ;
        RECT 1138.140 2496.630 1138.400 2496.950 ;
        RECT 1581.120 2496.630 1581.380 2496.950 ;
        RECT 1138.200 2059.565 1138.340 2496.630 ;
        RECT 1138.130 2059.195 1138.410 2059.565 ;
      LAYER via2 ;
        RECT 1138.130 2059.240 1138.410 2059.520 ;
      LAYER met3 ;
        RECT 1138.105 2059.530 1138.435 2059.545 ;
        RECT 1150.000 2059.530 1154.000 2059.680 ;
        RECT 1138.105 2059.230 1154.000 2059.530 ;
        RECT 1138.105 2059.215 1138.435 2059.230 ;
        RECT 1150.000 2059.080 1154.000 2059.230 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1138.110 268.840 1138.430 268.900 ;
        RECT 2900.830 268.840 2901.150 268.900 ;
        RECT 1138.110 268.700 2901.150 268.840 ;
        RECT 1138.110 268.640 1138.430 268.700 ;
        RECT 2900.830 268.640 2901.150 268.700 ;
      LAYER via ;
        RECT 1138.140 268.640 1138.400 268.900 ;
        RECT 2900.860 268.640 2901.120 268.900 ;
      LAYER met2 ;
        RECT 1138.130 1739.595 1138.410 1739.965 ;
        RECT 1138.200 268.930 1138.340 1739.595 ;
        RECT 1138.140 268.610 1138.400 268.930 ;
        RECT 2900.860 268.610 2901.120 268.930 ;
        RECT 2900.920 264.365 2901.060 268.610 ;
        RECT 2900.850 263.995 2901.130 264.365 ;
      LAYER via2 ;
        RECT 1138.130 1739.640 1138.410 1739.920 ;
        RECT 2900.850 264.040 2901.130 264.320 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 263.580 2924.800 264.780 ;
=======
        RECT 1138.105 1739.930 1138.435 1739.945 ;
        RECT 1150.000 1739.930 1154.000 1740.080 ;
        RECT 1138.105 1739.630 1154.000 1739.930 ;
        RECT 1138.105 1739.615 1138.435 1739.630 ;
        RECT 1150.000 1739.480 1154.000 1739.630 ;
        RECT 2900.825 264.330 2901.155 264.345 ;
        RECT 2917.600 264.330 2924.800 264.780 ;
        RECT 2900.825 264.030 2924.800 264.330 ;
        RECT 2900.825 264.015 2901.155 264.030 ;
        RECT 2917.600 263.580 2924.800 264.030 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1293.665 2496.365 1293.835 2509.115 ;
      LAYER mcon ;
        RECT 1293.665 2508.945 1293.835 2509.115 ;
      LAYER met1 ;
        RECT 1257.250 3498.500 1257.570 3498.560 ;
        RECT 1262.310 3498.500 1262.630 3498.560 ;
        RECT 1257.250 3498.360 1262.630 3498.500 ;
        RECT 1257.250 3498.300 1257.570 3498.360 ;
        RECT 1262.310 3498.300 1262.630 3498.360 ;
        RECT 1262.310 2509.100 1262.630 2509.160 ;
        RECT 1293.605 2509.100 1293.895 2509.145 ;
        RECT 1262.310 2508.960 1293.895 2509.100 ;
        RECT 1262.310 2508.900 1262.630 2508.960 ;
        RECT 1293.605 2508.915 1293.895 2508.960 ;
        RECT 1293.605 2496.520 1293.895 2496.565 ;
        RECT 1959.670 2496.520 1959.990 2496.580 ;
        RECT 1293.605 2496.380 1959.990 2496.520 ;
        RECT 1293.605 2496.335 1293.895 2496.380 ;
        RECT 1959.670 2496.320 1959.990 2496.380 ;
      LAYER via ;
        RECT 1257.280 3498.300 1257.540 3498.560 ;
        RECT 1262.340 3498.300 1262.600 3498.560 ;
        RECT 1262.340 2508.900 1262.600 2509.160 ;
        RECT 1959.700 2496.320 1959.960 2496.580 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1257.130 3519.700 1257.690 3524.800 ;
=======
        RECT 1257.130 3517.600 1257.690 3524.800 ;
        RECT 1257.340 3498.590 1257.480 3517.600 ;
        RECT 1257.280 3498.270 1257.540 3498.590 ;
        RECT 1262.340 3498.270 1262.600 3498.590 ;
        RECT 1262.400 2509.190 1262.540 3498.270 ;
        RECT 1262.340 2508.870 1262.600 2509.190 ;
        RECT 1959.700 2496.290 1959.960 2496.610 ;
        RECT 1959.760 2167.005 1959.900 2496.290 ;
        RECT 1959.690 2166.635 1959.970 2167.005 ;
      LAYER via2 ;
        RECT 1959.690 2166.680 1959.970 2166.960 ;
      LAYER met3 ;
        RECT 1946.000 2166.970 1950.000 2167.120 ;
        RECT 1959.665 2166.970 1959.995 2166.985 ;
        RECT 1946.000 2166.670 1959.995 2166.970 ;
        RECT 1946.000 2166.520 1950.000 2166.670 ;
        RECT 1959.665 2166.655 1959.995 2166.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.490 3498.500 932.810 3498.560 ;
        RECT 938.010 3498.500 938.330 3498.560 ;
        RECT 932.490 3498.360 938.330 3498.500 ;
        RECT 932.490 3498.300 932.810 3498.360 ;
        RECT 938.010 3498.300 938.330 3498.360 ;
        RECT 938.010 1696.840 938.330 1696.900 ;
        RECT 1948.630 1696.840 1948.950 1696.900 ;
        RECT 938.010 1696.700 1948.950 1696.840 ;
        RECT 938.010 1696.640 938.330 1696.700 ;
        RECT 1948.630 1696.640 1948.950 1696.700 ;
      LAYER via ;
        RECT 932.520 3498.300 932.780 3498.560 ;
        RECT 938.040 3498.300 938.300 3498.560 ;
        RECT 938.040 1696.640 938.300 1696.900 ;
        RECT 1948.660 1696.640 1948.920 1696.900 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 932.370 3519.700 932.930 3524.800 ;
=======
        RECT 932.370 3517.600 932.930 3524.800 ;
        RECT 932.580 3498.590 932.720 3517.600 ;
        RECT 932.520 3498.270 932.780 3498.590 ;
        RECT 938.040 3498.270 938.300 3498.590 ;
        RECT 938.100 1696.930 938.240 3498.270 ;
        RECT 1948.650 1700.000 1948.930 1704.000 ;
        RECT 1948.720 1696.930 1948.860 1700.000 ;
        RECT 938.040 1696.610 938.300 1696.930 ;
        RECT 1948.660 1696.610 1948.920 1696.930 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 608.190 3498.500 608.510 3498.560 ;
        RECT 613.710 3498.500 614.030 3498.560 ;
        RECT 608.190 3498.360 614.030 3498.500 ;
        RECT 608.190 3498.300 608.510 3498.360 ;
        RECT 613.710 3498.300 614.030 3498.360 ;
        RECT 613.710 2522.020 614.030 2522.080 ;
        RECT 1939.890 2522.020 1940.210 2522.080 ;
        RECT 613.710 2521.880 1940.210 2522.020 ;
        RECT 613.710 2521.820 614.030 2521.880 ;
        RECT 1939.890 2521.820 1940.210 2521.880 ;
      LAYER via ;
        RECT 608.220 3498.300 608.480 3498.560 ;
        RECT 613.740 3498.300 614.000 3498.560 ;
        RECT 613.740 2521.820 614.000 2522.080 ;
        RECT 1939.920 2521.820 1940.180 2522.080 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 608.070 3519.700 608.630 3524.800 ;
=======
        RECT 608.070 3517.600 608.630 3524.800 ;
        RECT 608.280 3498.590 608.420 3517.600 ;
        RECT 608.220 3498.270 608.480 3498.590 ;
        RECT 613.740 3498.270 614.000 3498.590 ;
        RECT 613.800 2522.110 613.940 3498.270 ;
        RECT 613.740 2521.790 614.000 2522.110 ;
        RECT 1939.920 2521.790 1940.180 2522.110 ;
        RECT 1939.980 2500.000 1940.120 2521.790 ;
        RECT 1939.910 2496.000 1940.190 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 283.890 3500.880 284.210 3500.940 ;
        RECT 289.410 3500.880 289.730 3500.940 ;
        RECT 283.890 3500.740 289.730 3500.880 ;
        RECT 283.890 3500.680 284.210 3500.740 ;
        RECT 289.410 3500.680 289.730 3500.740 ;
        RECT 289.410 2145.640 289.730 2145.700 ;
        RECT 1131.670 2145.640 1131.990 2145.700 ;
        RECT 289.410 2145.500 1131.990 2145.640 ;
        RECT 289.410 2145.440 289.730 2145.500 ;
        RECT 1131.670 2145.440 1131.990 2145.500 ;
      LAYER via ;
        RECT 283.920 3500.680 284.180 3500.940 ;
        RECT 289.440 3500.680 289.700 3500.940 ;
        RECT 289.440 2145.440 289.700 2145.700 ;
        RECT 1131.700 2145.440 1131.960 2145.700 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 283.770 3519.700 284.330 3524.800 ;
=======
        RECT 283.770 3517.600 284.330 3524.800 ;
        RECT 283.980 3500.970 284.120 3517.600 ;
        RECT 283.920 3500.650 284.180 3500.970 ;
        RECT 289.440 3500.650 289.700 3500.970 ;
        RECT 289.500 2145.730 289.640 3500.650 ;
        RECT 289.440 2145.410 289.700 2145.730 ;
        RECT 1131.700 2145.410 1131.960 2145.730 ;
        RECT 1131.760 2139.805 1131.900 2145.410 ;
        RECT 1131.690 2139.435 1131.970 2139.805 ;
      LAYER via2 ;
        RECT 1131.690 2139.480 1131.970 2139.760 ;
      LAYER met3 ;
        RECT 1131.665 2139.770 1131.995 2139.785 ;
        RECT 1150.000 2139.770 1154.000 2139.920 ;
        RECT 1131.665 2139.470 1154.000 2139.770 ;
        RECT 1131.665 2139.455 1131.995 2139.470 ;
        RECT 1150.000 2139.320 1154.000 2139.470 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1569.680 3477.960 1582.700 3478.100 ;
        RECT 17.090 3477.760 17.410 3477.820 ;
        RECT 1569.680 3477.760 1569.820 3477.960 ;
        RECT 17.090 3477.620 1569.820 3477.760 ;
        RECT 1582.560 3477.760 1582.700 3477.960 ;
        RECT 1728.290 3477.760 1728.610 3477.820 ;
        RECT 1582.560 3477.620 1728.610 3477.760 ;
        RECT 17.090 3477.560 17.410 3477.620 ;
        RECT 1728.290 3477.560 1728.610 3477.620 ;
        RECT 1728.290 2517.940 1728.610 2518.000 ;
        RECT 1946.330 2517.940 1946.650 2518.000 ;
        RECT 1728.290 2517.800 1946.650 2517.940 ;
        RECT 1728.290 2517.740 1728.610 2517.800 ;
        RECT 1946.330 2517.740 1946.650 2517.800 ;
      LAYER via ;
        RECT 17.120 3477.560 17.380 3477.820 ;
        RECT 1728.320 3477.560 1728.580 3477.820 ;
        RECT 1728.320 2517.740 1728.580 2518.000 ;
        RECT 1946.360 2517.740 1946.620 2518.000 ;
      LAYER met2 ;
        RECT 17.110 3483.115 17.390 3483.485 ;
        RECT 17.180 3477.850 17.320 3483.115 ;
        RECT 17.120 3477.530 17.380 3477.850 ;
        RECT 1728.320 3477.530 1728.580 3477.850 ;
        RECT 1728.380 2518.030 1728.520 3477.530 ;
        RECT 1728.320 2517.710 1728.580 2518.030 ;
        RECT 1946.360 2517.710 1946.620 2518.030 ;
        RECT 1946.420 2500.000 1946.560 2517.710 ;
        RECT 1946.350 2496.000 1946.630 2500.000 ;
      LAYER via2 ;
        RECT 17.110 3483.160 17.390 3483.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3482.700 0.300 3483.900 ;
=======
        RECT -4.800 3483.450 2.400 3483.900 ;
        RECT 17.085 3483.450 17.415 3483.465 ;
        RECT -4.800 3483.150 17.415 3483.450 ;
        RECT -4.800 3482.700 2.400 3483.150 ;
        RECT 17.085 3483.135 17.415 3483.150 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3194.880 17.410 3194.940 ;
        RECT 1947.250 3194.880 1947.570 3194.940 ;
        RECT 17.090 3194.740 1947.570 3194.880 ;
        RECT 17.090 3194.680 17.410 3194.740 ;
        RECT 1947.250 3194.680 1947.570 3194.740 ;
      LAYER via ;
        RECT 17.120 3194.680 17.380 3194.940 ;
        RECT 1947.280 3194.680 1947.540 3194.940 ;
      LAYER met2 ;
        RECT 17.110 3195.475 17.390 3195.845 ;
        RECT 17.180 3194.970 17.320 3195.475 ;
        RECT 17.120 3194.650 17.380 3194.970 ;
        RECT 1947.280 3194.650 1947.540 3194.970 ;
        RECT 1947.340 2302.325 1947.480 3194.650 ;
        RECT 1947.270 2301.955 1947.550 2302.325 ;
      LAYER via2 ;
        RECT 17.110 3195.520 17.390 3195.800 ;
        RECT 1947.270 2302.000 1947.550 2302.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3195.060 0.300 3196.260 ;
=======
        RECT -4.800 3195.810 2.400 3196.260 ;
        RECT 17.085 3195.810 17.415 3195.825 ;
        RECT -4.800 3195.510 17.415 3195.810 ;
        RECT -4.800 3195.060 2.400 3195.510 ;
        RECT 17.085 3195.495 17.415 3195.510 ;
        RECT 1947.245 2302.290 1947.575 2302.305 ;
        RECT 1947.030 2301.975 1947.575 2302.290 ;
        RECT 1947.030 2300.400 1947.330 2301.975 ;
        RECT 1946.000 2299.800 1950.000 2300.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2905.200 17.410 2905.260 ;
        RECT 51.590 2905.200 51.910 2905.260 ;
        RECT 17.090 2905.060 51.910 2905.200 ;
        RECT 17.090 2905.000 17.410 2905.060 ;
        RECT 51.590 2905.000 51.910 2905.060 ;
        RECT 51.590 2221.800 51.910 2221.860 ;
        RECT 1131.670 2221.800 1131.990 2221.860 ;
        RECT 51.590 2221.660 1131.990 2221.800 ;
        RECT 51.590 2221.600 51.910 2221.660 ;
        RECT 1131.670 2221.600 1131.990 2221.660 ;
      LAYER via ;
        RECT 17.120 2905.000 17.380 2905.260 ;
        RECT 51.620 2905.000 51.880 2905.260 ;
        RECT 51.620 2221.600 51.880 2221.860 ;
        RECT 1131.700 2221.600 1131.960 2221.860 ;
      LAYER met2 ;
        RECT 17.110 2908.515 17.390 2908.885 ;
        RECT 17.180 2905.290 17.320 2908.515 ;
        RECT 17.120 2904.970 17.380 2905.290 ;
        RECT 51.620 2904.970 51.880 2905.290 ;
        RECT 51.680 2221.890 51.820 2904.970 ;
        RECT 51.620 2221.570 51.880 2221.890 ;
        RECT 1131.700 2221.570 1131.960 2221.890 ;
        RECT 1131.760 2219.365 1131.900 2221.570 ;
        RECT 1131.690 2218.995 1131.970 2219.365 ;
      LAYER via2 ;
        RECT 17.110 2908.560 17.390 2908.840 ;
        RECT 1131.690 2219.040 1131.970 2219.320 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2908.100 0.300 2909.300 ;
=======
        RECT -4.800 2908.850 2.400 2909.300 ;
        RECT 17.085 2908.850 17.415 2908.865 ;
        RECT -4.800 2908.550 17.415 2908.850 ;
        RECT -4.800 2908.100 2.400 2908.550 ;
        RECT 17.085 2908.535 17.415 2908.550 ;
        RECT 1131.665 2219.330 1131.995 2219.345 ;
        RECT 1150.000 2219.330 1154.000 2219.480 ;
        RECT 1131.665 2219.030 1154.000 2219.330 ;
        RECT 1131.665 2219.015 1131.995 2219.030 ;
        RECT 1150.000 2218.880 1154.000 2219.030 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 2615.180 16.490 2615.240 ;
        RECT 65.390 2615.180 65.710 2615.240 ;
        RECT 16.170 2615.040 65.710 2615.180 ;
        RECT 16.170 2614.980 16.490 2615.040 ;
        RECT 65.390 2614.980 65.710 2615.040 ;
        RECT 65.390 2304.420 65.710 2304.480 ;
        RECT 1131.670 2304.420 1131.990 2304.480 ;
        RECT 65.390 2304.280 1131.990 2304.420 ;
        RECT 65.390 2304.220 65.710 2304.280 ;
        RECT 1131.670 2304.220 1131.990 2304.280 ;
      LAYER via ;
        RECT 16.200 2614.980 16.460 2615.240 ;
        RECT 65.420 2614.980 65.680 2615.240 ;
        RECT 65.420 2304.220 65.680 2304.480 ;
        RECT 1131.700 2304.220 1131.960 2304.480 ;
      LAYER met2 ;
        RECT 16.190 2620.875 16.470 2621.245 ;
        RECT 16.260 2615.270 16.400 2620.875 ;
        RECT 16.200 2614.950 16.460 2615.270 ;
        RECT 65.420 2614.950 65.680 2615.270 ;
        RECT 65.480 2304.510 65.620 2614.950 ;
        RECT 65.420 2304.190 65.680 2304.510 ;
        RECT 1131.700 2304.190 1131.960 2304.510 ;
        RECT 1131.760 2299.605 1131.900 2304.190 ;
        RECT 1131.690 2299.235 1131.970 2299.605 ;
      LAYER via2 ;
        RECT 16.190 2620.920 16.470 2621.200 ;
        RECT 1131.690 2299.280 1131.970 2299.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2620.460 0.300 2621.660 ;
=======
        RECT -4.800 2621.210 2.400 2621.660 ;
        RECT 16.165 2621.210 16.495 2621.225 ;
        RECT -4.800 2620.910 16.495 2621.210 ;
        RECT -4.800 2620.460 2.400 2620.910 ;
        RECT 16.165 2620.895 16.495 2620.910 ;
        RECT 1131.665 2299.570 1131.995 2299.585 ;
        RECT 1150.000 2299.570 1154.000 2299.720 ;
        RECT 1131.665 2299.270 1154.000 2299.570 ;
        RECT 1131.665 2299.255 1131.995 2299.270 ;
        RECT 1150.000 2299.120 1154.000 2299.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2333.500 0.300 2334.700 ;
=======
        RECT 1946.000 2433.530 1950.000 2433.680 ;
        RECT 1959.870 2433.530 1960.250 2433.540 ;
        RECT 1946.000 2433.230 1960.250 2433.530 ;
        RECT 1946.000 2433.080 1950.000 2433.230 ;
        RECT 1959.870 2433.220 1960.250 2433.230 ;
        RECT 290.070 2341.050 290.450 2341.060 ;
        RECT 336.990 2341.050 337.370 2341.060 ;
        RECT 290.070 2340.750 337.370 2341.050 ;
        RECT 290.070 2340.740 290.450 2340.750 ;
        RECT 336.990 2340.740 337.370 2340.750 ;
        RECT 386.670 2341.050 387.050 2341.060 ;
        RECT 433.590 2341.050 433.970 2341.060 ;
        RECT 386.670 2340.750 433.970 2341.050 ;
        RECT 386.670 2340.740 387.050 2340.750 ;
        RECT 433.590 2340.740 433.970 2340.750 ;
        RECT 483.270 2341.050 483.650 2341.060 ;
        RECT 530.190 2341.050 530.570 2341.060 ;
        RECT 483.270 2340.750 530.570 2341.050 ;
        RECT 483.270 2340.740 483.650 2340.750 ;
        RECT 530.190 2340.740 530.570 2340.750 ;
        RECT 773.070 2341.050 773.450 2341.060 ;
        RECT 819.990 2341.050 820.370 2341.060 ;
        RECT 773.070 2340.750 820.370 2341.050 ;
        RECT 773.070 2340.740 773.450 2340.750 ;
        RECT 819.990 2340.740 820.370 2340.750 ;
        RECT 966.270 2341.050 966.650 2341.060 ;
        RECT 980.990 2341.050 981.370 2341.060 ;
        RECT 966.270 2340.750 981.370 2341.050 ;
        RECT 966.270 2340.740 966.650 2340.750 ;
        RECT 980.990 2340.740 981.370 2340.750 ;
        RECT 1062.870 2341.050 1063.250 2341.060 ;
        RECT 1109.790 2341.050 1110.170 2341.060 ;
        RECT 1062.870 2340.750 1110.170 2341.050 ;
        RECT 1062.870 2340.740 1063.250 2340.750 ;
        RECT 1109.790 2340.740 1110.170 2340.750 ;
        RECT -4.800 2334.250 2.400 2334.700 ;
        RECT 26.030 2334.250 26.410 2334.260 ;
        RECT -4.800 2333.950 26.410 2334.250 ;
        RECT -4.800 2333.500 2.400 2333.950 ;
        RECT 26.030 2333.940 26.410 2333.950 ;
      LAYER via3 ;
        RECT 1959.900 2433.220 1960.220 2433.540 ;
        RECT 290.100 2340.740 290.420 2341.060 ;
        RECT 337.020 2340.740 337.340 2341.060 ;
        RECT 386.700 2340.740 387.020 2341.060 ;
        RECT 433.620 2340.740 433.940 2341.060 ;
        RECT 483.300 2340.740 483.620 2341.060 ;
        RECT 530.220 2340.740 530.540 2341.060 ;
        RECT 773.100 2340.740 773.420 2341.060 ;
        RECT 820.020 2340.740 820.340 2341.060 ;
        RECT 966.300 2340.740 966.620 2341.060 ;
        RECT 981.020 2340.740 981.340 2341.060 ;
        RECT 1062.900 2340.740 1063.220 2341.060 ;
        RECT 1109.820 2340.740 1110.140 2341.060 ;
        RECT 26.060 2333.940 26.380 2334.260 ;
      LAYER met4 ;
        RECT 1959.895 2433.215 1960.225 2433.545 ;
        RECT 289.670 2340.310 290.850 2341.490 ;
        RECT 336.590 2340.310 337.770 2341.490 ;
        RECT 386.270 2340.310 387.450 2341.490 ;
        RECT 433.190 2340.310 434.370 2341.490 ;
        RECT 482.870 2340.310 484.050 2341.490 ;
        RECT 529.790 2340.310 530.970 2341.490 ;
        RECT 772.670 2340.310 773.850 2341.490 ;
        RECT 820.015 2340.735 820.345 2341.065 ;
        RECT 820.030 2334.690 820.330 2340.735 ;
        RECT 965.870 2340.310 967.050 2341.490 ;
        RECT 980.590 2340.310 981.770 2341.490 ;
        RECT 1062.470 2340.310 1063.650 2341.490 ;
        RECT 1109.815 2340.735 1110.145 2341.065 ;
        RECT 1109.830 2334.690 1110.130 2340.735 ;
        RECT 1159.990 2340.310 1161.170 2341.490 ;
        RECT 1182.990 2340.310 1184.170 2341.490 ;
        RECT 25.630 2333.510 26.810 2334.690 ;
        RECT 819.590 2333.510 820.770 2334.690 ;
        RECT 1109.390 2333.510 1110.570 2334.690 ;
        RECT 1160.430 2327.890 1160.730 2340.310 ;
        RECT 1183.430 2327.890 1183.730 2340.310 ;
        RECT 1959.910 2334.690 1960.210 2433.215 ;
        RECT 1959.470 2333.510 1960.650 2334.690 ;
        RECT 1159.990 2326.710 1161.170 2327.890 ;
        RECT 1182.990 2326.710 1184.170 2327.890 ;
      LAYER met5 ;
        RECT 59.460 2340.100 97.860 2341.700 ;
        RECT 59.460 2334.900 61.060 2340.100 ;
        RECT 25.420 2333.300 61.060 2334.900 ;
        RECT 96.260 2334.900 97.860 2340.100 ;
        RECT 143.180 2340.100 194.460 2341.700 ;
        RECT 143.180 2334.900 144.780 2340.100 ;
        RECT 96.260 2333.300 144.780 2334.900 ;
        RECT 192.860 2334.900 194.460 2340.100 ;
        RECT 239.780 2340.100 291.060 2341.700 ;
        RECT 336.380 2340.100 387.660 2341.700 ;
        RECT 432.980 2340.100 484.260 2341.700 ;
        RECT 529.580 2340.100 580.860 2341.700 ;
        RECT 239.780 2334.900 241.380 2340.100 ;
        RECT 192.860 2333.300 241.380 2334.900 ;
        RECT 579.260 2334.900 580.860 2340.100 ;
        RECT 626.180 2340.100 677.460 2341.700 ;
        RECT 626.180 2334.900 627.780 2340.100 ;
        RECT 579.260 2333.300 627.780 2334.900 ;
        RECT 675.860 2334.900 677.460 2340.100 ;
        RECT 722.780 2340.100 774.060 2341.700 ;
        RECT 833.180 2340.100 871.580 2341.700 ;
        RECT 722.780 2334.900 724.380 2340.100 ;
        RECT 833.180 2334.900 834.780 2340.100 ;
        RECT 675.860 2333.300 724.380 2334.900 ;
        RECT 819.380 2333.300 834.780 2334.900 ;
        RECT 869.980 2328.100 871.580 2340.100 ;
        RECT 929.780 2340.100 967.260 2341.700 ;
        RECT 980.380 2340.100 1014.180 2341.700 ;
        RECT 929.780 2334.900 931.380 2340.100 ;
        RECT 915.980 2333.300 931.380 2334.900 ;
        RECT 1012.580 2334.900 1014.180 2340.100 ;
        RECT 1026.380 2340.100 1063.860 2341.700 ;
        RECT 1122.980 2340.100 1161.380 2341.700 ;
        RECT 1182.780 2340.100 1207.380 2341.700 ;
        RECT 1026.380 2334.900 1027.980 2340.100 ;
        RECT 1122.980 2334.900 1124.580 2340.100 ;
        RECT 1205.780 2338.300 1207.380 2340.100 ;
        RECT 1217.740 2340.100 1257.060 2341.700 ;
        RECT 1217.740 2338.300 1219.340 2340.100 ;
        RECT 1205.780 2336.700 1219.340 2338.300 ;
        RECT 1255.460 2338.300 1257.060 2340.100 ;
        RECT 1316.180 2340.100 1354.580 2341.700 ;
        RECT 1255.460 2336.700 1303.980 2338.300 ;
        RECT 1012.580 2333.300 1027.980 2334.900 ;
        RECT 1109.180 2333.300 1124.580 2334.900 ;
        RECT 1302.380 2334.900 1303.980 2336.700 ;
        RECT 1316.180 2334.900 1317.780 2340.100 ;
        RECT 1302.380 2333.300 1317.780 2334.900 ;
        RECT 915.980 2328.100 917.580 2333.300 ;
        RECT 1352.980 2328.100 1354.580 2340.100 ;
        RECT 1412.780 2340.100 1451.180 2341.700 ;
        RECT 1412.780 2334.900 1414.380 2340.100 ;
        RECT 1398.980 2333.300 1414.380 2334.900 ;
        RECT 1398.980 2328.100 1400.580 2333.300 ;
        RECT 869.980 2326.500 917.580 2328.100 ;
        RECT 1159.780 2326.500 1184.380 2328.100 ;
        RECT 1352.980 2326.500 1400.580 2328.100 ;
        RECT 1449.580 2328.100 1451.180 2340.100 ;
        RECT 1509.380 2340.100 1547.780 2341.700 ;
        RECT 1509.380 2334.900 1510.980 2340.100 ;
        RECT 1495.580 2333.300 1510.980 2334.900 ;
        RECT 1495.580 2328.100 1497.180 2333.300 ;
        RECT 1449.580 2326.500 1497.180 2328.100 ;
        RECT 1546.180 2328.100 1547.780 2340.100 ;
        RECT 1605.980 2340.100 1644.380 2341.700 ;
        RECT 1605.980 2334.900 1607.580 2340.100 ;
        RECT 1592.180 2333.300 1607.580 2334.900 ;
        RECT 1592.180 2328.100 1593.780 2333.300 ;
        RECT 1546.180 2326.500 1593.780 2328.100 ;
        RECT 1642.780 2328.100 1644.380 2340.100 ;
        RECT 1702.580 2340.100 1740.980 2341.700 ;
        RECT 1702.580 2334.900 1704.180 2340.100 ;
        RECT 1688.780 2333.300 1704.180 2334.900 ;
        RECT 1688.780 2328.100 1690.380 2333.300 ;
        RECT 1642.780 2326.500 1690.380 2328.100 ;
        RECT 1739.380 2328.100 1740.980 2340.100 ;
        RECT 1799.180 2340.100 1837.580 2341.700 ;
        RECT 1799.180 2334.900 1800.780 2340.100 ;
        RECT 1785.380 2333.300 1800.780 2334.900 ;
        RECT 1785.380 2328.100 1786.980 2333.300 ;
        RECT 1739.380 2326.500 1786.980 2328.100 ;
        RECT 1835.980 2328.100 1837.580 2340.100 ;
        RECT 1895.780 2340.100 1933.260 2341.700 ;
        RECT 1895.780 2334.900 1897.380 2340.100 ;
        RECT 1881.980 2333.300 1897.380 2334.900 ;
        RECT 1931.660 2334.900 1933.260 2340.100 ;
        RECT 1931.660 2333.300 1960.860 2334.900 ;
        RECT 1881.980 2328.100 1883.580 2333.300 ;
        RECT 1835.980 2326.500 1883.580 2328.100 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 79.190 2373.780 79.510 2373.840 ;
        RECT 1137.650 2373.780 1137.970 2373.840 ;
        RECT 79.190 2373.640 1137.970 2373.780 ;
        RECT 79.190 2373.580 79.510 2373.640 ;
        RECT 1137.650 2373.580 1137.970 2373.640 ;
        RECT 14.330 2049.080 14.650 2049.140 ;
        RECT 79.190 2049.080 79.510 2049.140 ;
        RECT 14.330 2048.940 79.510 2049.080 ;
        RECT 14.330 2048.880 14.650 2048.940 ;
        RECT 79.190 2048.880 79.510 2048.940 ;
      LAYER via ;
        RECT 79.220 2373.580 79.480 2373.840 ;
        RECT 1137.680 2373.580 1137.940 2373.840 ;
        RECT 14.360 2048.880 14.620 2049.140 ;
        RECT 79.220 2048.880 79.480 2049.140 ;
      LAYER met2 ;
        RECT 1137.670 2378.795 1137.950 2379.165 ;
        RECT 1137.740 2373.870 1137.880 2378.795 ;
        RECT 79.220 2373.550 79.480 2373.870 ;
        RECT 1137.680 2373.550 1137.940 2373.870 ;
        RECT 79.280 2049.170 79.420 2373.550 ;
        RECT 14.360 2048.850 14.620 2049.170 ;
        RECT 79.220 2048.850 79.480 2049.170 ;
        RECT 14.420 2046.645 14.560 2048.850 ;
        RECT 14.350 2046.275 14.630 2046.645 ;
      LAYER via2 ;
        RECT 1137.670 2378.840 1137.950 2379.120 ;
        RECT 14.350 2046.320 14.630 2046.600 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2045.860 0.300 2047.060 ;
=======
        RECT 1137.645 2379.130 1137.975 2379.145 ;
        RECT 1150.000 2379.130 1154.000 2379.280 ;
        RECT 1137.645 2378.830 1154.000 2379.130 ;
        RECT 1137.645 2378.815 1137.975 2378.830 ;
        RECT 1150.000 2378.680 1154.000 2378.830 ;
        RECT -4.800 2046.610 2.400 2047.060 ;
        RECT 14.325 2046.610 14.655 2046.625 ;
        RECT -4.800 2046.310 14.655 2046.610 ;
        RECT -4.800 2045.860 2.400 2046.310 ;
        RECT 14.325 2046.295 14.655 2046.310 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1962.890 503.440 1963.210 503.500 ;
        RECT 2900.830 503.440 2901.150 503.500 ;
        RECT 1962.890 503.300 2901.150 503.440 ;
        RECT 1962.890 503.240 1963.210 503.300 ;
        RECT 2900.830 503.240 2901.150 503.300 ;
      LAYER via ;
        RECT 1962.920 503.240 1963.180 503.500 ;
        RECT 2900.860 503.240 2901.120 503.500 ;
      LAYER met2 ;
        RECT 1962.910 1766.795 1963.190 1767.165 ;
        RECT 1962.980 503.530 1963.120 1766.795 ;
        RECT 1962.920 503.210 1963.180 503.530 ;
        RECT 2900.860 503.210 2901.120 503.530 ;
        RECT 2900.920 498.965 2901.060 503.210 ;
        RECT 2900.850 498.595 2901.130 498.965 ;
      LAYER via2 ;
        RECT 1962.910 1766.840 1963.190 1767.120 ;
        RECT 2900.850 498.640 2901.130 498.920 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 498.180 2924.800 499.380 ;
=======
        RECT 1946.000 1767.130 1950.000 1767.280 ;
        RECT 1962.885 1767.130 1963.215 1767.145 ;
        RECT 1946.000 1766.830 1963.215 1767.130 ;
        RECT 1946.000 1766.680 1950.000 1766.830 ;
        RECT 1962.885 1766.815 1963.215 1766.830 ;
        RECT 2900.825 498.930 2901.155 498.945 ;
        RECT 2917.600 498.930 2924.800 499.380 ;
        RECT 2900.825 498.630 2924.800 498.930 ;
        RECT 2900.825 498.615 2901.155 498.630 ;
        RECT 2917.600 498.180 2924.800 498.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 86.090 2456.740 86.410 2456.800 ;
        RECT 1131.670 2456.740 1131.990 2456.800 ;
        RECT 86.090 2456.600 1131.990 2456.740 ;
        RECT 86.090 2456.540 86.410 2456.600 ;
        RECT 1131.670 2456.540 1131.990 2456.600 ;
        RECT 15.710 1766.200 16.030 1766.260 ;
        RECT 86.090 1766.200 86.410 1766.260 ;
        RECT 15.710 1766.060 86.410 1766.200 ;
        RECT 15.710 1766.000 16.030 1766.060 ;
        RECT 86.090 1766.000 86.410 1766.060 ;
      LAYER via ;
        RECT 86.120 2456.540 86.380 2456.800 ;
        RECT 1131.700 2456.540 1131.960 2456.800 ;
        RECT 15.740 1766.000 16.000 1766.260 ;
        RECT 86.120 1766.000 86.380 1766.260 ;
      LAYER met2 ;
        RECT 1131.690 2459.035 1131.970 2459.405 ;
        RECT 1131.760 2456.830 1131.900 2459.035 ;
        RECT 86.120 2456.510 86.380 2456.830 ;
        RECT 1131.700 2456.510 1131.960 2456.830 ;
        RECT 86.180 1766.290 86.320 2456.510 ;
        RECT 15.740 1765.970 16.000 1766.290 ;
        RECT 86.120 1765.970 86.380 1766.290 ;
        RECT 15.800 1759.685 15.940 1765.970 ;
        RECT 15.730 1759.315 16.010 1759.685 ;
      LAYER via2 ;
        RECT 1131.690 2459.080 1131.970 2459.360 ;
        RECT 15.730 1759.360 16.010 1759.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1758.900 0.300 1760.100 ;
=======
        RECT 1131.665 2459.370 1131.995 2459.385 ;
        RECT 1150.000 2459.370 1154.000 2459.520 ;
        RECT 1131.665 2459.070 1154.000 2459.370 ;
        RECT 1131.665 2459.055 1131.995 2459.070 ;
        RECT 1150.000 2458.920 1154.000 2459.070 ;
        RECT -4.800 1759.650 2.400 1760.100 ;
        RECT 15.705 1759.650 16.035 1759.665 ;
        RECT -4.800 1759.350 16.035 1759.650 ;
        RECT -4.800 1758.900 2.400 1759.350 ;
        RECT 15.705 1759.335 16.035 1759.350 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1937.590 738.040 1937.910 738.100 ;
        RECT 2900.830 738.040 2901.150 738.100 ;
        RECT 1937.590 737.900 2901.150 738.040 ;
        RECT 1937.590 737.840 1937.910 737.900 ;
        RECT 2900.830 737.840 2901.150 737.900 ;
      LAYER via ;
        RECT 1937.620 737.840 1937.880 738.100 ;
        RECT 2900.860 737.840 2901.120 738.100 ;
      LAYER met2 ;
        RECT 1937.610 1700.000 1937.890 1704.000 ;
        RECT 1937.680 738.130 1937.820 1700.000 ;
        RECT 1937.620 737.810 1937.880 738.130 ;
        RECT 2900.860 737.810 2901.120 738.130 ;
        RECT 2900.920 733.565 2901.060 737.810 ;
        RECT 2900.850 733.195 2901.130 733.565 ;
      LAYER via2 ;
        RECT 2900.850 733.240 2901.130 733.520 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 732.780 2924.800 733.980 ;
=======
        RECT 2900.825 733.530 2901.155 733.545 ;
        RECT 2917.600 733.530 2924.800 733.980 ;
        RECT 2900.825 733.230 2924.800 733.530 ;
        RECT 2900.825 733.215 2901.155 733.230 ;
        RECT 2917.600 732.780 2924.800 733.230 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1137.650 972.640 1137.970 972.700 ;
        RECT 2900.830 972.640 2901.150 972.700 ;
        RECT 1137.650 972.500 2901.150 972.640 ;
        RECT 1137.650 972.440 1137.970 972.500 ;
        RECT 2900.830 972.440 2901.150 972.500 ;
      LAYER via ;
        RECT 1137.680 972.440 1137.940 972.700 ;
        RECT 2900.860 972.440 2901.120 972.700 ;
      LAYER met2 ;
        RECT 1137.670 1819.155 1137.950 1819.525 ;
        RECT 1137.740 972.730 1137.880 1819.155 ;
        RECT 1137.680 972.410 1137.940 972.730 ;
        RECT 2900.860 972.410 2901.120 972.730 ;
        RECT 2900.920 968.165 2901.060 972.410 ;
        RECT 2900.850 967.795 2901.130 968.165 ;
      LAYER via2 ;
        RECT 1137.670 1819.200 1137.950 1819.480 ;
        RECT 2900.850 967.840 2901.130 968.120 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 967.380 2924.800 968.580 ;
=======
        RECT 1137.645 1819.490 1137.975 1819.505 ;
        RECT 1150.000 1819.490 1154.000 1819.640 ;
        RECT 1137.645 1819.190 1154.000 1819.490 ;
        RECT 1137.645 1819.175 1137.975 1819.190 ;
        RECT 1150.000 1819.040 1154.000 1819.190 ;
        RECT 2900.825 968.130 2901.155 968.145 ;
        RECT 2917.600 968.130 2924.800 968.580 ;
        RECT 2900.825 967.830 2924.800 968.130 ;
        RECT 2900.825 967.815 2901.155 967.830 ;
        RECT 2917.600 967.380 2924.800 967.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1913.210 2511.820 1913.530 2511.880 ;
        RECT 2604.590 2511.820 2604.910 2511.880 ;
        RECT 1913.210 2511.680 2604.910 2511.820 ;
        RECT 1913.210 2511.620 1913.530 2511.680 ;
        RECT 2604.590 2511.620 2604.910 2511.680 ;
        RECT 2604.590 1207.240 2604.910 1207.300 ;
        RECT 2900.830 1207.240 2901.150 1207.300 ;
        RECT 2604.590 1207.100 2901.150 1207.240 ;
        RECT 2604.590 1207.040 2604.910 1207.100 ;
        RECT 2900.830 1207.040 2901.150 1207.100 ;
      LAYER via ;
        RECT 1913.240 2511.620 1913.500 2511.880 ;
        RECT 2604.620 2511.620 2604.880 2511.880 ;
        RECT 2604.620 1207.040 2604.880 1207.300 ;
        RECT 2900.860 1207.040 2901.120 1207.300 ;
      LAYER met2 ;
        RECT 1913.240 2511.590 1913.500 2511.910 ;
        RECT 2604.620 2511.590 2604.880 2511.910 ;
        RECT 1913.300 2500.000 1913.440 2511.590 ;
        RECT 1913.230 2496.000 1913.510 2500.000 ;
        RECT 2604.680 1207.330 2604.820 2511.590 ;
        RECT 2604.620 1207.010 2604.880 1207.330 ;
        RECT 2900.860 1207.010 2901.120 1207.330 ;
        RECT 2900.920 1202.765 2901.060 1207.010 ;
        RECT 2900.850 1202.395 2901.130 1202.765 ;
      LAYER via2 ;
        RECT 2900.850 1202.440 2901.130 1202.720 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1201.980 2924.800 1203.180 ;
=======
        RECT 2900.825 1202.730 2901.155 1202.745 ;
        RECT 2917.600 1202.730 2924.800 1203.180 ;
        RECT 2900.825 1202.430 2924.800 1202.730 ;
        RECT 2900.825 1202.415 2901.155 1202.430 ;
        RECT 2917.600 1201.980 2924.800 1202.430 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1137.190 1441.840 1137.510 1441.900 ;
        RECT 2900.830 1441.840 2901.150 1441.900 ;
        RECT 1137.190 1441.700 2901.150 1441.840 ;
        RECT 1137.190 1441.640 1137.510 1441.700 ;
        RECT 2900.830 1441.640 2901.150 1441.700 ;
      LAYER via ;
        RECT 1137.220 1441.640 1137.480 1441.900 ;
        RECT 2900.860 1441.640 2901.120 1441.900 ;
      LAYER met2 ;
        RECT 1137.210 1899.395 1137.490 1899.765 ;
        RECT 1137.280 1441.930 1137.420 1899.395 ;
        RECT 1137.220 1441.610 1137.480 1441.930 ;
        RECT 2900.860 1441.610 2901.120 1441.930 ;
        RECT 2900.920 1437.365 2901.060 1441.610 ;
        RECT 2900.850 1436.995 2901.130 1437.365 ;
      LAYER via2 ;
        RECT 1137.210 1899.440 1137.490 1899.720 ;
        RECT 2900.850 1437.040 2901.130 1437.320 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1436.580 2924.800 1437.780 ;
=======
        RECT 1137.185 1899.730 1137.515 1899.745 ;
        RECT 1150.000 1899.730 1154.000 1899.880 ;
        RECT 1137.185 1899.430 1154.000 1899.730 ;
        RECT 1137.185 1899.415 1137.515 1899.430 ;
        RECT 1150.000 1899.280 1154.000 1899.430 ;
        RECT 2900.825 1437.330 2901.155 1437.345 ;
        RECT 2917.600 1437.330 2924.800 1437.780 ;
        RECT 2900.825 1437.030 2924.800 1437.330 ;
        RECT 2900.825 1437.015 2901.155 1437.030 ;
        RECT 2917.600 1436.580 2924.800 1437.030 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1938.970 1676.440 1939.290 1676.500 ;
        RECT 2900.830 1676.440 2901.150 1676.500 ;
        RECT 1938.970 1676.300 2901.150 1676.440 ;
        RECT 1938.970 1676.240 1939.290 1676.300 ;
        RECT 2900.830 1676.240 2901.150 1676.300 ;
      LAYER via ;
        RECT 1939.000 1676.240 1939.260 1676.500 ;
        RECT 2900.860 1676.240 2901.120 1676.500 ;
      LAYER met2 ;
        RECT 1938.990 1700.000 1939.270 1704.000 ;
        RECT 1939.060 1676.530 1939.200 1700.000 ;
        RECT 1939.000 1676.210 1939.260 1676.530 ;
        RECT 2900.860 1676.210 2901.120 1676.530 ;
        RECT 2900.920 1671.965 2901.060 1676.210 ;
        RECT 2900.850 1671.595 2901.130 1671.965 ;
      LAYER via2 ;
        RECT 2900.850 1671.640 2901.130 1671.920 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1671.180 2924.800 1672.380 ;
=======
        RECT 2900.825 1671.930 2901.155 1671.945 ;
        RECT 2917.600 1671.930 2924.800 1672.380 ;
        RECT 2900.825 1671.630 2924.800 1671.930 ;
        RECT 2900.825 1671.615 2901.155 1671.630 ;
        RECT 2917.600 1671.180 2924.800 1671.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1905.780 2924.800 1906.980 ;
=======
        RECT 1136.470 1979.290 1136.850 1979.300 ;
        RECT 1150.000 1979.290 1154.000 1979.440 ;
        RECT 1136.470 1978.990 1154.000 1979.290 ;
        RECT 1136.470 1978.980 1136.850 1978.990 ;
        RECT 1150.000 1978.840 1154.000 1978.990 ;
        RECT 2898.270 1906.530 2898.650 1906.540 ;
        RECT 2917.600 1906.530 2924.800 1906.980 ;
        RECT 2898.270 1906.230 2924.800 1906.530 ;
        RECT 2898.270 1906.220 2898.650 1906.230 ;
        RECT 2917.600 1905.780 2924.800 1906.230 ;
      LAYER via3 ;
        RECT 1136.500 1978.980 1136.820 1979.300 ;
        RECT 2898.300 1906.220 2898.620 1906.540 ;
      LAYER met4 ;
        RECT 1136.495 1978.975 1136.825 1979.305 ;
        RECT 1136.510 1906.290 1136.810 1978.975 ;
        RECT 2897.870 1908.510 2899.050 1909.690 ;
        RECT 2898.310 1906.545 2898.610 1908.510 ;
        RECT 1136.070 1905.110 1137.250 1906.290 ;
        RECT 2898.295 1906.215 2898.625 1906.545 ;
      LAYER met5 ;
        RECT 1192.900 1911.700 1269.940 1913.300 ;
        RECT 1192.900 1906.500 1194.500 1911.700 ;
        RECT 1135.860 1904.900 1194.500 1906.500 ;
        RECT 1268.340 1906.500 1269.940 1911.700 ;
        RECT 1289.500 1911.700 1318.700 1913.300 ;
        RECT 1289.500 1906.500 1291.100 1911.700 ;
        RECT 1268.340 1904.900 1291.100 1906.500 ;
        RECT 1317.100 1906.500 1318.700 1911.700 ;
        RECT 1364.020 1911.700 1415.300 1913.300 ;
        RECT 1364.020 1906.500 1365.620 1911.700 ;
        RECT 1317.100 1904.900 1365.620 1906.500 ;
        RECT 1413.700 1906.500 1415.300 1911.700 ;
        RECT 1460.620 1911.700 1511.900 1913.300 ;
        RECT 1460.620 1906.500 1462.220 1911.700 ;
        RECT 1413.700 1904.900 1462.220 1906.500 ;
        RECT 1510.300 1906.500 1511.900 1911.700 ;
        RECT 1557.220 1911.700 1608.500 1913.300 ;
        RECT 1557.220 1906.500 1558.820 1911.700 ;
        RECT 1510.300 1904.900 1558.820 1906.500 ;
        RECT 1606.900 1906.500 1608.500 1911.700 ;
        RECT 1653.820 1911.700 1705.100 1913.300 ;
        RECT 1653.820 1906.500 1655.420 1911.700 ;
        RECT 1606.900 1904.900 1655.420 1906.500 ;
        RECT 1703.500 1906.500 1705.100 1911.700 ;
        RECT 1750.420 1911.700 1801.700 1913.300 ;
        RECT 1750.420 1906.500 1752.020 1911.700 ;
        RECT 1703.500 1904.900 1752.020 1906.500 ;
        RECT 1800.100 1906.500 1801.700 1911.700 ;
        RECT 1847.020 1911.700 1898.300 1913.300 ;
        RECT 1847.020 1906.500 1848.620 1911.700 ;
        RECT 1800.100 1904.900 1848.620 1906.500 ;
        RECT 1896.700 1906.500 1898.300 1911.700 ;
        RECT 1943.620 1911.700 1994.900 1913.300 ;
        RECT 1943.620 1906.500 1945.220 1911.700 ;
        RECT 1896.700 1904.900 1945.220 1906.500 ;
        RECT 1993.300 1906.500 1994.900 1911.700 ;
        RECT 2040.220 1911.700 2091.500 1913.300 ;
        RECT 2040.220 1906.500 2041.820 1911.700 ;
        RECT 1993.300 1904.900 2041.820 1906.500 ;
        RECT 2089.900 1906.500 2091.500 1911.700 ;
        RECT 2136.820 1911.700 2188.100 1913.300 ;
        RECT 2136.820 1906.500 2138.420 1911.700 ;
        RECT 2089.900 1904.900 2138.420 1906.500 ;
        RECT 2186.500 1906.500 2188.100 1911.700 ;
        RECT 2233.420 1911.700 2284.700 1913.300 ;
        RECT 2233.420 1906.500 2235.020 1911.700 ;
        RECT 2186.500 1904.900 2235.020 1906.500 ;
        RECT 2283.100 1906.500 2284.700 1911.700 ;
        RECT 2330.020 1911.700 2381.300 1913.300 ;
        RECT 2330.020 1906.500 2331.620 1911.700 ;
        RECT 2283.100 1904.900 2331.620 1906.500 ;
        RECT 2379.700 1906.500 2381.300 1911.700 ;
        RECT 2426.620 1911.700 2477.900 1913.300 ;
        RECT 2426.620 1906.500 2428.220 1911.700 ;
        RECT 2379.700 1904.900 2428.220 1906.500 ;
        RECT 2476.300 1906.500 2477.900 1911.700 ;
        RECT 2523.220 1911.700 2574.500 1913.300 ;
        RECT 2523.220 1906.500 2524.820 1911.700 ;
        RECT 2476.300 1904.900 2524.820 1906.500 ;
        RECT 2572.900 1906.500 2574.500 1911.700 ;
        RECT 2620.740 1911.700 2740.100 1913.300 ;
        RECT 2620.740 1906.500 2622.340 1911.700 ;
        RECT 2572.900 1904.900 2622.340 1906.500 ;
        RECT 2738.500 1906.500 2740.100 1911.700 ;
        RECT 2766.100 1911.700 2837.620 1913.300 ;
        RECT 2766.100 1906.500 2767.700 1911.700 ;
        RECT 2738.500 1904.900 2767.700 1906.500 ;
        RECT 2836.020 1906.500 2837.620 1911.700 ;
        RECT 2882.940 1911.700 2899.260 1913.300 ;
        RECT 2882.940 1906.500 2884.540 1911.700 ;
        RECT 2897.660 1908.300 2899.260 1911.700 ;
        RECT 2836.020 1904.900 2884.540 1906.500 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1920.110 2512.500 1920.430 2512.560 ;
        RECT 1951.390 2512.500 1951.710 2512.560 ;
        RECT 1920.110 2512.360 1951.710 2512.500 ;
        RECT 1920.110 2512.300 1920.430 2512.360 ;
        RECT 1951.390 2512.300 1951.710 2512.360 ;
        RECT 1951.390 2145.640 1951.710 2145.700 ;
        RECT 2900.830 2145.640 2901.150 2145.700 ;
        RECT 1951.390 2145.500 2901.150 2145.640 ;
        RECT 1951.390 2145.440 1951.710 2145.500 ;
        RECT 2900.830 2145.440 2901.150 2145.500 ;
      LAYER via ;
        RECT 1920.140 2512.300 1920.400 2512.560 ;
        RECT 1951.420 2512.300 1951.680 2512.560 ;
        RECT 1951.420 2145.440 1951.680 2145.700 ;
        RECT 2900.860 2145.440 2901.120 2145.700 ;
      LAYER met2 ;
        RECT 1920.140 2512.270 1920.400 2512.590 ;
        RECT 1951.420 2512.270 1951.680 2512.590 ;
        RECT 1920.200 2500.000 1920.340 2512.270 ;
        RECT 1920.130 2496.000 1920.410 2500.000 ;
        RECT 1951.480 2145.730 1951.620 2512.270 ;
        RECT 1951.420 2145.410 1951.680 2145.730 ;
        RECT 2900.860 2145.410 2901.120 2145.730 ;
        RECT 2900.920 2141.165 2901.060 2145.410 ;
        RECT 2900.850 2140.795 2901.130 2141.165 ;
      LAYER via2 ;
        RECT 2900.850 2140.840 2901.130 2141.120 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2140.380 2924.800 2141.580 ;
=======
        RECT 2900.825 2141.130 2901.155 2141.145 ;
        RECT 2917.600 2141.130 2924.800 2141.580 ;
        RECT 2900.825 2140.830 2924.800 2141.130 ;
        RECT 2900.825 2140.815 2901.155 2140.830 ;
        RECT 2917.600 2140.380 2924.800 2140.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1787.170 84.560 1787.490 84.620 ;
        RECT 1800.970 84.560 1801.290 84.620 ;
        RECT 1787.170 84.420 1801.290 84.560 ;
        RECT 1787.170 84.360 1787.490 84.420 ;
        RECT 1800.970 84.360 1801.290 84.420 ;
        RECT 1593.970 84.220 1594.290 84.280 ;
        RECT 1607.770 84.220 1608.090 84.280 ;
        RECT 1593.970 84.080 1608.090 84.220 ;
        RECT 1593.970 84.020 1594.290 84.080 ;
        RECT 1607.770 84.020 1608.090 84.080 ;
        RECT 1702.070 84.220 1702.390 84.280 ;
        RECT 1704.370 84.220 1704.690 84.280 ;
        RECT 1702.070 84.080 1704.690 84.220 ;
        RECT 1702.070 84.020 1702.390 84.080 ;
        RECT 1704.370 84.020 1704.690 84.080 ;
        RECT 2090.310 84.220 2090.630 84.280 ;
        RECT 2124.810 84.220 2125.130 84.280 ;
        RECT 2090.310 84.080 2125.130 84.220 ;
        RECT 2090.310 84.020 2090.630 84.080 ;
        RECT 2124.810 84.020 2125.130 84.080 ;
        RECT 1932.070 83.540 1932.390 83.600 ;
        RECT 1946.330 83.540 1946.650 83.600 ;
        RECT 1932.070 83.400 1946.650 83.540 ;
        RECT 1932.070 83.340 1932.390 83.400 ;
        RECT 1946.330 83.340 1946.650 83.400 ;
      LAYER via ;
        RECT 1787.200 84.360 1787.460 84.620 ;
        RECT 1801.000 84.360 1801.260 84.620 ;
        RECT 1594.000 84.020 1594.260 84.280 ;
        RECT 1607.800 84.020 1608.060 84.280 ;
        RECT 1702.100 84.020 1702.360 84.280 ;
        RECT 1704.400 84.020 1704.660 84.280 ;
        RECT 2090.340 84.020 2090.600 84.280 ;
        RECT 2124.840 84.020 2125.100 84.280 ;
        RECT 1932.100 83.340 1932.360 83.600 ;
        RECT 1946.360 83.340 1946.620 83.600 ;
      LAYER met2 ;
        RECT 1153.310 2498.050 1153.590 2500.000 ;
        RECT 1155.150 2498.050 1155.430 2498.165 ;
        RECT 1153.310 2497.910 1155.430 2498.050 ;
        RECT 1153.310 2496.000 1153.590 2497.910 ;
        RECT 1155.150 2497.795 1155.430 2497.910 ;
        RECT 1907.710 86.515 1907.990 86.885 ;
        RECT 1787.190 84.475 1787.470 84.845 ;
        RECT 1800.990 84.475 1801.270 84.845 ;
        RECT 1787.200 84.330 1787.460 84.475 ;
        RECT 1801.000 84.330 1801.260 84.475 ;
        RECT 1594.000 84.165 1594.260 84.310 ;
        RECT 1607.800 84.165 1608.060 84.310 ;
        RECT 1702.100 84.165 1702.360 84.310 ;
        RECT 1704.400 84.165 1704.660 84.310 ;
        RECT 1593.990 83.795 1594.270 84.165 ;
        RECT 1607.790 83.795 1608.070 84.165 ;
        RECT 1702.090 83.795 1702.370 84.165 ;
        RECT 1704.390 83.795 1704.670 84.165 ;
        RECT 1907.780 83.485 1907.920 86.515 ;
        RECT 2028.230 85.835 2028.510 86.205 ;
        RECT 1946.350 84.475 1946.630 84.845 ;
        RECT 1946.420 83.630 1946.560 84.475 ;
        RECT 2028.300 84.165 2028.440 85.835 ;
        RECT 2124.830 84.475 2125.110 84.845 ;
        RECT 2124.900 84.310 2125.040 84.475 ;
        RECT 2090.340 84.165 2090.600 84.310 ;
        RECT 2028.230 83.795 2028.510 84.165 ;
        RECT 2042.030 83.795 2042.310 84.165 ;
        RECT 2090.330 83.795 2090.610 84.165 ;
        RECT 2124.840 83.990 2125.100 84.310 ;
        RECT 1932.100 83.485 1932.360 83.630 ;
        RECT 1907.710 83.115 1907.990 83.485 ;
        RECT 1932.090 83.115 1932.370 83.485 ;
        RECT 1946.360 83.310 1946.620 83.630 ;
        RECT 2042.100 83.370 2042.240 83.795 ;
        RECT 2042.950 83.370 2043.230 83.485 ;
        RECT 2042.100 83.230 2043.230 83.370 ;
        RECT 2042.950 83.115 2043.230 83.230 ;
      LAYER via2 ;
        RECT 1155.150 2497.840 1155.430 2498.120 ;
        RECT 1907.710 86.560 1907.990 86.840 ;
        RECT 1787.190 84.520 1787.470 84.800 ;
        RECT 1800.990 84.520 1801.270 84.800 ;
        RECT 1593.990 83.840 1594.270 84.120 ;
        RECT 1607.790 83.840 1608.070 84.120 ;
        RECT 1702.090 83.840 1702.370 84.120 ;
        RECT 1704.390 83.840 1704.670 84.120 ;
        RECT 2028.230 85.880 2028.510 86.160 ;
        RECT 1946.350 84.520 1946.630 84.800 ;
        RECT 2124.830 84.520 2125.110 84.800 ;
        RECT 2028.230 83.840 2028.510 84.120 ;
        RECT 2042.030 83.840 2042.310 84.120 ;
        RECT 2090.330 83.840 2090.610 84.120 ;
        RECT 1907.710 83.160 1907.990 83.440 ;
        RECT 1932.090 83.160 1932.370 83.440 ;
        RECT 2042.950 83.160 2043.230 83.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 87.460 2924.800 88.660 ;
=======
        RECT 1155.125 2498.130 1155.455 2498.145 ;
        RECT 1158.550 2498.130 1158.930 2498.140 ;
        RECT 1155.125 2497.830 1158.930 2498.130 ;
        RECT 1155.125 2497.815 1155.455 2497.830 ;
        RECT 1158.550 2497.820 1158.930 2497.830 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2916.710 87.910 2924.800 88.210 ;
        RECT 1883.510 86.850 1883.890 86.860 ;
        RECT 1907.685 86.850 1908.015 86.865 ;
        RECT 1883.510 86.550 1908.015 86.850 ;
        RECT 1883.510 86.540 1883.890 86.550 ;
        RECT 1907.685 86.535 1908.015 86.550 ;
        RECT 1980.110 86.170 1980.490 86.180 ;
        RECT 2028.205 86.170 2028.535 86.185 ;
        RECT 1980.110 85.870 2028.535 86.170 ;
        RECT 1980.110 85.860 1980.490 85.870 ;
        RECT 2028.205 85.855 2028.535 85.870 ;
        RECT 1883.510 85.490 1883.890 85.500 ;
        RECT 1873.430 85.190 1883.890 85.490 ;
        RECT 1787.165 84.810 1787.495 84.825 ;
        RECT 1752.910 84.510 1787.495 84.810 ;
        RECT 1593.965 84.130 1594.295 84.145 ;
        RECT 1559.710 83.830 1594.295 84.130 ;
        RECT 1158.550 83.450 1158.930 83.460 ;
        RECT 1559.710 83.450 1560.010 83.830 ;
        RECT 1593.965 83.815 1594.295 83.830 ;
        RECT 1607.765 84.130 1608.095 84.145 ;
        RECT 1702.065 84.130 1702.395 84.145 ;
        RECT 1607.765 83.830 1641.890 84.130 ;
        RECT 1607.765 83.815 1608.095 83.830 ;
        RECT 1158.550 83.150 1560.010 83.450 ;
        RECT 1641.590 83.450 1641.890 83.830 ;
        RECT 1656.310 83.830 1702.395 84.130 ;
        RECT 1656.310 83.450 1656.610 83.830 ;
        RECT 1702.065 83.815 1702.395 83.830 ;
        RECT 1704.365 84.130 1704.695 84.145 ;
        RECT 1704.365 83.830 1738.490 84.130 ;
        RECT 1704.365 83.815 1704.695 83.830 ;
        RECT 1641.590 83.150 1656.610 83.450 ;
        RECT 1738.190 83.450 1738.490 83.830 ;
        RECT 1752.910 83.450 1753.210 84.510 ;
        RECT 1787.165 84.495 1787.495 84.510 ;
        RECT 1800.965 84.810 1801.295 84.825 ;
        RECT 1800.965 84.510 1835.090 84.810 ;
        RECT 1800.965 84.495 1801.295 84.510 ;
        RECT 1834.790 84.130 1835.090 84.510 ;
        RECT 1873.430 84.130 1873.730 85.190 ;
        RECT 1883.510 85.180 1883.890 85.190 ;
        RECT 1946.325 84.810 1946.655 84.825 ;
        RECT 1980.110 84.810 1980.490 84.820 ;
        RECT 1946.325 84.510 1980.490 84.810 ;
        RECT 1946.325 84.495 1946.655 84.510 ;
        RECT 1980.110 84.500 1980.490 84.510 ;
        RECT 2124.805 84.810 2125.135 84.825 ;
        RECT 2124.805 84.510 2159.850 84.810 ;
        RECT 2124.805 84.495 2125.135 84.510 ;
        RECT 1834.790 83.830 1873.730 84.130 ;
        RECT 2028.205 84.130 2028.535 84.145 ;
        RECT 2042.005 84.130 2042.335 84.145 ;
        RECT 2090.305 84.130 2090.635 84.145 ;
        RECT 2028.205 83.830 2042.335 84.130 ;
        RECT 2028.205 83.815 2028.535 83.830 ;
        RECT 2042.005 83.815 2042.335 83.830 ;
        RECT 2076.750 83.830 2090.635 84.130 ;
        RECT 2159.550 84.130 2159.850 84.510 ;
        RECT 2208.310 84.510 2256.450 84.810 ;
        RECT 2159.550 83.830 2207.690 84.130 ;
        RECT 1738.190 83.150 1753.210 83.450 ;
        RECT 1907.685 83.450 1908.015 83.465 ;
        RECT 1932.065 83.450 1932.395 83.465 ;
        RECT 1907.685 83.150 1932.395 83.450 ;
        RECT 1158.550 83.140 1158.930 83.150 ;
        RECT 1907.685 83.135 1908.015 83.150 ;
        RECT 1932.065 83.135 1932.395 83.150 ;
        RECT 2042.925 83.450 2043.255 83.465 ;
        RECT 2076.750 83.450 2077.050 83.830 ;
        RECT 2090.305 83.815 2090.635 83.830 ;
        RECT 2042.925 83.150 2077.050 83.450 ;
        RECT 2207.390 83.450 2207.690 83.830 ;
        RECT 2208.310 83.450 2208.610 84.510 ;
        RECT 2256.150 84.130 2256.450 84.510 ;
        RECT 2304.910 84.510 2353.050 84.810 ;
        RECT 2256.150 83.830 2304.290 84.130 ;
        RECT 2207.390 83.150 2208.610 83.450 ;
        RECT 2303.990 83.450 2304.290 83.830 ;
        RECT 2304.910 83.450 2305.210 84.510 ;
        RECT 2352.750 84.130 2353.050 84.510 ;
        RECT 2401.510 84.510 2449.650 84.810 ;
        RECT 2352.750 83.830 2400.890 84.130 ;
        RECT 2303.990 83.150 2305.210 83.450 ;
        RECT 2400.590 83.450 2400.890 83.830 ;
        RECT 2401.510 83.450 2401.810 84.510 ;
        RECT 2449.350 84.130 2449.650 84.510 ;
        RECT 2498.110 84.510 2546.250 84.810 ;
        RECT 2449.350 83.830 2497.490 84.130 ;
        RECT 2400.590 83.150 2401.810 83.450 ;
        RECT 2497.190 83.450 2497.490 83.830 ;
        RECT 2498.110 83.450 2498.410 84.510 ;
        RECT 2545.950 84.130 2546.250 84.510 ;
        RECT 2594.710 84.510 2642.850 84.810 ;
        RECT 2545.950 83.830 2594.090 84.130 ;
        RECT 2497.190 83.150 2498.410 83.450 ;
        RECT 2593.790 83.450 2594.090 83.830 ;
        RECT 2594.710 83.450 2595.010 84.510 ;
        RECT 2642.550 84.130 2642.850 84.510 ;
        RECT 2691.310 84.510 2739.450 84.810 ;
        RECT 2642.550 83.830 2690.690 84.130 ;
        RECT 2593.790 83.150 2595.010 83.450 ;
        RECT 2690.390 83.450 2690.690 83.830 ;
        RECT 2691.310 83.450 2691.610 84.510 ;
        RECT 2739.150 84.130 2739.450 84.510 ;
        RECT 2787.910 84.510 2836.050 84.810 ;
        RECT 2739.150 83.830 2787.290 84.130 ;
        RECT 2690.390 83.150 2691.610 83.450 ;
        RECT 2786.990 83.450 2787.290 83.830 ;
        RECT 2787.910 83.450 2788.210 84.510 ;
        RECT 2835.750 84.130 2836.050 84.510 ;
        RECT 2916.710 84.130 2917.010 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
        RECT 2835.750 83.830 2883.890 84.130 ;
        RECT 2786.990 83.150 2788.210 83.450 ;
        RECT 2883.590 83.450 2883.890 83.830 ;
        RECT 2884.510 83.830 2917.010 84.130 ;
        RECT 2884.510 83.450 2884.810 83.830 ;
        RECT 2883.590 83.150 2884.810 83.450 ;
        RECT 2042.925 83.135 2043.255 83.150 ;
      LAYER via3 ;
        RECT 1158.580 2497.820 1158.900 2498.140 ;
        RECT 1883.540 86.540 1883.860 86.860 ;
        RECT 1980.140 85.860 1980.460 86.180 ;
        RECT 1158.580 83.140 1158.900 83.460 ;
        RECT 1883.540 85.180 1883.860 85.500 ;
        RECT 1980.140 84.500 1980.460 84.820 ;
      LAYER met4 ;
        RECT 1158.575 2497.815 1158.905 2498.145 ;
        RECT 1158.590 83.465 1158.890 2497.815 ;
        RECT 1883.535 86.535 1883.865 86.865 ;
        RECT 1883.550 85.505 1883.850 86.535 ;
        RECT 1980.135 85.855 1980.465 86.185 ;
        RECT 1883.535 85.175 1883.865 85.505 ;
        RECT 1980.150 84.825 1980.450 85.855 ;
        RECT 1980.135 84.495 1980.465 84.825 ;
        RECT 1158.575 83.135 1158.905 83.465 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1352.085 2495.685 1352.255 2497.215 ;
      LAYER mcon ;
        RECT 1352.085 2497.045 1352.255 2497.215 ;
      LAYER met1 ;
        RECT 1352.010 2497.200 1352.330 2497.260 ;
        RECT 1351.815 2497.060 1352.330 2497.200 ;
        RECT 1352.010 2497.000 1352.330 2497.060 ;
        RECT 1352.025 2495.840 1352.315 2495.885 ;
        RECT 2901.750 2495.840 2902.070 2495.900 ;
        RECT 1352.025 2495.700 2902.070 2495.840 ;
        RECT 1352.025 2495.655 1352.315 2495.700 ;
        RECT 2901.750 2495.640 2902.070 2495.700 ;
      LAYER via ;
        RECT 1352.040 2497.000 1352.300 2497.260 ;
        RECT 2901.780 2495.640 2902.040 2495.900 ;
      LAYER met2 ;
        RECT 1351.570 2497.370 1351.850 2500.000 ;
        RECT 1351.570 2497.290 1352.240 2497.370 ;
        RECT 1351.570 2497.230 1352.300 2497.290 ;
        RECT 1351.570 2496.000 1351.850 2497.230 ;
        RECT 1352.040 2496.970 1352.300 2497.230 ;
        RECT 2901.780 2495.610 2902.040 2495.930 ;
        RECT 2901.840 2434.245 2901.980 2495.610 ;
        RECT 2901.770 2433.875 2902.050 2434.245 ;
      LAYER via2 ;
        RECT 2901.770 2433.920 2902.050 2434.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2433.460 2924.800 2434.660 ;
=======
        RECT 2901.745 2434.210 2902.075 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2901.745 2433.910 2924.800 2434.210 ;
        RECT 2901.745 2433.895 2902.075 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1372.710 2663.800 1373.030 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 1372.710 2663.660 2901.150 2663.800 ;
        RECT 1372.710 2663.600 1373.030 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
      LAYER via ;
        RECT 1372.740 2663.600 1373.000 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 1372.740 2663.570 1373.000 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 1371.350 2499.410 1371.630 2500.000 ;
        RECT 1372.800 2499.410 1372.940 2663.570 ;
        RECT 1371.350 2499.270 1372.940 2499.410 ;
        RECT 1371.350 2496.000 1371.630 2499.270 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2668.740 2924.800 2669.940 ;
=======
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1393.410 2898.400 1393.730 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 1393.410 2898.260 2901.150 2898.400 ;
        RECT 1393.410 2898.200 1393.730 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
      LAYER via ;
        RECT 1393.440 2898.200 1393.700 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 1393.440 2898.170 1393.700 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 1391.130 2498.730 1391.410 2500.000 ;
        RECT 1393.500 2498.730 1393.640 2898.170 ;
        RECT 1391.130 2498.590 1393.640 2498.730 ;
        RECT 1391.130 2496.000 1391.410 2498.590 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2903.340 2924.800 2904.540 ;
=======
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1414.110 3133.000 1414.430 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 1414.110 3132.860 2901.150 3133.000 ;
        RECT 1414.110 3132.800 1414.430 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 1414.140 3132.800 1414.400 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 1414.140 3132.770 1414.400 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 1410.910 2498.730 1411.190 2500.000 ;
        RECT 1414.200 2499.410 1414.340 3132.770 ;
        RECT 1413.740 2499.270 1414.340 2499.410 ;
        RECT 1413.740 2498.730 1413.880 2499.270 ;
        RECT 1410.910 2498.590 1413.880 2498.730 ;
        RECT 1410.910 2496.000 1411.190 2498.590 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3137.940 2924.800 3139.140 ;
=======
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1434.810 3367.600 1435.130 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1434.810 3367.460 2901.150 3367.600 ;
        RECT 1434.810 3367.400 1435.130 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 1430.670 2514.880 1430.990 2514.940 ;
        RECT 1434.810 2514.880 1435.130 2514.940 ;
        RECT 1430.670 2514.740 1435.130 2514.880 ;
        RECT 1430.670 2514.680 1430.990 2514.740 ;
        RECT 1434.810 2514.680 1435.130 2514.740 ;
      LAYER via ;
        RECT 1434.840 3367.400 1435.100 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 1430.700 2514.680 1430.960 2514.940 ;
        RECT 1434.840 2514.680 1435.100 2514.940 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1434.840 3367.370 1435.100 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1434.900 2514.970 1435.040 3367.370 ;
        RECT 1430.700 2514.650 1430.960 2514.970 ;
        RECT 1434.840 2514.650 1435.100 2514.970 ;
        RECT 1430.760 2500.000 1430.900 2514.650 ;
        RECT 1430.690 2496.000 1430.970 2500.000 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3372.540 2924.800 3373.740 ;
=======
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1455.510 3501.900 1455.830 3501.960 ;
        RECT 2798.250 3501.900 2798.570 3501.960 ;
        RECT 1455.510 3501.760 2798.570 3501.900 ;
        RECT 1455.510 3501.700 1455.830 3501.760 ;
        RECT 2798.250 3501.700 2798.570 3501.760 ;
        RECT 1450.450 2514.880 1450.770 2514.940 ;
        RECT 1455.510 2514.880 1455.830 2514.940 ;
        RECT 1450.450 2514.740 1455.830 2514.880 ;
        RECT 1450.450 2514.680 1450.770 2514.740 ;
        RECT 1455.510 2514.680 1455.830 2514.740 ;
      LAYER via ;
        RECT 1455.540 3501.700 1455.800 3501.960 ;
        RECT 2798.280 3501.700 2798.540 3501.960 ;
        RECT 1450.480 2514.680 1450.740 2514.940 ;
        RECT 1455.540 2514.680 1455.800 2514.940 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2798.130 3519.700 2798.690 3524.800 ;
=======
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.990 2798.480 3517.600 ;
        RECT 1455.540 3501.670 1455.800 3501.990 ;
        RECT 2798.280 3501.670 2798.540 3501.990 ;
        RECT 1455.600 2514.970 1455.740 3501.670 ;
        RECT 1450.480 2514.650 1450.740 2514.970 ;
        RECT 1455.540 2514.650 1455.800 2514.970 ;
        RECT 1450.540 2500.000 1450.680 2514.650 ;
        RECT 1450.470 2496.000 1450.750 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1476.210 3503.600 1476.530 3503.660 ;
        RECT 2473.950 3503.600 2474.270 3503.660 ;
        RECT 1476.210 3503.460 2474.270 3503.600 ;
        RECT 1476.210 3503.400 1476.530 3503.460 ;
        RECT 2473.950 3503.400 2474.270 3503.460 ;
        RECT 1470.230 2514.880 1470.550 2514.940 ;
        RECT 1476.210 2514.880 1476.530 2514.940 ;
        RECT 1470.230 2514.740 1476.530 2514.880 ;
        RECT 1470.230 2514.680 1470.550 2514.740 ;
        RECT 1476.210 2514.680 1476.530 2514.740 ;
      LAYER via ;
        RECT 1476.240 3503.400 1476.500 3503.660 ;
        RECT 2473.980 3503.400 2474.240 3503.660 ;
        RECT 1470.260 2514.680 1470.520 2514.940 ;
        RECT 1476.240 2514.680 1476.500 2514.940 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2473.830 3519.700 2474.390 3524.800 ;
=======
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3503.690 2474.180 3517.600 ;
        RECT 1476.240 3503.370 1476.500 3503.690 ;
        RECT 2473.980 3503.370 2474.240 3503.690 ;
        RECT 1476.300 2514.970 1476.440 3503.370 ;
        RECT 1470.260 2514.650 1470.520 2514.970 ;
        RECT 1476.240 2514.650 1476.500 2514.970 ;
        RECT 1470.320 2500.000 1470.460 2514.650 ;
        RECT 1470.250 2496.000 1470.530 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3422.355 ;
        RECT 2147.425 3139.645 2147.595 3187.755 ;
        RECT 2146.965 3088.645 2147.135 3132.675 ;
        RECT 2147.885 2946.525 2148.055 3035.775 ;
        RECT 2146.505 2753.065 2146.675 2801.175 ;
      LAYER mcon ;
        RECT 2147.885 3422.185 2148.055 3422.355 ;
        RECT 2147.425 3187.585 2147.595 3187.755 ;
        RECT 2146.965 3132.505 2147.135 3132.675 ;
        RECT 2147.885 3035.605 2148.055 3035.775 ;
        RECT 2146.505 2801.005 2146.675 2801.175 ;
      LAYER met1 ;
        RECT 2146.890 3443.080 2147.210 3443.140 ;
        RECT 2149.190 3443.080 2149.510 3443.140 ;
        RECT 2146.890 3442.940 2149.510 3443.080 ;
        RECT 2146.890 3442.880 2147.210 3442.940 ;
        RECT 2149.190 3442.880 2149.510 3442.940 ;
        RECT 2146.430 3422.340 2146.750 3422.400 ;
        RECT 2147.825 3422.340 2148.115 3422.385 ;
        RECT 2146.430 3422.200 2148.115 3422.340 ;
        RECT 2146.430 3422.140 2146.750 3422.200 ;
        RECT 2147.825 3422.155 2148.115 3422.200 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2147.350 3187.740 2147.670 3187.800 ;
        RECT 2147.155 3187.600 2147.670 3187.740 ;
        RECT 2147.350 3187.540 2147.670 3187.600 ;
        RECT 2147.365 3139.800 2147.655 3139.845 ;
        RECT 2147.810 3139.800 2148.130 3139.860 ;
        RECT 2147.365 3139.660 2148.130 3139.800 ;
        RECT 2147.365 3139.615 2147.655 3139.660 ;
        RECT 2147.810 3139.600 2148.130 3139.660 ;
        RECT 2146.905 3132.660 2147.195 3132.705 ;
        RECT 2147.810 3132.660 2148.130 3132.720 ;
        RECT 2146.905 3132.520 2148.130 3132.660 ;
        RECT 2146.905 3132.475 2147.195 3132.520 ;
        RECT 2147.810 3132.460 2148.130 3132.520 ;
        RECT 2146.890 3088.800 2147.210 3088.860 ;
        RECT 2146.695 3088.660 2147.210 3088.800 ;
        RECT 2146.890 3088.600 2147.210 3088.660 ;
        RECT 2147.350 3036.440 2147.670 3036.500 ;
        RECT 2147.810 3036.440 2148.130 3036.500 ;
        RECT 2147.350 3036.300 2148.130 3036.440 ;
        RECT 2147.350 3036.240 2147.670 3036.300 ;
        RECT 2147.810 3036.240 2148.130 3036.300 ;
        RECT 2147.810 3035.760 2148.130 3035.820 ;
        RECT 2147.615 3035.620 2148.130 3035.760 ;
        RECT 2147.810 3035.560 2148.130 3035.620 ;
        RECT 2147.825 2946.680 2148.115 2946.725 ;
        RECT 2148.270 2946.680 2148.590 2946.740 ;
        RECT 2147.825 2946.540 2148.590 2946.680 ;
        RECT 2147.825 2946.495 2148.115 2946.540 ;
        RECT 2148.270 2946.480 2148.590 2946.540 ;
        RECT 2148.270 2912.340 2148.590 2912.400 ;
        RECT 2147.900 2912.200 2148.590 2912.340 ;
        RECT 2147.900 2911.720 2148.040 2912.200 ;
        RECT 2148.270 2912.140 2148.590 2912.200 ;
        RECT 2147.810 2911.460 2148.130 2911.720 ;
        RECT 2146.430 2815.580 2146.750 2815.840 ;
        RECT 2146.520 2815.160 2146.660 2815.580 ;
        RECT 2146.430 2814.900 2146.750 2815.160 ;
        RECT 2146.430 2801.160 2146.750 2801.220 ;
        RECT 2146.235 2801.020 2146.750 2801.160 ;
        RECT 2146.430 2800.960 2146.750 2801.020 ;
        RECT 2146.445 2753.220 2146.735 2753.265 ;
        RECT 2147.350 2753.220 2147.670 2753.280 ;
        RECT 2146.445 2753.080 2147.670 2753.220 ;
        RECT 2146.445 2753.035 2146.735 2753.080 ;
        RECT 2147.350 2753.020 2147.670 2753.080 ;
        RECT 2146.430 2718.200 2146.750 2718.260 ;
        RECT 2147.350 2718.200 2147.670 2718.260 ;
        RECT 2146.430 2718.060 2147.670 2718.200 ;
        RECT 2146.430 2718.000 2146.750 2718.060 ;
        RECT 2147.350 2718.000 2147.670 2718.060 ;
        RECT 2146.430 2670.260 2146.750 2670.320 ;
        RECT 2147.350 2670.260 2147.670 2670.320 ;
        RECT 2146.430 2670.120 2147.670 2670.260 ;
        RECT 2146.430 2670.060 2146.750 2670.120 ;
        RECT 2147.350 2670.060 2147.670 2670.120 ;
        RECT 2147.350 2622.120 2147.670 2622.380 ;
        RECT 2147.440 2621.980 2147.580 2622.120 ;
        RECT 2147.810 2621.980 2148.130 2622.040 ;
        RECT 2147.440 2621.840 2148.130 2621.980 ;
        RECT 2147.810 2621.780 2148.130 2621.840 ;
        RECT 2146.890 2560.100 2147.210 2560.160 ;
        RECT 2148.270 2560.100 2148.590 2560.160 ;
        RECT 2146.890 2559.960 2148.590 2560.100 ;
        RECT 2146.890 2559.900 2147.210 2559.960 ;
        RECT 2148.270 2559.900 2148.590 2559.960 ;
        RECT 1490.010 2522.360 1490.330 2522.420 ;
        RECT 2148.270 2522.360 2148.590 2522.420 ;
        RECT 1490.010 2522.220 2148.590 2522.360 ;
        RECT 1490.010 2522.160 1490.330 2522.220 ;
        RECT 2148.270 2522.160 2148.590 2522.220 ;
      LAYER via ;
        RECT 2146.920 3442.880 2147.180 3443.140 ;
        RECT 2149.220 3442.880 2149.480 3443.140 ;
        RECT 2146.460 3422.140 2146.720 3422.400 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2147.380 3187.540 2147.640 3187.800 ;
        RECT 2147.840 3139.600 2148.100 3139.860 ;
        RECT 2147.840 3132.460 2148.100 3132.720 ;
        RECT 2146.920 3088.600 2147.180 3088.860 ;
        RECT 2147.380 3036.240 2147.640 3036.500 ;
        RECT 2147.840 3036.240 2148.100 3036.500 ;
        RECT 2147.840 3035.560 2148.100 3035.820 ;
        RECT 2148.300 2946.480 2148.560 2946.740 ;
        RECT 2148.300 2912.140 2148.560 2912.400 ;
        RECT 2147.840 2911.460 2148.100 2911.720 ;
        RECT 2146.460 2815.580 2146.720 2815.840 ;
        RECT 2146.460 2814.900 2146.720 2815.160 ;
        RECT 2146.460 2800.960 2146.720 2801.220 ;
        RECT 2147.380 2753.020 2147.640 2753.280 ;
        RECT 2146.460 2718.000 2146.720 2718.260 ;
        RECT 2147.380 2718.000 2147.640 2718.260 ;
        RECT 2146.460 2670.060 2146.720 2670.320 ;
        RECT 2147.380 2670.060 2147.640 2670.320 ;
        RECT 2147.380 2622.120 2147.640 2622.380 ;
        RECT 2147.840 2621.780 2148.100 2622.040 ;
        RECT 2146.920 2559.900 2147.180 2560.160 ;
        RECT 2148.300 2559.900 2148.560 2560.160 ;
        RECT 1490.040 2522.160 1490.300 2522.420 ;
        RECT 2148.300 2522.160 2148.560 2522.420 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2149.070 3519.700 2149.630 3524.800 ;
=======
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3443.170 2149.420 3517.600 ;
        RECT 2146.920 3442.850 2147.180 3443.170 ;
        RECT 2149.220 3442.850 2149.480 3443.170 ;
        RECT 2146.980 3429.650 2147.120 3442.850 ;
        RECT 2146.520 3429.510 2147.120 3429.650 ;
        RECT 2146.520 3422.430 2146.660 3429.510 ;
        RECT 2146.460 3422.110 2146.720 3422.430 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3236.450 2147.580 3298.270 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3201.850 2147.120 3236.130 ;
        RECT 2146.980 3201.710 2147.580 3201.850 ;
        RECT 2147.440 3187.830 2147.580 3201.710 ;
        RECT 2147.380 3187.510 2147.640 3187.830 ;
        RECT 2147.840 3139.570 2148.100 3139.890 ;
        RECT 2147.900 3132.750 2148.040 3139.570 ;
        RECT 2147.840 3132.430 2148.100 3132.750 ;
        RECT 2146.920 3088.570 2147.180 3088.890 ;
        RECT 2146.980 3084.325 2147.120 3088.570 ;
        RECT 2146.910 3083.955 2147.190 3084.325 ;
        RECT 2147.830 3083.955 2148.110 3084.325 ;
        RECT 2147.900 3036.530 2148.040 3083.955 ;
        RECT 2147.380 3036.210 2147.640 3036.530 ;
        RECT 2147.840 3036.210 2148.100 3036.530 ;
        RECT 2147.440 3035.930 2147.580 3036.210 ;
        RECT 2147.440 3035.850 2148.040 3035.930 ;
        RECT 2147.440 3035.790 2148.100 3035.850 ;
        RECT 2147.840 3035.530 2148.100 3035.790 ;
        RECT 2148.300 2946.450 2148.560 2946.770 ;
        RECT 2148.360 2912.430 2148.500 2946.450 ;
        RECT 2148.300 2912.110 2148.560 2912.430 ;
        RECT 2147.840 2911.430 2148.100 2911.750 ;
        RECT 2147.900 2863.210 2148.040 2911.430 ;
        RECT 2146.980 2863.070 2148.040 2863.210 ;
        RECT 2146.980 2849.610 2147.120 2863.070 ;
        RECT 2146.520 2849.470 2147.120 2849.610 ;
        RECT 2146.520 2815.870 2146.660 2849.470 ;
        RECT 2146.460 2815.550 2146.720 2815.870 ;
        RECT 2146.460 2814.870 2146.720 2815.190 ;
        RECT 2146.520 2801.250 2146.660 2814.870 ;
        RECT 2146.460 2800.930 2146.720 2801.250 ;
        RECT 2147.380 2752.990 2147.640 2753.310 ;
        RECT 2147.440 2718.290 2147.580 2752.990 ;
        RECT 2146.460 2717.970 2146.720 2718.290 ;
        RECT 2147.380 2717.970 2147.640 2718.290 ;
        RECT 2146.520 2670.350 2146.660 2717.970 ;
        RECT 2146.460 2670.030 2146.720 2670.350 ;
        RECT 2147.380 2670.030 2147.640 2670.350 ;
        RECT 2147.440 2622.410 2147.580 2670.030 ;
        RECT 2147.380 2622.090 2147.640 2622.410 ;
        RECT 2147.840 2621.750 2148.100 2622.070 ;
        RECT 2147.900 2608.325 2148.040 2621.750 ;
        RECT 2146.910 2607.955 2147.190 2608.325 ;
        RECT 2147.830 2607.955 2148.110 2608.325 ;
        RECT 2146.980 2560.190 2147.120 2607.955 ;
        RECT 2146.920 2559.870 2147.180 2560.190 ;
        RECT 2148.300 2559.870 2148.560 2560.190 ;
        RECT 2148.360 2522.450 2148.500 2559.870 ;
        RECT 1490.040 2522.130 1490.300 2522.450 ;
        RECT 2148.300 2522.130 2148.560 2522.450 ;
        RECT 1490.100 2500.000 1490.240 2522.130 ;
        RECT 1490.030 2496.000 1490.310 2500.000 ;
      LAYER via2 ;
        RECT 2146.910 3084.000 2147.190 3084.280 ;
        RECT 2147.830 3084.000 2148.110 3084.280 ;
        RECT 2146.910 2608.000 2147.190 2608.280 ;
        RECT 2147.830 2608.000 2148.110 2608.280 ;
      LAYER met3 ;
        RECT 2146.885 3084.290 2147.215 3084.305 ;
        RECT 2147.805 3084.290 2148.135 3084.305 ;
        RECT 2146.885 3083.990 2148.135 3084.290 ;
        RECT 2146.885 3083.975 2147.215 3083.990 ;
        RECT 2147.805 3083.975 2148.135 3083.990 ;
        RECT 2146.885 2608.290 2147.215 2608.305 ;
        RECT 2147.805 2608.290 2148.135 2608.305 ;
        RECT 2146.885 2607.990 2148.135 2608.290 ;
        RECT 2146.885 2607.975 2147.215 2607.990 ;
        RECT 2147.805 2607.975 2148.135 2607.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1510.710 3499.860 1511.030 3499.920 ;
        RECT 1824.890 3499.860 1825.210 3499.920 ;
        RECT 1510.710 3499.720 1825.210 3499.860 ;
        RECT 1510.710 3499.660 1511.030 3499.720 ;
        RECT 1824.890 3499.660 1825.210 3499.720 ;
      LAYER via ;
        RECT 1510.740 3499.660 1511.000 3499.920 ;
        RECT 1824.920 3499.660 1825.180 3499.920 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1824.770 3519.700 1825.330 3524.800 ;
=======
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3499.950 1825.120 3517.600 ;
        RECT 1510.740 3499.630 1511.000 3499.950 ;
        RECT 1824.920 3499.630 1825.180 3499.950 ;
        RECT 1510.270 2499.410 1510.550 2500.000 ;
        RECT 1510.800 2499.410 1510.940 3499.630 ;
        RECT 1510.270 2499.270 1510.940 2499.410 ;
        RECT 1510.270 2496.000 1510.550 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3499.180 1500.910 3499.240 ;
        RECT 1524.970 3499.180 1525.290 3499.240 ;
        RECT 1500.590 3499.040 1525.290 3499.180 ;
        RECT 1500.590 3498.980 1500.910 3499.040 ;
        RECT 1524.970 3498.980 1525.290 3499.040 ;
      LAYER via ;
        RECT 1500.620 3498.980 1500.880 3499.240 ;
        RECT 1525.000 3498.980 1525.260 3499.240 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1500.470 3519.700 1501.030 3524.800 ;
=======
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3499.270 1500.820 3517.600 ;
        RECT 1500.620 3498.950 1500.880 3499.270 ;
        RECT 1525.000 3498.950 1525.260 3499.270 ;
        RECT 1525.060 2498.730 1525.200 3498.950 ;
        RECT 1530.050 2498.730 1530.330 2500.000 ;
        RECT 1525.060 2498.590 1530.330 2498.730 ;
        RECT 1530.050 2496.000 1530.330 2498.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1587.070 319.160 1587.390 319.220 ;
        RECT 1608.230 319.160 1608.550 319.220 ;
        RECT 1587.070 319.020 1608.550 319.160 ;
        RECT 1587.070 318.960 1587.390 319.020 ;
        RECT 1608.230 318.960 1608.550 319.020 ;
        RECT 1702.070 318.820 1702.390 318.880 ;
        RECT 1704.370 318.820 1704.690 318.880 ;
        RECT 1702.070 318.680 1704.690 318.820 ;
        RECT 1702.070 318.620 1702.390 318.680 ;
        RECT 1704.370 318.620 1704.690 318.680 ;
        RECT 1798.670 318.820 1798.990 318.880 ;
        RECT 1801.890 318.820 1802.210 318.880 ;
        RECT 1798.670 318.680 1802.210 318.820 ;
        RECT 1798.670 318.620 1798.990 318.680 ;
        RECT 1801.890 318.620 1802.210 318.680 ;
        RECT 2090.310 318.820 2090.630 318.880 ;
        RECT 2124.810 318.820 2125.130 318.880 ;
        RECT 2090.310 318.680 2125.130 318.820 ;
        RECT 2090.310 318.620 2090.630 318.680 ;
        RECT 2124.810 318.620 2125.130 318.680 ;
        RECT 1932.070 318.140 1932.390 318.200 ;
        RECT 1946.330 318.140 1946.650 318.200 ;
        RECT 1932.070 318.000 1946.650 318.140 ;
        RECT 1932.070 317.940 1932.390 318.000 ;
        RECT 1946.330 317.940 1946.650 318.000 ;
      LAYER via ;
        RECT 1587.100 318.960 1587.360 319.220 ;
        RECT 1608.260 318.960 1608.520 319.220 ;
        RECT 1702.100 318.620 1702.360 318.880 ;
        RECT 1704.400 318.620 1704.660 318.880 ;
        RECT 1798.700 318.620 1798.960 318.880 ;
        RECT 1801.920 318.620 1802.180 318.880 ;
        RECT 2090.340 318.620 2090.600 318.880 ;
        RECT 2124.840 318.620 2125.100 318.880 ;
        RECT 1932.100 317.940 1932.360 318.200 ;
        RECT 1946.360 317.940 1946.620 318.200 ;
      LAYER met2 ;
        RECT 1173.090 2498.730 1173.370 2500.000 ;
        RECT 1174.470 2498.730 1174.750 2498.845 ;
        RECT 1173.090 2498.590 1174.750 2498.730 ;
        RECT 1173.090 2496.000 1173.370 2498.590 ;
        RECT 1174.470 2498.475 1174.750 2498.590 ;
        RECT 2028.230 320.435 2028.510 320.805 ;
        RECT 1283.490 319.075 1283.770 319.445 ;
        RECT 1587.090 319.075 1587.370 319.445 ;
        RECT 1283.560 318.085 1283.700 319.075 ;
        RECT 1587.100 318.930 1587.360 319.075 ;
        RECT 1608.260 318.930 1608.520 319.250 ;
        RECT 1946.350 319.075 1946.630 319.445 ;
        RECT 1608.320 318.765 1608.460 318.930 ;
        RECT 1702.100 318.765 1702.360 318.910 ;
        RECT 1704.400 318.765 1704.660 318.910 ;
        RECT 1798.700 318.765 1798.960 318.910 ;
        RECT 1801.920 318.765 1802.180 318.910 ;
        RECT 1482.670 318.650 1482.950 318.765 ;
        RECT 1483.590 318.650 1483.870 318.765 ;
        RECT 1482.670 318.510 1483.870 318.650 ;
        RECT 1482.670 318.395 1482.950 318.510 ;
        RECT 1483.590 318.395 1483.870 318.510 ;
        RECT 1608.250 318.395 1608.530 318.765 ;
        RECT 1702.090 318.395 1702.370 318.765 ;
        RECT 1704.390 318.395 1704.670 318.765 ;
        RECT 1798.690 318.395 1798.970 318.765 ;
        RECT 1801.910 318.395 1802.190 318.765 ;
        RECT 1895.290 318.395 1895.570 318.765 ;
        RECT 1283.490 317.715 1283.770 318.085 ;
        RECT 1895.360 316.725 1895.500 318.395 ;
        RECT 1946.420 318.230 1946.560 319.075 ;
        RECT 2028.300 318.765 2028.440 320.435 ;
        RECT 2052.610 319.755 2052.890 320.125 ;
        RECT 2028.230 318.395 2028.510 318.765 ;
        RECT 1932.100 318.085 1932.360 318.230 ;
        RECT 1932.090 317.715 1932.370 318.085 ;
        RECT 1946.360 317.910 1946.620 318.230 ;
        RECT 2052.680 318.085 2052.820 319.755 ;
        RECT 2124.830 319.075 2125.110 319.445 ;
        RECT 2124.900 318.910 2125.040 319.075 ;
        RECT 2090.340 318.765 2090.600 318.910 ;
        RECT 2090.330 318.395 2090.610 318.765 ;
        RECT 2124.840 318.590 2125.100 318.910 ;
        RECT 2052.610 317.715 2052.890 318.085 ;
        RECT 1895.290 316.355 1895.570 316.725 ;
      LAYER via2 ;
        RECT 1174.470 2498.520 1174.750 2498.800 ;
        RECT 2028.230 320.480 2028.510 320.760 ;
        RECT 1283.490 319.120 1283.770 319.400 ;
        RECT 1587.090 319.120 1587.370 319.400 ;
        RECT 1946.350 319.120 1946.630 319.400 ;
        RECT 1482.670 318.440 1482.950 318.720 ;
        RECT 1483.590 318.440 1483.870 318.720 ;
        RECT 1608.250 318.440 1608.530 318.720 ;
        RECT 1702.090 318.440 1702.370 318.720 ;
        RECT 1704.390 318.440 1704.670 318.720 ;
        RECT 1798.690 318.440 1798.970 318.720 ;
        RECT 1801.910 318.440 1802.190 318.720 ;
        RECT 1895.290 318.440 1895.570 318.720 ;
        RECT 1283.490 317.760 1283.770 318.040 ;
        RECT 2052.610 319.800 2052.890 320.080 ;
        RECT 2028.230 318.440 2028.510 318.720 ;
        RECT 1932.090 317.760 1932.370 318.040 ;
        RECT 2124.830 319.120 2125.110 319.400 ;
        RECT 2090.330 318.440 2090.610 318.720 ;
        RECT 2052.610 317.760 2052.890 318.040 ;
        RECT 1895.290 316.400 1895.570 316.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 322.060 2924.800 323.260 ;
=======
        RECT 1174.445 2498.810 1174.775 2498.825 ;
        RECT 1178.790 2498.810 1179.170 2498.820 ;
        RECT 1174.445 2498.510 1179.170 2498.810 ;
        RECT 1174.445 2498.495 1174.775 2498.510 ;
        RECT 1178.790 2498.500 1179.170 2498.510 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2916.710 322.510 2924.800 322.810 ;
        RECT 1980.110 320.770 1980.490 320.780 ;
        RECT 2028.205 320.770 2028.535 320.785 ;
        RECT 1538.550 320.470 1559.090 320.770 ;
        RECT 1178.790 319.410 1179.170 319.420 ;
        RECT 1248.710 319.410 1249.090 319.420 ;
        RECT 1283.465 319.410 1283.795 319.425 ;
        RECT 1538.550 319.410 1538.850 320.470 ;
        RECT 1178.790 319.110 1222.370 319.410 ;
        RECT 1178.790 319.100 1179.170 319.110 ;
        RECT 1222.070 318.050 1222.370 319.110 ;
        RECT 1248.710 319.110 1283.795 319.410 ;
        RECT 1248.710 319.100 1249.090 319.110 ;
        RECT 1283.465 319.095 1283.795 319.110 ;
        RECT 1384.910 319.240 1427.530 319.410 ;
        RECT 1428.150 319.240 1445.930 319.410 ;
        RECT 1384.910 319.110 1445.930 319.240 ;
        RECT 1248.710 318.050 1249.090 318.060 ;
        RECT 1222.070 317.750 1249.090 318.050 ;
        RECT 1248.710 317.740 1249.090 317.750 ;
        RECT 1283.465 318.050 1283.795 318.065 ;
        RECT 1384.910 318.050 1385.210 319.110 ;
        RECT 1427.230 318.940 1428.450 319.110 ;
        RECT 1445.630 318.730 1445.930 319.110 ;
        RECT 1500.830 319.110 1538.850 319.410 ;
        RECT 1558.790 319.410 1559.090 320.470 ;
        RECT 1980.110 320.470 2028.535 320.770 ;
        RECT 1980.110 320.460 1980.490 320.470 ;
        RECT 2028.205 320.455 2028.535 320.470 ;
        RECT 2052.585 320.090 2052.915 320.105 ;
        RECT 2028.910 319.790 2052.915 320.090 ;
        RECT 1587.065 319.410 1587.395 319.425 ;
        RECT 1558.790 319.110 1587.395 319.410 ;
        RECT 1482.645 318.730 1482.975 318.745 ;
        RECT 1445.630 318.430 1482.975 318.730 ;
        RECT 1482.645 318.415 1482.975 318.430 ;
        RECT 1483.565 318.730 1483.895 318.745 ;
        RECT 1500.830 318.730 1501.130 319.110 ;
        RECT 1587.065 319.095 1587.395 319.110 ;
        RECT 1946.325 319.410 1946.655 319.425 ;
        RECT 1980.110 319.410 1980.490 319.420 ;
        RECT 1946.325 319.110 1980.490 319.410 ;
        RECT 1946.325 319.095 1946.655 319.110 ;
        RECT 1980.110 319.100 1980.490 319.110 ;
        RECT 1483.565 318.430 1501.130 318.730 ;
        RECT 1608.225 318.730 1608.555 318.745 ;
        RECT 1702.065 318.730 1702.395 318.745 ;
        RECT 1608.225 318.430 1641.890 318.730 ;
        RECT 1483.565 318.415 1483.895 318.430 ;
        RECT 1608.225 318.415 1608.555 318.430 ;
        RECT 1283.465 317.750 1385.210 318.050 ;
        RECT 1641.590 318.050 1641.890 318.430 ;
        RECT 1656.310 318.430 1702.395 318.730 ;
        RECT 1656.310 318.050 1656.610 318.430 ;
        RECT 1702.065 318.415 1702.395 318.430 ;
        RECT 1704.365 318.730 1704.695 318.745 ;
        RECT 1798.665 318.730 1798.995 318.745 ;
        RECT 1704.365 318.430 1738.490 318.730 ;
        RECT 1704.365 318.415 1704.695 318.430 ;
        RECT 1641.590 317.750 1656.610 318.050 ;
        RECT 1738.190 318.050 1738.490 318.430 ;
        RECT 1752.910 318.430 1798.995 318.730 ;
        RECT 1752.910 318.050 1753.210 318.430 ;
        RECT 1798.665 318.415 1798.995 318.430 ;
        RECT 1801.885 318.730 1802.215 318.745 ;
        RECT 1895.265 318.730 1895.595 318.745 ;
        RECT 1801.885 318.430 1835.090 318.730 ;
        RECT 1801.885 318.415 1802.215 318.430 ;
        RECT 1738.190 317.750 1753.210 318.050 ;
        RECT 1834.790 318.050 1835.090 318.430 ;
        RECT 1849.510 318.430 1895.595 318.730 ;
        RECT 1849.510 318.050 1849.810 318.430 ;
        RECT 1895.265 318.415 1895.595 318.430 ;
        RECT 2028.205 318.730 2028.535 318.745 ;
        RECT 2028.910 318.730 2029.210 319.790 ;
        RECT 2052.585 319.775 2052.915 319.790 ;
        RECT 2124.805 319.410 2125.135 319.425 ;
        RECT 2124.805 319.110 2159.850 319.410 ;
        RECT 2124.805 319.095 2125.135 319.110 ;
        RECT 2090.305 318.730 2090.635 318.745 ;
        RECT 2028.205 318.430 2029.210 318.730 ;
        RECT 2076.750 318.430 2090.635 318.730 ;
        RECT 2159.550 318.730 2159.850 319.110 ;
        RECT 2208.310 319.110 2256.450 319.410 ;
        RECT 2159.550 318.430 2207.690 318.730 ;
        RECT 2028.205 318.415 2028.535 318.430 ;
        RECT 1932.065 318.050 1932.395 318.065 ;
        RECT 1834.790 317.750 1849.810 318.050 ;
        RECT 1931.390 317.750 1932.395 318.050 ;
        RECT 1283.465 317.735 1283.795 317.750 ;
        RECT 1895.265 316.690 1895.595 316.705 ;
        RECT 1931.390 316.690 1931.690 317.750 ;
        RECT 1932.065 317.735 1932.395 317.750 ;
        RECT 2052.585 318.050 2052.915 318.065 ;
        RECT 2076.750 318.050 2077.050 318.430 ;
        RECT 2090.305 318.415 2090.635 318.430 ;
        RECT 2052.585 317.750 2077.050 318.050 ;
        RECT 2207.390 318.050 2207.690 318.430 ;
        RECT 2208.310 318.050 2208.610 319.110 ;
        RECT 2256.150 318.730 2256.450 319.110 ;
        RECT 2304.910 319.110 2353.050 319.410 ;
        RECT 2256.150 318.430 2304.290 318.730 ;
        RECT 2207.390 317.750 2208.610 318.050 ;
        RECT 2303.990 318.050 2304.290 318.430 ;
        RECT 2304.910 318.050 2305.210 319.110 ;
        RECT 2352.750 318.730 2353.050 319.110 ;
        RECT 2401.510 319.110 2449.650 319.410 ;
        RECT 2352.750 318.430 2400.890 318.730 ;
        RECT 2303.990 317.750 2305.210 318.050 ;
        RECT 2400.590 318.050 2400.890 318.430 ;
        RECT 2401.510 318.050 2401.810 319.110 ;
        RECT 2449.350 318.730 2449.650 319.110 ;
        RECT 2498.110 319.110 2546.250 319.410 ;
        RECT 2449.350 318.430 2497.490 318.730 ;
        RECT 2400.590 317.750 2401.810 318.050 ;
        RECT 2497.190 318.050 2497.490 318.430 ;
        RECT 2498.110 318.050 2498.410 319.110 ;
        RECT 2545.950 318.730 2546.250 319.110 ;
        RECT 2594.710 319.110 2642.850 319.410 ;
        RECT 2545.950 318.430 2594.090 318.730 ;
        RECT 2497.190 317.750 2498.410 318.050 ;
        RECT 2593.790 318.050 2594.090 318.430 ;
        RECT 2594.710 318.050 2595.010 319.110 ;
        RECT 2642.550 318.730 2642.850 319.110 ;
        RECT 2691.310 319.110 2739.450 319.410 ;
        RECT 2642.550 318.430 2690.690 318.730 ;
        RECT 2593.790 317.750 2595.010 318.050 ;
        RECT 2690.390 318.050 2690.690 318.430 ;
        RECT 2691.310 318.050 2691.610 319.110 ;
        RECT 2739.150 318.730 2739.450 319.110 ;
        RECT 2787.910 319.110 2836.050 319.410 ;
        RECT 2739.150 318.430 2787.290 318.730 ;
        RECT 2690.390 317.750 2691.610 318.050 ;
        RECT 2786.990 318.050 2787.290 318.430 ;
        RECT 2787.910 318.050 2788.210 319.110 ;
        RECT 2835.750 318.730 2836.050 319.110 ;
        RECT 2916.710 318.730 2917.010 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
        RECT 2835.750 318.430 2883.890 318.730 ;
        RECT 2786.990 317.750 2788.210 318.050 ;
        RECT 2883.590 318.050 2883.890 318.430 ;
        RECT 2884.510 318.430 2917.010 318.730 ;
        RECT 2884.510 318.050 2884.810 318.430 ;
        RECT 2883.590 317.750 2884.810 318.050 ;
        RECT 2052.585 317.735 2052.915 317.750 ;
        RECT 1895.265 316.390 1931.690 316.690 ;
        RECT 1895.265 316.375 1895.595 316.390 ;
      LAYER via3 ;
        RECT 1178.820 2498.500 1179.140 2498.820 ;
        RECT 1178.820 319.100 1179.140 319.420 ;
        RECT 1248.740 319.100 1249.060 319.420 ;
        RECT 1248.740 317.740 1249.060 318.060 ;
        RECT 1980.140 320.460 1980.460 320.780 ;
        RECT 1980.140 319.100 1980.460 319.420 ;
      LAYER met4 ;
        RECT 1178.815 2498.495 1179.145 2498.825 ;
        RECT 1178.830 319.425 1179.130 2498.495 ;
        RECT 1980.135 320.455 1980.465 320.785 ;
        RECT 1980.150 319.425 1980.450 320.455 ;
        RECT 1178.815 319.095 1179.145 319.425 ;
        RECT 1248.735 319.095 1249.065 319.425 ;
        RECT 1980.135 319.095 1980.465 319.425 ;
        RECT 1248.750 318.065 1249.050 319.095 ;
        RECT 1248.735 317.735 1249.065 318.065 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3500.200 1176.150 3500.260 ;
        RECT 1545.670 3500.200 1545.990 3500.260 ;
        RECT 1175.830 3500.060 1545.990 3500.200 ;
        RECT 1175.830 3500.000 1176.150 3500.060 ;
        RECT 1545.670 3500.000 1545.990 3500.060 ;
      LAYER via ;
        RECT 1175.860 3500.000 1176.120 3500.260 ;
        RECT 1545.700 3500.000 1545.960 3500.260 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1175.710 3519.700 1176.270 3524.800 ;
=======
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3500.290 1176.060 3517.600 ;
        RECT 1175.860 3499.970 1176.120 3500.290 ;
        RECT 1545.700 3499.970 1545.960 3500.290 ;
        RECT 1545.760 2498.730 1545.900 3499.970 ;
        RECT 1549.830 2498.730 1550.110 2500.000 ;
        RECT 1545.760 2498.590 1550.110 2498.730 ;
        RECT 1549.830 2496.000 1550.110 2498.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 851.530 3504.960 851.850 3505.020 ;
        RECT 1566.370 3504.960 1566.690 3505.020 ;
        RECT 851.530 3504.820 1566.690 3504.960 ;
        RECT 851.530 3504.760 851.850 3504.820 ;
        RECT 1566.370 3504.760 1566.690 3504.820 ;
      LAYER via ;
        RECT 851.560 3504.760 851.820 3505.020 ;
        RECT 1566.400 3504.760 1566.660 3505.020 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 851.410 3519.700 851.970 3524.800 ;
=======
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3505.050 851.760 3517.600 ;
        RECT 851.560 3504.730 851.820 3505.050 ;
        RECT 1566.400 3504.730 1566.660 3505.050 ;
        RECT 1566.460 2498.730 1566.600 3504.730 ;
        RECT 1569.610 2498.730 1569.890 2500.000 ;
        RECT 1566.460 2498.590 1569.890 2498.730 ;
        RECT 1569.610 2496.000 1569.890 2498.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.230 3503.260 527.550 3503.320 ;
        RECT 1587.070 3503.260 1587.390 3503.320 ;
        RECT 527.230 3503.120 1587.390 3503.260 ;
        RECT 527.230 3503.060 527.550 3503.120 ;
        RECT 1587.070 3503.060 1587.390 3503.120 ;
      LAYER via ;
        RECT 527.260 3503.060 527.520 3503.320 ;
        RECT 1587.100 3503.060 1587.360 3503.320 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 527.110 3519.700 527.670 3524.800 ;
=======
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.350 527.460 3517.600 ;
        RECT 527.260 3503.030 527.520 3503.350 ;
        RECT 1587.100 3503.030 1587.360 3503.350 ;
        RECT 1587.160 2499.410 1587.300 3503.030 ;
        RECT 1589.390 2499.410 1589.670 2500.000 ;
        RECT 1587.160 2499.270 1589.670 2499.410 ;
        RECT 1589.390 2496.000 1589.670 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.560 202.790 3501.620 ;
        RECT 1607.770 3501.560 1608.090 3501.620 ;
        RECT 202.470 3501.420 1608.090 3501.560 ;
        RECT 202.470 3501.360 202.790 3501.420 ;
        RECT 1607.770 3501.360 1608.090 3501.420 ;
      LAYER via ;
        RECT 202.500 3501.360 202.760 3501.620 ;
        RECT 1607.800 3501.360 1608.060 3501.620 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 202.350 3519.700 202.910 3524.800 ;
=======
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.650 202.700 3517.600 ;
        RECT 202.500 3501.330 202.760 3501.650 ;
        RECT 1607.800 3501.330 1608.060 3501.650 ;
        RECT 1607.860 2499.410 1608.000 3501.330 ;
        RECT 1609.170 2499.410 1609.450 2500.000 ;
        RECT 1607.860 2499.270 1609.450 2499.410 ;
        RECT 1609.170 2496.000 1609.450 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 1628.470 3408.740 1628.790 3408.800 ;
        RECT 17.550 3408.600 1628.790 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 1628.470 3408.540 1628.790 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 1628.500 3408.540 1628.760 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 1628.500 3408.510 1628.760 3408.830 ;
        RECT 1628.560 2499.410 1628.700 3408.510 ;
        RECT 1628.950 2499.410 1629.230 2500.000 ;
        RECT 1628.560 2499.270 1629.230 2499.410 ;
        RECT 1628.950 2496.000 1629.230 2499.270 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3410.620 0.300 3411.820 ;
=======
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3119.060 17.410 3119.120 ;
        RECT 1642.730 3119.060 1643.050 3119.120 ;
        RECT 17.090 3118.920 1643.050 3119.060 ;
        RECT 17.090 3118.860 17.410 3118.920 ;
        RECT 1642.730 3118.860 1643.050 3118.920 ;
      LAYER via ;
        RECT 17.120 3118.860 17.380 3119.120 ;
        RECT 1642.760 3118.860 1643.020 3119.120 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 3119.150 17.320 3124.075 ;
        RECT 17.120 3118.830 17.380 3119.150 ;
        RECT 1642.760 3118.830 1643.020 3119.150 ;
        RECT 1642.820 2500.090 1642.960 3118.830 ;
        RECT 1642.820 2499.950 1645.720 2500.090 ;
        RECT 1645.580 2498.730 1645.720 2499.950 ;
        RECT 1648.730 2498.730 1649.010 2500.000 ;
        RECT 1645.580 2498.590 1649.010 2498.730 ;
        RECT 1648.730 2496.000 1649.010 2498.590 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3123.660 0.300 3124.860 ;
=======
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2836.180 17.410 2836.240 ;
        RECT 1662.970 2836.180 1663.290 2836.240 ;
        RECT 17.090 2836.040 1663.290 2836.180 ;
        RECT 17.090 2835.980 17.410 2836.040 ;
        RECT 1662.970 2835.980 1663.290 2836.040 ;
      LAYER via ;
        RECT 17.120 2835.980 17.380 2836.240 ;
        RECT 1663.000 2835.980 1663.260 2836.240 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2836.270 17.320 2836.435 ;
        RECT 17.120 2835.950 17.380 2836.270 ;
        RECT 1663.000 2835.950 1663.260 2836.270 ;
        RECT 1663.060 2501.450 1663.200 2835.950 ;
        RECT 1663.060 2501.310 1665.960 2501.450 ;
        RECT 1665.820 2498.730 1665.960 2501.310 ;
        RECT 1668.970 2498.730 1669.250 2500.000 ;
        RECT 1665.820 2498.590 1669.250 2498.730 ;
        RECT 1668.970 2496.000 1669.250 2498.590 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2836.020 0.300 2837.220 ;
=======
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2546.500 16.030 2546.560 ;
        RECT 1683.670 2546.500 1683.990 2546.560 ;
        RECT 15.710 2546.360 1683.990 2546.500 ;
        RECT 15.710 2546.300 16.030 2546.360 ;
        RECT 1683.670 2546.300 1683.990 2546.360 ;
      LAYER via ;
        RECT 15.740 2546.300 16.000 2546.560 ;
        RECT 1683.700 2546.300 1683.960 2546.560 ;
      LAYER met2 ;
        RECT 15.730 2549.475 16.010 2549.845 ;
        RECT 15.800 2546.590 15.940 2549.475 ;
        RECT 15.740 2546.270 16.000 2546.590 ;
        RECT 1683.700 2546.270 1683.960 2546.590 ;
        RECT 1683.760 2500.090 1683.900 2546.270 ;
        RECT 1683.760 2499.950 1686.200 2500.090 ;
        RECT 1686.060 2499.410 1686.200 2499.950 ;
        RECT 1688.750 2499.410 1689.030 2500.000 ;
        RECT 1686.060 2499.270 1689.030 2499.410 ;
        RECT 1688.750 2496.000 1689.030 2499.270 ;
      LAYER via2 ;
        RECT 15.730 2549.520 16.010 2549.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2549.060 0.300 2550.260 ;
=======
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 15.705 2549.810 16.035 2549.825 ;
        RECT -4.800 2549.510 16.035 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 15.705 2549.495 16.035 2549.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.530 2514.115 1708.810 2514.485 ;
        RECT 1708.600 2500.000 1708.740 2514.115 ;
        RECT 1708.530 2496.000 1708.810 2500.000 ;
      LAYER via2 ;
        RECT 1708.530 2514.160 1708.810 2514.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2261.420 0.300 2262.620 ;
=======
        RECT 1272.630 2514.450 1273.010 2514.460 ;
        RECT 1708.505 2514.450 1708.835 2514.465 ;
        RECT 1272.630 2514.150 1708.835 2514.450 ;
        RECT 1272.630 2514.140 1273.010 2514.150 ;
        RECT 1708.505 2514.135 1708.835 2514.150 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 19.590 2262.170 19.970 2262.180 ;
        RECT -4.800 2261.870 19.970 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 19.590 2261.860 19.970 2261.870 ;
      LAYER via3 ;
        RECT 1272.660 2514.140 1272.980 2514.460 ;
        RECT 19.620 2261.860 19.940 2262.180 ;
      LAYER met4 ;
        RECT 1272.655 2514.135 1272.985 2514.465 ;
        RECT 1272.670 2273.490 1272.970 2514.135 ;
        RECT 1272.230 2272.310 1273.410 2273.490 ;
        RECT 19.190 2265.510 20.370 2266.690 ;
        RECT 19.630 2262.185 19.930 2265.510 ;
        RECT 19.615 2261.855 19.945 2262.185 ;
      LAYER met5 ;
        RECT 82.460 2272.100 130.980 2273.700 ;
        RECT 82.460 2266.900 84.060 2272.100 ;
        RECT 18.980 2265.300 84.060 2266.900 ;
        RECT 129.380 2266.900 130.980 2272.100 ;
        RECT 179.060 2272.100 227.580 2273.700 ;
        RECT 179.060 2266.900 180.660 2272.100 ;
        RECT 129.380 2265.300 180.660 2266.900 ;
        RECT 225.980 2266.900 227.580 2272.100 ;
        RECT 275.660 2272.100 324.180 2273.700 ;
        RECT 275.660 2266.900 277.260 2272.100 ;
        RECT 225.980 2265.300 277.260 2266.900 ;
        RECT 322.580 2266.900 324.180 2272.100 ;
        RECT 372.260 2272.100 420.780 2273.700 ;
        RECT 372.260 2266.900 373.860 2272.100 ;
        RECT 322.580 2265.300 373.860 2266.900 ;
        RECT 419.180 2266.900 420.780 2272.100 ;
        RECT 468.860 2272.100 517.380 2273.700 ;
        RECT 468.860 2266.900 470.460 2272.100 ;
        RECT 419.180 2265.300 470.460 2266.900 ;
        RECT 515.780 2266.900 517.380 2272.100 ;
        RECT 565.460 2272.100 613.980 2273.700 ;
        RECT 565.460 2266.900 567.060 2272.100 ;
        RECT 515.780 2265.300 567.060 2266.900 ;
        RECT 612.380 2266.900 613.980 2272.100 ;
        RECT 662.060 2272.100 710.580 2273.700 ;
        RECT 662.060 2266.900 663.660 2272.100 ;
        RECT 612.380 2265.300 663.660 2266.900 ;
        RECT 708.980 2266.900 710.580 2272.100 ;
        RECT 758.660 2272.100 807.180 2273.700 ;
        RECT 758.660 2266.900 760.260 2272.100 ;
        RECT 708.980 2265.300 760.260 2266.900 ;
        RECT 805.580 2266.900 807.180 2272.100 ;
        RECT 855.260 2272.100 903.780 2273.700 ;
        RECT 855.260 2266.900 856.860 2272.100 ;
        RECT 805.580 2265.300 856.860 2266.900 ;
        RECT 902.180 2266.900 903.780 2272.100 ;
        RECT 951.860 2272.100 1000.380 2273.700 ;
        RECT 951.860 2266.900 953.460 2272.100 ;
        RECT 902.180 2265.300 953.460 2266.900 ;
        RECT 998.780 2266.900 1000.380 2272.100 ;
        RECT 1048.460 2272.100 1096.980 2273.700 ;
        RECT 1048.460 2266.900 1050.060 2272.100 ;
        RECT 998.780 2265.300 1050.060 2266.900 ;
        RECT 1095.380 2266.900 1096.980 2272.100 ;
        RECT 1145.060 2272.100 1193.580 2273.700 ;
        RECT 1145.060 2266.900 1146.660 2272.100 ;
        RECT 1095.380 2265.300 1146.660 2266.900 ;
        RECT 1191.980 2266.900 1193.580 2272.100 ;
        RECT 1241.660 2272.100 1273.620 2273.700 ;
        RECT 1241.660 2266.900 1243.260 2272.100 ;
        RECT 1191.980 2265.300 1243.260 2266.900 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1726.985 2495.005 1727.155 2496.875 ;
      LAYER mcon ;
        RECT 1726.985 2496.705 1727.155 2496.875 ;
      LAYER met1 ;
        RECT 1726.910 2496.860 1727.230 2496.920 ;
        RECT 1726.715 2496.720 1727.230 2496.860 ;
        RECT 1726.910 2496.660 1727.230 2496.720 ;
        RECT 14.790 2495.160 15.110 2495.220 ;
        RECT 1726.925 2495.160 1727.215 2495.205 ;
        RECT 14.790 2495.020 1727.215 2495.160 ;
        RECT 14.790 2494.960 15.110 2495.020 ;
        RECT 1726.925 2494.975 1727.215 2495.020 ;
      LAYER via ;
        RECT 1726.940 2496.660 1727.200 2496.920 ;
        RECT 14.820 2494.960 15.080 2495.220 ;
      LAYER met2 ;
        RECT 1726.940 2496.690 1727.200 2496.950 ;
        RECT 1728.310 2496.690 1728.590 2500.000 ;
        RECT 1726.940 2496.630 1728.590 2496.690 ;
        RECT 1727.000 2496.550 1728.590 2496.630 ;
        RECT 1728.310 2496.000 1728.590 2496.550 ;
        RECT 14.820 2494.930 15.080 2495.250 ;
        RECT 14.880 1975.245 15.020 2494.930 ;
        RECT 14.810 1974.875 15.090 1975.245 ;
      LAYER via2 ;
        RECT 14.810 1974.920 15.090 1975.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1974.460 0.300 1975.660 ;
=======
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 14.785 1975.210 15.115 1975.225 ;
        RECT -4.800 1974.910 15.115 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 14.785 1974.895 15.115 1974.910 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1269.210 554.440 1269.530 554.500 ;
        RECT 1273.350 554.440 1273.670 554.500 ;
        RECT 1269.210 554.300 1273.670 554.440 ;
        RECT 1269.210 554.240 1269.530 554.300 ;
        RECT 1273.350 554.240 1273.670 554.300 ;
        RECT 1365.810 553.760 1366.130 553.820 ;
        RECT 1393.410 553.760 1393.730 553.820 ;
        RECT 1365.810 553.620 1393.730 553.760 ;
        RECT 1365.810 553.560 1366.130 553.620 ;
        RECT 1393.410 553.560 1393.730 553.620 ;
        RECT 1702.070 553.420 1702.390 553.480 ;
        RECT 1704.370 553.420 1704.690 553.480 ;
        RECT 1702.070 553.280 1704.690 553.420 ;
        RECT 1702.070 553.220 1702.390 553.280 ;
        RECT 1704.370 553.220 1704.690 553.280 ;
        RECT 1798.670 553.420 1798.990 553.480 ;
        RECT 1801.890 553.420 1802.210 553.480 ;
        RECT 1798.670 553.280 1802.210 553.420 ;
        RECT 1798.670 553.220 1798.990 553.280 ;
        RECT 1801.890 553.220 1802.210 553.280 ;
        RECT 2090.310 553.420 2090.630 553.480 ;
        RECT 2124.810 553.420 2125.130 553.480 ;
        RECT 2090.310 553.280 2125.130 553.420 ;
        RECT 2090.310 553.220 2090.630 553.280 ;
        RECT 2124.810 553.220 2125.130 553.280 ;
        RECT 1606.390 553.080 1606.710 553.140 ;
        RECT 1607.770 553.080 1608.090 553.140 ;
        RECT 1606.390 552.940 1608.090 553.080 ;
        RECT 1606.390 552.880 1606.710 552.940 ;
        RECT 1607.770 552.880 1608.090 552.940 ;
        RECT 1932.070 552.740 1932.390 552.800 ;
        RECT 1946.330 552.740 1946.650 552.800 ;
        RECT 1932.070 552.600 1946.650 552.740 ;
        RECT 1932.070 552.540 1932.390 552.600 ;
        RECT 1946.330 552.540 1946.650 552.600 ;
      LAYER via ;
        RECT 1269.240 554.240 1269.500 554.500 ;
        RECT 1273.380 554.240 1273.640 554.500 ;
        RECT 1365.840 553.560 1366.100 553.820 ;
        RECT 1393.440 553.560 1393.700 553.820 ;
        RECT 1702.100 553.220 1702.360 553.480 ;
        RECT 1704.400 553.220 1704.660 553.480 ;
        RECT 1798.700 553.220 1798.960 553.480 ;
        RECT 1801.920 553.220 1802.180 553.480 ;
        RECT 2090.340 553.220 2090.600 553.480 ;
        RECT 2124.840 553.220 2125.100 553.480 ;
        RECT 1606.420 552.880 1606.680 553.140 ;
        RECT 1607.800 552.880 1608.060 553.140 ;
        RECT 1932.100 552.540 1932.360 552.800 ;
        RECT 1946.360 552.540 1946.620 552.800 ;
      LAYER met2 ;
        RECT 1191.490 2498.050 1191.770 2498.165 ;
        RECT 1192.870 2498.050 1193.150 2500.000 ;
        RECT 1191.490 2497.910 1193.150 2498.050 ;
        RECT 1191.490 2497.795 1191.770 2497.910 ;
        RECT 1192.870 2496.000 1193.150 2497.910 ;
        RECT 2028.230 555.035 2028.510 555.405 ;
        RECT 1269.230 554.355 1269.510 554.725 ;
        RECT 1273.370 554.355 1273.650 554.725 ;
        RECT 1269.240 554.210 1269.500 554.355 ;
        RECT 1273.380 554.210 1273.640 554.355 ;
        RECT 1365.830 553.675 1366.110 554.045 ;
        RECT 1365.840 553.530 1366.100 553.675 ;
        RECT 1393.440 553.530 1393.700 553.850 ;
        RECT 1946.350 553.675 1946.630 554.045 ;
        RECT 1393.500 553.365 1393.640 553.530 ;
        RECT 1702.100 553.365 1702.360 553.510 ;
        RECT 1704.400 553.365 1704.660 553.510 ;
        RECT 1798.700 553.365 1798.960 553.510 ;
        RECT 1801.920 553.365 1802.180 553.510 ;
        RECT 1393.430 552.995 1393.710 553.365 ;
        RECT 1606.410 552.995 1606.690 553.365 ;
        RECT 1607.790 552.995 1608.070 553.365 ;
        RECT 1702.090 552.995 1702.370 553.365 ;
        RECT 1704.390 552.995 1704.670 553.365 ;
        RECT 1798.690 552.995 1798.970 553.365 ;
        RECT 1801.910 552.995 1802.190 553.365 ;
        RECT 1895.290 552.995 1895.570 553.365 ;
        RECT 1606.420 552.850 1606.680 552.995 ;
        RECT 1607.800 552.850 1608.060 552.995 ;
        RECT 1895.360 551.325 1895.500 552.995 ;
        RECT 1946.420 552.830 1946.560 553.675 ;
        RECT 2028.300 553.365 2028.440 555.035 ;
        RECT 2052.610 554.355 2052.890 554.725 ;
        RECT 2028.230 552.995 2028.510 553.365 ;
        RECT 1932.100 552.685 1932.360 552.830 ;
        RECT 1932.090 552.315 1932.370 552.685 ;
        RECT 1946.360 552.510 1946.620 552.830 ;
        RECT 2052.680 552.685 2052.820 554.355 ;
        RECT 2124.830 553.675 2125.110 554.045 ;
        RECT 2124.900 553.510 2125.040 553.675 ;
        RECT 2090.340 553.365 2090.600 553.510 ;
        RECT 2090.330 552.995 2090.610 553.365 ;
        RECT 2124.840 553.190 2125.100 553.510 ;
        RECT 2052.610 552.315 2052.890 552.685 ;
        RECT 1895.290 550.955 1895.570 551.325 ;
      LAYER via2 ;
        RECT 1191.490 2497.840 1191.770 2498.120 ;
        RECT 2028.230 555.080 2028.510 555.360 ;
        RECT 1269.230 554.400 1269.510 554.680 ;
        RECT 1273.370 554.400 1273.650 554.680 ;
        RECT 1365.830 553.720 1366.110 554.000 ;
        RECT 1946.350 553.720 1946.630 554.000 ;
        RECT 1393.430 553.040 1393.710 553.320 ;
        RECT 1606.410 553.040 1606.690 553.320 ;
        RECT 1607.790 553.040 1608.070 553.320 ;
        RECT 1702.090 553.040 1702.370 553.320 ;
        RECT 1704.390 553.040 1704.670 553.320 ;
        RECT 1798.690 553.040 1798.970 553.320 ;
        RECT 1801.910 553.040 1802.190 553.320 ;
        RECT 1895.290 553.040 1895.570 553.320 ;
        RECT 2052.610 554.400 2052.890 554.680 ;
        RECT 2028.230 553.040 2028.510 553.320 ;
        RECT 1932.090 552.360 1932.370 552.640 ;
        RECT 2124.830 553.720 2125.110 554.000 ;
        RECT 2090.330 553.040 2090.610 553.320 ;
        RECT 2052.610 552.360 2052.890 552.640 ;
        RECT 1895.290 551.000 1895.570 551.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 556.660 2924.800 557.860 ;
=======
        RECT 1190.750 2498.130 1191.130 2498.140 ;
        RECT 1191.465 2498.130 1191.795 2498.145 ;
        RECT 1190.750 2497.830 1191.795 2498.130 ;
        RECT 1190.750 2497.820 1191.130 2497.830 ;
        RECT 1191.465 2497.815 1191.795 2497.830 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2916.710 557.110 2924.800 557.410 ;
        RECT 1980.110 555.370 1980.490 555.380 ;
        RECT 2028.205 555.370 2028.535 555.385 ;
        RECT 1980.110 555.070 2028.535 555.370 ;
        RECT 1980.110 555.060 1980.490 555.070 ;
        RECT 2028.205 555.055 2028.535 555.070 ;
        RECT 1190.750 554.690 1191.130 554.700 ;
        RECT 1269.205 554.690 1269.535 554.705 ;
        RECT 1190.750 554.390 1269.535 554.690 ;
        RECT 1190.750 554.380 1191.130 554.390 ;
        RECT 1269.205 554.375 1269.535 554.390 ;
        RECT 1273.345 554.690 1273.675 554.705 ;
        RECT 2052.585 554.690 2052.915 554.705 ;
        RECT 1273.345 554.390 1321.730 554.690 ;
        RECT 1273.345 554.375 1273.675 554.390 ;
        RECT 1321.430 554.010 1321.730 554.390 ;
        RECT 2028.910 554.390 2052.915 554.690 ;
        RECT 1365.805 554.010 1366.135 554.025 ;
        RECT 1946.325 554.010 1946.655 554.025 ;
        RECT 1980.110 554.010 1980.490 554.020 ;
        RECT 1321.430 553.710 1366.135 554.010 ;
        RECT 1365.805 553.695 1366.135 553.710 ;
        RECT 1441.030 553.710 1511.250 554.010 ;
        RECT 1393.405 553.330 1393.735 553.345 ;
        RECT 1441.030 553.330 1441.330 553.710 ;
        RECT 1393.405 553.030 1394.410 553.330 ;
        RECT 1393.405 553.015 1393.735 553.030 ;
        RECT 1394.110 552.650 1394.410 553.030 ;
        RECT 1395.030 553.030 1441.330 553.330 ;
        RECT 1395.030 552.650 1395.330 553.030 ;
        RECT 1394.110 552.350 1395.330 552.650 ;
        RECT 1510.950 552.650 1511.250 553.710 ;
        RECT 1946.325 553.710 1980.490 554.010 ;
        RECT 1946.325 553.695 1946.655 553.710 ;
        RECT 1980.110 553.700 1980.490 553.710 ;
        RECT 1606.385 553.330 1606.715 553.345 ;
        RECT 1559.710 553.030 1606.715 553.330 ;
        RECT 1559.710 552.650 1560.010 553.030 ;
        RECT 1606.385 553.015 1606.715 553.030 ;
        RECT 1607.765 553.330 1608.095 553.345 ;
        RECT 1702.065 553.330 1702.395 553.345 ;
        RECT 1607.765 553.030 1641.890 553.330 ;
        RECT 1607.765 553.015 1608.095 553.030 ;
        RECT 1510.950 552.350 1560.010 552.650 ;
        RECT 1641.590 552.650 1641.890 553.030 ;
        RECT 1656.310 553.030 1702.395 553.330 ;
        RECT 1656.310 552.650 1656.610 553.030 ;
        RECT 1702.065 553.015 1702.395 553.030 ;
        RECT 1704.365 553.330 1704.695 553.345 ;
        RECT 1798.665 553.330 1798.995 553.345 ;
        RECT 1704.365 553.030 1738.490 553.330 ;
        RECT 1704.365 553.015 1704.695 553.030 ;
        RECT 1641.590 552.350 1656.610 552.650 ;
        RECT 1738.190 552.650 1738.490 553.030 ;
        RECT 1752.910 553.030 1798.995 553.330 ;
        RECT 1752.910 552.650 1753.210 553.030 ;
        RECT 1798.665 553.015 1798.995 553.030 ;
        RECT 1801.885 553.330 1802.215 553.345 ;
        RECT 1895.265 553.330 1895.595 553.345 ;
        RECT 1801.885 553.030 1835.090 553.330 ;
        RECT 1801.885 553.015 1802.215 553.030 ;
        RECT 1738.190 552.350 1753.210 552.650 ;
        RECT 1834.790 552.650 1835.090 553.030 ;
        RECT 1849.510 553.030 1895.595 553.330 ;
        RECT 1849.510 552.650 1849.810 553.030 ;
        RECT 1895.265 553.015 1895.595 553.030 ;
        RECT 2028.205 553.330 2028.535 553.345 ;
        RECT 2028.910 553.330 2029.210 554.390 ;
        RECT 2052.585 554.375 2052.915 554.390 ;
        RECT 2124.805 554.010 2125.135 554.025 ;
        RECT 2124.805 553.710 2159.850 554.010 ;
        RECT 2124.805 553.695 2125.135 553.710 ;
        RECT 2090.305 553.330 2090.635 553.345 ;
        RECT 2028.205 553.030 2029.210 553.330 ;
        RECT 2076.750 553.030 2090.635 553.330 ;
        RECT 2159.550 553.330 2159.850 553.710 ;
        RECT 2208.310 553.710 2256.450 554.010 ;
        RECT 2159.550 553.030 2207.690 553.330 ;
        RECT 2028.205 553.015 2028.535 553.030 ;
        RECT 1932.065 552.650 1932.395 552.665 ;
        RECT 1834.790 552.350 1849.810 552.650 ;
        RECT 1931.390 552.350 1932.395 552.650 ;
        RECT 1895.265 551.290 1895.595 551.305 ;
        RECT 1931.390 551.290 1931.690 552.350 ;
        RECT 1932.065 552.335 1932.395 552.350 ;
        RECT 2052.585 552.650 2052.915 552.665 ;
        RECT 2076.750 552.650 2077.050 553.030 ;
        RECT 2090.305 553.015 2090.635 553.030 ;
        RECT 2052.585 552.350 2077.050 552.650 ;
        RECT 2207.390 552.650 2207.690 553.030 ;
        RECT 2208.310 552.650 2208.610 553.710 ;
        RECT 2256.150 553.330 2256.450 553.710 ;
        RECT 2304.910 553.710 2353.050 554.010 ;
        RECT 2256.150 553.030 2304.290 553.330 ;
        RECT 2207.390 552.350 2208.610 552.650 ;
        RECT 2303.990 552.650 2304.290 553.030 ;
        RECT 2304.910 552.650 2305.210 553.710 ;
        RECT 2352.750 553.330 2353.050 553.710 ;
        RECT 2401.510 553.710 2449.650 554.010 ;
        RECT 2352.750 553.030 2400.890 553.330 ;
        RECT 2303.990 552.350 2305.210 552.650 ;
        RECT 2400.590 552.650 2400.890 553.030 ;
        RECT 2401.510 552.650 2401.810 553.710 ;
        RECT 2449.350 553.330 2449.650 553.710 ;
        RECT 2498.110 553.710 2546.250 554.010 ;
        RECT 2449.350 553.030 2497.490 553.330 ;
        RECT 2400.590 552.350 2401.810 552.650 ;
        RECT 2497.190 552.650 2497.490 553.030 ;
        RECT 2498.110 552.650 2498.410 553.710 ;
        RECT 2545.950 553.330 2546.250 553.710 ;
        RECT 2594.710 553.710 2642.850 554.010 ;
        RECT 2545.950 553.030 2594.090 553.330 ;
        RECT 2497.190 552.350 2498.410 552.650 ;
        RECT 2593.790 552.650 2594.090 553.030 ;
        RECT 2594.710 552.650 2595.010 553.710 ;
        RECT 2642.550 553.330 2642.850 553.710 ;
        RECT 2691.310 553.710 2739.450 554.010 ;
        RECT 2642.550 553.030 2690.690 553.330 ;
        RECT 2593.790 552.350 2595.010 552.650 ;
        RECT 2690.390 552.650 2690.690 553.030 ;
        RECT 2691.310 552.650 2691.610 553.710 ;
        RECT 2739.150 553.330 2739.450 553.710 ;
        RECT 2787.910 553.710 2836.050 554.010 ;
        RECT 2739.150 553.030 2787.290 553.330 ;
        RECT 2690.390 552.350 2691.610 552.650 ;
        RECT 2786.990 552.650 2787.290 553.030 ;
        RECT 2787.910 552.650 2788.210 553.710 ;
        RECT 2835.750 553.330 2836.050 553.710 ;
        RECT 2916.710 553.330 2917.010 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2835.750 553.030 2883.890 553.330 ;
        RECT 2786.990 552.350 2788.210 552.650 ;
        RECT 2883.590 552.650 2883.890 553.030 ;
        RECT 2884.510 553.030 2917.010 553.330 ;
        RECT 2884.510 552.650 2884.810 553.030 ;
        RECT 2883.590 552.350 2884.810 552.650 ;
        RECT 2052.585 552.335 2052.915 552.350 ;
        RECT 1895.265 550.990 1931.690 551.290 ;
        RECT 1895.265 550.975 1895.595 550.990 ;
      LAYER via3 ;
        RECT 1190.780 2497.820 1191.100 2498.140 ;
        RECT 1980.140 555.060 1980.460 555.380 ;
        RECT 1190.780 554.380 1191.100 554.700 ;
        RECT 1980.140 553.700 1980.460 554.020 ;
      LAYER met4 ;
        RECT 1190.775 2497.815 1191.105 2498.145 ;
        RECT 1190.790 554.705 1191.090 2497.815 ;
        RECT 1980.135 555.055 1980.465 555.385 ;
        RECT 1190.775 554.375 1191.105 554.705 ;
        RECT 1980.150 554.025 1980.450 555.055 ;
        RECT 1980.135 553.695 1980.465 554.025 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1746.305 2494.665 1746.475 2496.875 ;
      LAYER mcon ;
        RECT 1746.305 2496.705 1746.475 2496.875 ;
      LAYER met1 ;
        RECT 1746.230 2496.860 1746.550 2496.920 ;
        RECT 1746.035 2496.720 1746.550 2496.860 ;
        RECT 1746.230 2496.660 1746.550 2496.720 ;
        RECT 16.170 2494.820 16.490 2494.880 ;
        RECT 1746.245 2494.820 1746.535 2494.865 ;
        RECT 16.170 2494.680 1746.535 2494.820 ;
        RECT 16.170 2494.620 16.490 2494.680 ;
        RECT 1746.245 2494.635 1746.535 2494.680 ;
      LAYER via ;
        RECT 1746.260 2496.660 1746.520 2496.920 ;
        RECT 16.200 2494.620 16.460 2494.880 ;
      LAYER met2 ;
        RECT 1746.260 2496.690 1746.520 2496.950 ;
        RECT 1748.090 2496.690 1748.370 2500.000 ;
        RECT 1746.260 2496.630 1748.370 2496.690 ;
        RECT 1746.320 2496.550 1748.370 2496.630 ;
        RECT 1748.090 2496.000 1748.370 2496.550 ;
        RECT 16.200 2494.590 16.460 2494.910 ;
        RECT 16.260 1687.605 16.400 2494.590 ;
        RECT 16.190 1687.235 16.470 1687.605 ;
      LAYER via2 ;
        RECT 16.190 1687.280 16.470 1687.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1686.820 0.300 1688.020 ;
=======
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 16.165 1687.570 16.495 1687.585 ;
        RECT -4.800 1687.270 16.495 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 16.165 1687.255 16.495 1687.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1766.545 2493.985 1766.715 2496.875 ;
      LAYER mcon ;
        RECT 1766.545 2496.705 1766.715 2496.875 ;
      LAYER met1 ;
        RECT 1766.470 2496.860 1766.790 2496.920 ;
        RECT 1766.275 2496.720 1766.790 2496.860 ;
        RECT 1766.470 2496.660 1766.790 2496.720 ;
        RECT 20.310 2494.140 20.630 2494.200 ;
        RECT 1766.485 2494.140 1766.775 2494.185 ;
        RECT 20.310 2494.000 1766.775 2494.140 ;
        RECT 20.310 2493.940 20.630 2494.000 ;
        RECT 1766.485 2493.955 1766.775 2494.000 ;
      LAYER via ;
        RECT 1766.500 2496.660 1766.760 2496.920 ;
        RECT 20.340 2493.940 20.600 2494.200 ;
      LAYER met2 ;
        RECT 1766.500 2496.690 1766.760 2496.950 ;
        RECT 1767.870 2496.690 1768.150 2500.000 ;
        RECT 1766.500 2496.630 1768.150 2496.690 ;
        RECT 1766.560 2496.550 1768.150 2496.630 ;
        RECT 1767.870 2496.000 1768.150 2496.550 ;
        RECT 20.340 2493.910 20.600 2494.230 ;
        RECT 20.400 1472.045 20.540 2493.910 ;
        RECT 20.330 1471.675 20.610 1472.045 ;
      LAYER via2 ;
        RECT 20.330 1471.720 20.610 1472.000 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1471.260 0.300 1472.460 ;
=======
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 20.305 1472.010 20.635 1472.025 ;
        RECT -4.800 1471.710 20.635 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 20.305 1471.695 20.635 1471.710 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1787.245 2493.305 1787.415 2496.875 ;
      LAYER mcon ;
        RECT 1787.245 2496.705 1787.415 2496.875 ;
      LAYER met1 ;
        RECT 1787.170 2496.860 1787.490 2496.920 ;
        RECT 1786.975 2496.720 1787.490 2496.860 ;
        RECT 1787.170 2496.660 1787.490 2496.720 ;
        RECT 19.850 2493.460 20.170 2493.520 ;
        RECT 1787.185 2493.460 1787.475 2493.505 ;
        RECT 19.850 2493.320 1787.475 2493.460 ;
        RECT 19.850 2493.260 20.170 2493.320 ;
        RECT 1787.185 2493.275 1787.475 2493.320 ;
      LAYER via ;
        RECT 1787.200 2496.660 1787.460 2496.920 ;
        RECT 19.880 2493.260 20.140 2493.520 ;
      LAYER met2 ;
        RECT 1787.200 2496.690 1787.460 2496.950 ;
        RECT 1787.650 2496.690 1787.930 2500.000 ;
        RECT 1787.200 2496.630 1787.930 2496.690 ;
        RECT 1787.260 2496.550 1787.930 2496.630 ;
        RECT 1787.650 2496.000 1787.930 2496.550 ;
        RECT 19.880 2493.230 20.140 2493.550 ;
        RECT 19.940 1256.485 20.080 2493.230 ;
        RECT 19.870 1256.115 20.150 1256.485 ;
      LAYER via2 ;
        RECT 19.870 1256.160 20.150 1256.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1255.700 0.300 1256.900 ;
=======
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 19.845 1256.450 20.175 1256.465 ;
        RECT -4.800 1256.150 20.175 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 19.845 1256.135 20.175 1256.150 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1806.105 2492.625 1806.275 2496.875 ;
      LAYER mcon ;
        RECT 1806.105 2496.705 1806.275 2496.875 ;
      LAYER met1 ;
        RECT 1806.030 2496.860 1806.350 2496.920 ;
        RECT 1805.835 2496.720 1806.350 2496.860 ;
        RECT 1806.030 2496.660 1806.350 2496.720 ;
        RECT 19.390 2492.780 19.710 2492.840 ;
        RECT 1806.045 2492.780 1806.335 2492.825 ;
        RECT 19.390 2492.640 1806.335 2492.780 ;
        RECT 19.390 2492.580 19.710 2492.640 ;
        RECT 1806.045 2492.595 1806.335 2492.640 ;
      LAYER via ;
        RECT 1806.060 2496.660 1806.320 2496.920 ;
        RECT 19.420 2492.580 19.680 2492.840 ;
      LAYER met2 ;
        RECT 1806.060 2496.690 1806.320 2496.950 ;
        RECT 1807.430 2496.690 1807.710 2500.000 ;
        RECT 1806.060 2496.630 1807.710 2496.690 ;
        RECT 1806.120 2496.550 1807.710 2496.630 ;
        RECT 1807.430 2496.000 1807.710 2496.550 ;
        RECT 19.420 2492.550 19.680 2492.870 ;
        RECT 19.480 1040.925 19.620 2492.550 ;
        RECT 19.410 1040.555 19.690 1040.925 ;
      LAYER via2 ;
        RECT 19.410 1040.600 19.690 1040.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1040.140 0.300 1041.340 ;
=======
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 19.385 1040.890 19.715 1040.905 ;
        RECT -4.800 1040.590 19.715 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 19.385 1040.575 19.715 1040.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1825.425 2491.945 1825.595 2496.875 ;
      LAYER mcon ;
        RECT 1825.425 2496.705 1825.595 2496.875 ;
      LAYER met1 ;
        RECT 1825.350 2496.860 1825.670 2496.920 ;
        RECT 1825.155 2496.720 1825.670 2496.860 ;
        RECT 1825.350 2496.660 1825.670 2496.720 ;
        RECT 18.930 2492.100 19.250 2492.160 ;
        RECT 1825.365 2492.100 1825.655 2492.145 ;
        RECT 18.930 2491.960 1825.655 2492.100 ;
        RECT 18.930 2491.900 19.250 2491.960 ;
        RECT 1825.365 2491.915 1825.655 2491.960 ;
      LAYER via ;
        RECT 1825.380 2496.660 1825.640 2496.920 ;
        RECT 18.960 2491.900 19.220 2492.160 ;
      LAYER met2 ;
        RECT 1825.380 2496.690 1825.640 2496.950 ;
        RECT 1827.210 2496.690 1827.490 2500.000 ;
        RECT 1825.380 2496.630 1827.490 2496.690 ;
        RECT 1825.440 2496.550 1827.490 2496.630 ;
        RECT 1827.210 2496.000 1827.490 2496.550 ;
        RECT 18.960 2491.870 19.220 2492.190 ;
        RECT 19.020 825.365 19.160 2491.870 ;
        RECT 18.950 824.995 19.230 825.365 ;
      LAYER via2 ;
        RECT 18.950 825.040 19.230 825.320 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 824.580 0.300 825.780 ;
=======
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 18.925 825.330 19.255 825.345 ;
        RECT -4.800 825.030 19.255 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 18.925 825.015 19.255 825.030 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1845.665 2491.265 1845.835 2496.875 ;
      LAYER mcon ;
        RECT 1845.665 2496.705 1845.835 2496.875 ;
      LAYER met1 ;
        RECT 1845.590 2496.860 1845.910 2496.920 ;
        RECT 1845.395 2496.720 1845.910 2496.860 ;
        RECT 1845.590 2496.660 1845.910 2496.720 ;
        RECT 18.010 2491.420 18.330 2491.480 ;
        RECT 1845.605 2491.420 1845.895 2491.465 ;
        RECT 18.010 2491.280 1845.895 2491.420 ;
        RECT 18.010 2491.220 18.330 2491.280 ;
        RECT 1845.605 2491.235 1845.895 2491.280 ;
      LAYER via ;
        RECT 1845.620 2496.660 1845.880 2496.920 ;
        RECT 18.040 2491.220 18.300 2491.480 ;
      LAYER met2 ;
        RECT 1845.620 2496.690 1845.880 2496.950 ;
        RECT 1847.450 2496.690 1847.730 2500.000 ;
        RECT 1845.620 2496.630 1847.730 2496.690 ;
        RECT 1845.680 2496.550 1847.730 2496.630 ;
        RECT 1847.450 2496.000 1847.730 2496.550 ;
        RECT 18.040 2491.190 18.300 2491.510 ;
        RECT 18.100 610.485 18.240 2491.190 ;
        RECT 18.030 610.115 18.310 610.485 ;
      LAYER via2 ;
        RECT 18.030 610.160 18.310 610.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 609.700 0.300 610.900 ;
=======
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 18.005 610.450 18.335 610.465 ;
        RECT -4.800 610.150 18.335 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 18.005 610.135 18.335 610.150 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.230 2513.435 1867.510 2513.805 ;
        RECT 1867.300 2500.000 1867.440 2513.435 ;
        RECT 1867.230 2496.000 1867.510 2500.000 ;
        RECT 17.570 399.995 17.850 400.365 ;
        RECT 17.640 394.925 17.780 399.995 ;
        RECT 17.570 394.555 17.850 394.925 ;
      LAYER via2 ;
        RECT 1867.230 2513.480 1867.510 2513.760 ;
        RECT 17.570 400.040 17.850 400.320 ;
        RECT 17.570 394.600 17.850 394.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 394.140 0.300 395.340 ;
=======
        RECT 1252.390 2513.770 1252.770 2513.780 ;
        RECT 1867.205 2513.770 1867.535 2513.785 ;
        RECT 1252.390 2513.470 1867.535 2513.770 ;
        RECT 1252.390 2513.460 1252.770 2513.470 ;
        RECT 1867.205 2513.455 1867.535 2513.470 ;
        RECT 17.545 400.330 17.875 400.345 ;
        RECT 1252.390 400.330 1252.770 400.340 ;
        RECT 17.545 400.030 1252.770 400.330 ;
        RECT 17.545 400.015 17.875 400.030 ;
        RECT 1252.390 400.020 1252.770 400.030 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.545 394.890 17.875 394.905 ;
        RECT -4.800 394.590 17.875 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.545 394.575 17.875 394.590 ;
      LAYER via3 ;
        RECT 1252.420 2513.460 1252.740 2513.780 ;
        RECT 1252.420 400.020 1252.740 400.340 ;
      LAYER met4 ;
        RECT 1252.415 2513.455 1252.745 2513.785 ;
        RECT 1252.430 400.345 1252.730 2513.455 ;
        RECT 1252.415 400.015 1252.745 400.345 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.010 2512.755 1887.290 2513.125 ;
        RECT 1887.080 2500.000 1887.220 2512.755 ;
        RECT 1887.010 2496.000 1887.290 2500.000 ;
      LAYER via2 ;
        RECT 1887.010 2512.800 1887.290 2513.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 178.580 0.300 179.780 ;
=======
        RECT 1251.470 2513.090 1251.850 2513.100 ;
        RECT 1886.985 2513.090 1887.315 2513.105 ;
        RECT 1251.470 2512.790 1887.315 2513.090 ;
        RECT 1251.470 2512.780 1251.850 2512.790 ;
        RECT 1886.985 2512.775 1887.315 2512.790 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 1251.470 179.330 1251.850 179.340 ;
        RECT -4.800 179.030 1251.850 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 1251.470 179.020 1251.850 179.030 ;
      LAYER via3 ;
        RECT 1251.500 2512.780 1251.820 2513.100 ;
        RECT 1251.500 179.020 1251.820 179.340 ;
      LAYER met4 ;
        RECT 1251.495 2512.775 1251.825 2513.105 ;
        RECT 1251.510 179.345 1251.810 2512.775 ;
        RECT 1251.495 179.015 1251.825 179.345 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1702.070 788.020 1702.390 788.080 ;
        RECT 1704.370 788.020 1704.690 788.080 ;
        RECT 1702.070 787.880 1704.690 788.020 ;
        RECT 1702.070 787.820 1702.390 787.880 ;
        RECT 1704.370 787.820 1704.690 787.880 ;
        RECT 1798.670 788.020 1798.990 788.080 ;
        RECT 1801.890 788.020 1802.210 788.080 ;
        RECT 1798.670 787.880 1802.210 788.020 ;
        RECT 1798.670 787.820 1798.990 787.880 ;
        RECT 1801.890 787.820 1802.210 787.880 ;
        RECT 2090.310 788.020 2090.630 788.080 ;
        RECT 2124.810 788.020 2125.130 788.080 ;
        RECT 2090.310 787.880 2125.130 788.020 ;
        RECT 2090.310 787.820 2090.630 787.880 ;
        RECT 2124.810 787.820 2125.130 787.880 ;
        RECT 1606.390 787.680 1606.710 787.740 ;
        RECT 1607.770 787.680 1608.090 787.740 ;
        RECT 1606.390 787.540 1608.090 787.680 ;
        RECT 1606.390 787.480 1606.710 787.540 ;
        RECT 1607.770 787.480 1608.090 787.540 ;
        RECT 1932.070 787.340 1932.390 787.400 ;
        RECT 1946.330 787.340 1946.650 787.400 ;
        RECT 1932.070 787.200 1946.650 787.340 ;
        RECT 1932.070 787.140 1932.390 787.200 ;
        RECT 1946.330 787.140 1946.650 787.200 ;
      LAYER via ;
        RECT 1702.100 787.820 1702.360 788.080 ;
        RECT 1704.400 787.820 1704.660 788.080 ;
        RECT 1798.700 787.820 1798.960 788.080 ;
        RECT 1801.920 787.820 1802.180 788.080 ;
        RECT 2090.340 787.820 2090.600 788.080 ;
        RECT 2124.840 787.820 2125.100 788.080 ;
        RECT 1606.420 787.480 1606.680 787.740 ;
        RECT 1607.800 787.480 1608.060 787.740 ;
        RECT 1932.100 787.140 1932.360 787.400 ;
        RECT 1946.360 787.140 1946.620 787.400 ;
      LAYER met2 ;
        RECT 1212.650 2498.050 1212.930 2500.000 ;
        RECT 1213.570 2498.050 1213.850 2498.165 ;
        RECT 1212.650 2497.910 1213.850 2498.050 ;
        RECT 1212.650 2496.000 1212.930 2497.910 ;
        RECT 1213.570 2497.795 1213.850 2497.910 ;
        RECT 2028.230 789.635 2028.510 790.005 ;
        RECT 1386.530 788.275 1386.810 788.645 ;
        RECT 1449.090 788.275 1449.370 788.645 ;
        RECT 1946.350 788.275 1946.630 788.645 ;
        RECT 1386.600 787.285 1386.740 788.275 ;
        RECT 1449.160 787.285 1449.300 788.275 ;
        RECT 1702.100 787.965 1702.360 788.110 ;
        RECT 1704.400 787.965 1704.660 788.110 ;
        RECT 1798.700 787.965 1798.960 788.110 ;
        RECT 1801.920 787.965 1802.180 788.110 ;
        RECT 1606.410 787.595 1606.690 787.965 ;
        RECT 1607.790 787.595 1608.070 787.965 ;
        RECT 1702.090 787.595 1702.370 787.965 ;
        RECT 1704.390 787.595 1704.670 787.965 ;
        RECT 1798.690 787.595 1798.970 787.965 ;
        RECT 1801.910 787.595 1802.190 787.965 ;
        RECT 1895.290 787.595 1895.570 787.965 ;
        RECT 1606.420 787.450 1606.680 787.595 ;
        RECT 1607.800 787.450 1608.060 787.595 ;
        RECT 1386.530 786.915 1386.810 787.285 ;
        RECT 1449.090 786.915 1449.370 787.285 ;
        RECT 1895.360 785.925 1895.500 787.595 ;
        RECT 1946.420 787.430 1946.560 788.275 ;
        RECT 2028.300 787.965 2028.440 789.635 ;
        RECT 2052.610 788.955 2052.890 789.325 ;
        RECT 2028.230 787.595 2028.510 787.965 ;
        RECT 1932.100 787.285 1932.360 787.430 ;
        RECT 1932.090 786.915 1932.370 787.285 ;
        RECT 1946.360 787.110 1946.620 787.430 ;
        RECT 2052.680 787.285 2052.820 788.955 ;
        RECT 2124.830 788.275 2125.110 788.645 ;
        RECT 2124.900 788.110 2125.040 788.275 ;
        RECT 2090.340 787.965 2090.600 788.110 ;
        RECT 2090.330 787.595 2090.610 787.965 ;
        RECT 2124.840 787.790 2125.100 788.110 ;
        RECT 2052.610 786.915 2052.890 787.285 ;
        RECT 1895.290 785.555 1895.570 785.925 ;
      LAYER via2 ;
        RECT 1213.570 2497.840 1213.850 2498.120 ;
        RECT 2028.230 789.680 2028.510 789.960 ;
        RECT 1386.530 788.320 1386.810 788.600 ;
        RECT 1449.090 788.320 1449.370 788.600 ;
        RECT 1946.350 788.320 1946.630 788.600 ;
        RECT 1606.410 787.640 1606.690 787.920 ;
        RECT 1607.790 787.640 1608.070 787.920 ;
        RECT 1702.090 787.640 1702.370 787.920 ;
        RECT 1704.390 787.640 1704.670 787.920 ;
        RECT 1798.690 787.640 1798.970 787.920 ;
        RECT 1801.910 787.640 1802.190 787.920 ;
        RECT 1895.290 787.640 1895.570 787.920 ;
        RECT 1386.530 786.960 1386.810 787.240 ;
        RECT 1449.090 786.960 1449.370 787.240 ;
        RECT 2052.610 789.000 2052.890 789.280 ;
        RECT 2028.230 787.640 2028.510 787.920 ;
        RECT 1932.090 786.960 1932.370 787.240 ;
        RECT 2124.830 788.320 2125.110 788.600 ;
        RECT 2090.330 787.640 2090.610 787.920 ;
        RECT 2052.610 786.960 2052.890 787.240 ;
        RECT 1895.290 785.600 1895.570 785.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 791.260 2924.800 792.460 ;
=======
        RECT 1213.545 2498.140 1213.875 2498.145 ;
        RECT 1213.545 2498.130 1214.130 2498.140 ;
        RECT 1213.545 2497.830 1214.330 2498.130 ;
        RECT 1213.545 2497.820 1214.130 2497.830 ;
        RECT 1213.545 2497.815 1213.875 2497.820 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2916.710 791.710 2924.800 792.010 ;
        RECT 1980.110 789.970 1980.490 789.980 ;
        RECT 2028.205 789.970 2028.535 789.985 ;
        RECT 1980.110 789.670 2028.535 789.970 ;
        RECT 1980.110 789.660 1980.490 789.670 ;
        RECT 2028.205 789.655 2028.535 789.670 ;
        RECT 2052.585 789.290 2052.915 789.305 ;
        RECT 2028.910 788.990 2052.915 789.290 ;
        RECT 1386.505 788.610 1386.835 788.625 ;
        RECT 1449.065 788.610 1449.395 788.625 ;
        RECT 1946.325 788.610 1946.655 788.625 ;
        RECT 1980.110 788.610 1980.490 788.620 ;
        RECT 1386.505 788.295 1387.050 788.610 ;
        RECT 1449.065 788.310 1559.090 788.610 ;
        RECT 1449.065 788.295 1449.395 788.310 ;
        RECT 1386.750 787.930 1387.050 788.295 ;
        RECT 1386.750 787.630 1387.970 787.930 ;
        RECT 1213.750 787.250 1214.130 787.260 ;
        RECT 1386.505 787.250 1386.835 787.265 ;
        RECT 1213.750 786.950 1248.130 787.250 ;
        RECT 1213.750 786.940 1214.130 786.950 ;
        RECT 1247.830 786.570 1248.130 786.950 ;
        RECT 1270.830 786.950 1386.835 787.250 ;
        RECT 1387.670 787.250 1387.970 787.630 ;
        RECT 1449.065 787.250 1449.395 787.265 ;
        RECT 1387.670 786.950 1449.395 787.250 ;
        RECT 1558.790 787.250 1559.090 788.310 ;
        RECT 1946.325 788.310 1980.490 788.610 ;
        RECT 1946.325 788.295 1946.655 788.310 ;
        RECT 1980.110 788.300 1980.490 788.310 ;
        RECT 1606.385 787.930 1606.715 787.945 ;
        RECT 1559.710 787.630 1606.715 787.930 ;
        RECT 1559.710 787.250 1560.010 787.630 ;
        RECT 1606.385 787.615 1606.715 787.630 ;
        RECT 1607.765 787.930 1608.095 787.945 ;
        RECT 1702.065 787.930 1702.395 787.945 ;
        RECT 1607.765 787.630 1641.890 787.930 ;
        RECT 1607.765 787.615 1608.095 787.630 ;
        RECT 1558.790 786.950 1560.010 787.250 ;
        RECT 1641.590 787.250 1641.890 787.630 ;
        RECT 1656.310 787.630 1702.395 787.930 ;
        RECT 1656.310 787.250 1656.610 787.630 ;
        RECT 1702.065 787.615 1702.395 787.630 ;
        RECT 1704.365 787.930 1704.695 787.945 ;
        RECT 1798.665 787.930 1798.995 787.945 ;
        RECT 1704.365 787.630 1738.490 787.930 ;
        RECT 1704.365 787.615 1704.695 787.630 ;
        RECT 1641.590 786.950 1656.610 787.250 ;
        RECT 1738.190 787.250 1738.490 787.630 ;
        RECT 1752.910 787.630 1798.995 787.930 ;
        RECT 1752.910 787.250 1753.210 787.630 ;
        RECT 1798.665 787.615 1798.995 787.630 ;
        RECT 1801.885 787.930 1802.215 787.945 ;
        RECT 1895.265 787.930 1895.595 787.945 ;
        RECT 1801.885 787.630 1835.090 787.930 ;
        RECT 1801.885 787.615 1802.215 787.630 ;
        RECT 1738.190 786.950 1753.210 787.250 ;
        RECT 1834.790 787.250 1835.090 787.630 ;
        RECT 1849.510 787.630 1895.595 787.930 ;
        RECT 1849.510 787.250 1849.810 787.630 ;
        RECT 1895.265 787.615 1895.595 787.630 ;
        RECT 2028.205 787.930 2028.535 787.945 ;
        RECT 2028.910 787.930 2029.210 788.990 ;
        RECT 2052.585 788.975 2052.915 788.990 ;
        RECT 2124.805 788.610 2125.135 788.625 ;
        RECT 2124.805 788.310 2159.850 788.610 ;
        RECT 2124.805 788.295 2125.135 788.310 ;
        RECT 2090.305 787.930 2090.635 787.945 ;
        RECT 2028.205 787.630 2029.210 787.930 ;
        RECT 2076.750 787.630 2090.635 787.930 ;
        RECT 2159.550 787.930 2159.850 788.310 ;
        RECT 2208.310 788.310 2256.450 788.610 ;
        RECT 2159.550 787.630 2207.690 787.930 ;
        RECT 2028.205 787.615 2028.535 787.630 ;
        RECT 1932.065 787.250 1932.395 787.265 ;
        RECT 1834.790 786.950 1849.810 787.250 ;
        RECT 1931.390 786.950 1932.395 787.250 ;
        RECT 1270.830 786.570 1271.130 786.950 ;
        RECT 1386.505 786.935 1386.835 786.950 ;
        RECT 1449.065 786.935 1449.395 786.950 ;
        RECT 1247.830 786.270 1271.130 786.570 ;
        RECT 1895.265 785.890 1895.595 785.905 ;
        RECT 1931.390 785.890 1931.690 786.950 ;
        RECT 1932.065 786.935 1932.395 786.950 ;
        RECT 2052.585 787.250 2052.915 787.265 ;
        RECT 2076.750 787.250 2077.050 787.630 ;
        RECT 2090.305 787.615 2090.635 787.630 ;
        RECT 2052.585 786.950 2077.050 787.250 ;
        RECT 2207.390 787.250 2207.690 787.630 ;
        RECT 2208.310 787.250 2208.610 788.310 ;
        RECT 2256.150 787.930 2256.450 788.310 ;
        RECT 2304.910 788.310 2353.050 788.610 ;
        RECT 2256.150 787.630 2304.290 787.930 ;
        RECT 2207.390 786.950 2208.610 787.250 ;
        RECT 2303.990 787.250 2304.290 787.630 ;
        RECT 2304.910 787.250 2305.210 788.310 ;
        RECT 2352.750 787.930 2353.050 788.310 ;
        RECT 2401.510 788.310 2449.650 788.610 ;
        RECT 2352.750 787.630 2400.890 787.930 ;
        RECT 2303.990 786.950 2305.210 787.250 ;
        RECT 2400.590 787.250 2400.890 787.630 ;
        RECT 2401.510 787.250 2401.810 788.310 ;
        RECT 2449.350 787.930 2449.650 788.310 ;
        RECT 2498.110 788.310 2546.250 788.610 ;
        RECT 2449.350 787.630 2497.490 787.930 ;
        RECT 2400.590 786.950 2401.810 787.250 ;
        RECT 2497.190 787.250 2497.490 787.630 ;
        RECT 2498.110 787.250 2498.410 788.310 ;
        RECT 2545.950 787.930 2546.250 788.310 ;
        RECT 2594.710 788.310 2642.850 788.610 ;
        RECT 2545.950 787.630 2594.090 787.930 ;
        RECT 2497.190 786.950 2498.410 787.250 ;
        RECT 2593.790 787.250 2594.090 787.630 ;
        RECT 2594.710 787.250 2595.010 788.310 ;
        RECT 2642.550 787.930 2642.850 788.310 ;
        RECT 2691.310 788.310 2739.450 788.610 ;
        RECT 2642.550 787.630 2690.690 787.930 ;
        RECT 2593.790 786.950 2595.010 787.250 ;
        RECT 2690.390 787.250 2690.690 787.630 ;
        RECT 2691.310 787.250 2691.610 788.310 ;
        RECT 2739.150 787.930 2739.450 788.310 ;
        RECT 2787.910 788.310 2836.050 788.610 ;
        RECT 2739.150 787.630 2787.290 787.930 ;
        RECT 2690.390 786.950 2691.610 787.250 ;
        RECT 2786.990 787.250 2787.290 787.630 ;
        RECT 2787.910 787.250 2788.210 788.310 ;
        RECT 2835.750 787.930 2836.050 788.310 ;
        RECT 2916.710 787.930 2917.010 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2835.750 787.630 2883.890 787.930 ;
        RECT 2786.990 786.950 2788.210 787.250 ;
        RECT 2883.590 787.250 2883.890 787.630 ;
        RECT 2884.510 787.630 2917.010 787.930 ;
        RECT 2884.510 787.250 2884.810 787.630 ;
        RECT 2883.590 786.950 2884.810 787.250 ;
        RECT 2052.585 786.935 2052.915 786.950 ;
        RECT 1895.265 785.590 1931.690 785.890 ;
        RECT 1895.265 785.575 1895.595 785.590 ;
      LAYER via3 ;
        RECT 1213.780 2497.820 1214.100 2498.140 ;
        RECT 1980.140 789.660 1980.460 789.980 ;
        RECT 1213.780 786.940 1214.100 787.260 ;
        RECT 1980.140 788.300 1980.460 788.620 ;
      LAYER met4 ;
        RECT 1213.775 2497.815 1214.105 2498.145 ;
        RECT 1213.790 787.265 1214.090 2497.815 ;
        RECT 1980.135 789.655 1980.465 789.985 ;
        RECT 1980.150 788.625 1980.450 789.655 ;
        RECT 1980.135 788.295 1980.465 788.625 ;
        RECT 1213.775 786.935 1214.105 787.265 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1365.810 1022.620 1366.130 1022.680 ;
        RECT 1369.950 1022.620 1370.270 1022.680 ;
        RECT 1365.810 1022.480 1370.270 1022.620 ;
        RECT 1365.810 1022.420 1366.130 1022.480 ;
        RECT 1369.950 1022.420 1370.270 1022.480 ;
        RECT 1702.070 1022.620 1702.390 1022.680 ;
        RECT 1704.370 1022.620 1704.690 1022.680 ;
        RECT 1702.070 1022.480 1704.690 1022.620 ;
        RECT 1702.070 1022.420 1702.390 1022.480 ;
        RECT 1704.370 1022.420 1704.690 1022.480 ;
        RECT 1798.670 1022.620 1798.990 1022.680 ;
        RECT 1801.890 1022.620 1802.210 1022.680 ;
        RECT 1798.670 1022.480 1802.210 1022.620 ;
        RECT 1798.670 1022.420 1798.990 1022.480 ;
        RECT 1801.890 1022.420 1802.210 1022.480 ;
        RECT 2090.310 1022.620 2090.630 1022.680 ;
        RECT 2124.810 1022.620 2125.130 1022.680 ;
        RECT 2090.310 1022.480 2125.130 1022.620 ;
        RECT 2090.310 1022.420 2090.630 1022.480 ;
        RECT 2124.810 1022.420 2125.130 1022.480 ;
        RECT 1606.390 1022.280 1606.710 1022.340 ;
        RECT 1607.770 1022.280 1608.090 1022.340 ;
        RECT 1606.390 1022.140 1608.090 1022.280 ;
        RECT 1606.390 1022.080 1606.710 1022.140 ;
        RECT 1607.770 1022.080 1608.090 1022.140 ;
        RECT 1932.070 1021.940 1932.390 1022.000 ;
        RECT 1946.330 1021.940 1946.650 1022.000 ;
        RECT 1932.070 1021.800 1946.650 1021.940 ;
        RECT 1932.070 1021.740 1932.390 1021.800 ;
        RECT 1946.330 1021.740 1946.650 1021.800 ;
      LAYER via ;
        RECT 1365.840 1022.420 1366.100 1022.680 ;
        RECT 1369.980 1022.420 1370.240 1022.680 ;
        RECT 1702.100 1022.420 1702.360 1022.680 ;
        RECT 1704.400 1022.420 1704.660 1022.680 ;
        RECT 1798.700 1022.420 1798.960 1022.680 ;
        RECT 1801.920 1022.420 1802.180 1022.680 ;
        RECT 2090.340 1022.420 2090.600 1022.680 ;
        RECT 2124.840 1022.420 2125.100 1022.680 ;
        RECT 1606.420 1022.080 1606.680 1022.340 ;
        RECT 1607.800 1022.080 1608.060 1022.340 ;
        RECT 1932.100 1021.740 1932.360 1022.000 ;
        RECT 1946.360 1021.740 1946.620 1022.000 ;
      LAYER met2 ;
        RECT 1232.430 2498.050 1232.710 2500.000 ;
        RECT 1233.810 2498.050 1234.090 2498.165 ;
        RECT 1232.430 2497.910 1234.090 2498.050 ;
        RECT 1232.430 2496.000 1232.710 2497.910 ;
        RECT 1233.810 2497.795 1234.090 2497.910 ;
        RECT 2028.230 1024.235 2028.510 1024.605 ;
        RECT 1466.110 1023.555 1466.390 1023.925 ;
        RECT 1365.840 1022.565 1366.100 1022.710 ;
        RECT 1369.980 1022.565 1370.240 1022.710 ;
        RECT 1365.830 1022.195 1366.110 1022.565 ;
        RECT 1369.970 1022.195 1370.250 1022.565 ;
        RECT 1466.180 1021.885 1466.320 1023.555 ;
        RECT 1496.930 1022.875 1497.210 1023.245 ;
        RECT 1946.350 1022.875 1946.630 1023.245 ;
        RECT 1497.000 1021.885 1497.140 1022.875 ;
        RECT 1702.100 1022.565 1702.360 1022.710 ;
        RECT 1704.400 1022.565 1704.660 1022.710 ;
        RECT 1798.700 1022.565 1798.960 1022.710 ;
        RECT 1801.920 1022.565 1802.180 1022.710 ;
        RECT 1606.410 1022.195 1606.690 1022.565 ;
        RECT 1607.790 1022.195 1608.070 1022.565 ;
        RECT 1702.090 1022.195 1702.370 1022.565 ;
        RECT 1704.390 1022.195 1704.670 1022.565 ;
        RECT 1798.690 1022.195 1798.970 1022.565 ;
        RECT 1801.910 1022.195 1802.190 1022.565 ;
        RECT 1895.290 1022.195 1895.570 1022.565 ;
        RECT 1606.420 1022.050 1606.680 1022.195 ;
        RECT 1607.800 1022.050 1608.060 1022.195 ;
        RECT 1466.110 1021.515 1466.390 1021.885 ;
        RECT 1496.930 1021.515 1497.210 1021.885 ;
        RECT 1895.360 1020.525 1895.500 1022.195 ;
        RECT 1946.420 1022.030 1946.560 1022.875 ;
        RECT 2028.300 1022.565 2028.440 1024.235 ;
        RECT 2052.610 1023.555 2052.890 1023.925 ;
        RECT 2028.230 1022.195 2028.510 1022.565 ;
        RECT 1932.100 1021.885 1932.360 1022.030 ;
        RECT 1932.090 1021.515 1932.370 1021.885 ;
        RECT 1946.360 1021.710 1946.620 1022.030 ;
        RECT 2052.680 1021.885 2052.820 1023.555 ;
        RECT 2124.830 1022.875 2125.110 1023.245 ;
        RECT 2124.900 1022.710 2125.040 1022.875 ;
        RECT 2090.340 1022.565 2090.600 1022.710 ;
        RECT 2090.330 1022.195 2090.610 1022.565 ;
        RECT 2124.840 1022.390 2125.100 1022.710 ;
        RECT 2052.610 1021.515 2052.890 1021.885 ;
        RECT 1895.290 1020.155 1895.570 1020.525 ;
      LAYER via2 ;
        RECT 1233.810 2497.840 1234.090 2498.120 ;
        RECT 2028.230 1024.280 2028.510 1024.560 ;
        RECT 1466.110 1023.600 1466.390 1023.880 ;
        RECT 1365.830 1022.240 1366.110 1022.520 ;
        RECT 1369.970 1022.240 1370.250 1022.520 ;
        RECT 1496.930 1022.920 1497.210 1023.200 ;
        RECT 1946.350 1022.920 1946.630 1023.200 ;
        RECT 1606.410 1022.240 1606.690 1022.520 ;
        RECT 1607.790 1022.240 1608.070 1022.520 ;
        RECT 1702.090 1022.240 1702.370 1022.520 ;
        RECT 1704.390 1022.240 1704.670 1022.520 ;
        RECT 1798.690 1022.240 1798.970 1022.520 ;
        RECT 1801.910 1022.240 1802.190 1022.520 ;
        RECT 1895.290 1022.240 1895.570 1022.520 ;
        RECT 1466.110 1021.560 1466.390 1021.840 ;
        RECT 1496.930 1021.560 1497.210 1021.840 ;
        RECT 2052.610 1023.600 2052.890 1023.880 ;
        RECT 2028.230 1022.240 2028.510 1022.520 ;
        RECT 1932.090 1021.560 1932.370 1021.840 ;
        RECT 2124.830 1022.920 2125.110 1023.200 ;
        RECT 2090.330 1022.240 2090.610 1022.520 ;
        RECT 2052.610 1021.560 2052.890 1021.840 ;
        RECT 1895.290 1020.200 1895.570 1020.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1025.860 2924.800 1027.060 ;
=======
        RECT 1233.785 2498.140 1234.115 2498.145 ;
        RECT 1233.785 2498.130 1234.370 2498.140 ;
        RECT 1233.785 2497.830 1234.570 2498.130 ;
        RECT 1233.785 2497.820 1234.370 2497.830 ;
        RECT 1233.785 2497.815 1234.115 2497.820 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2916.710 1026.310 2924.800 1026.610 ;
        RECT 1980.110 1024.570 1980.490 1024.580 ;
        RECT 2028.205 1024.570 2028.535 1024.585 ;
        RECT 1256.110 1024.270 1281.250 1024.570 ;
        RECT 1233.990 1023.890 1234.370 1023.900 ;
        RECT 1256.110 1023.890 1256.410 1024.270 ;
        RECT 1233.990 1023.590 1256.410 1023.890 ;
        RECT 1280.950 1023.890 1281.250 1024.270 ;
        RECT 1980.110 1024.270 2028.535 1024.570 ;
        RECT 1980.110 1024.260 1980.490 1024.270 ;
        RECT 2028.205 1024.255 2028.535 1024.270 ;
        RECT 1441.910 1023.890 1442.290 1023.900 ;
        RECT 1466.085 1023.890 1466.415 1023.905 ;
        RECT 2052.585 1023.890 2052.915 1023.905 ;
        RECT 1280.950 1023.590 1321.730 1023.890 ;
        RECT 1233.990 1023.580 1234.370 1023.590 ;
        RECT 1321.430 1023.210 1321.730 1023.590 ;
        RECT 1441.910 1023.590 1466.415 1023.890 ;
        RECT 1441.910 1023.580 1442.290 1023.590 ;
        RECT 1466.085 1023.575 1466.415 1023.590 ;
        RECT 2028.910 1023.590 2052.915 1023.890 ;
        RECT 1496.905 1023.210 1497.235 1023.225 ;
        RECT 1946.325 1023.210 1946.655 1023.225 ;
        RECT 1980.110 1023.210 1980.490 1023.220 ;
        RECT 1321.430 1022.910 1345.650 1023.210 ;
        RECT 1345.350 1022.530 1345.650 1022.910 ;
        RECT 1496.905 1022.910 1511.250 1023.210 ;
        RECT 1496.905 1022.895 1497.235 1022.910 ;
        RECT 1365.805 1022.530 1366.135 1022.545 ;
        RECT 1345.350 1022.230 1366.135 1022.530 ;
        RECT 1365.805 1022.215 1366.135 1022.230 ;
        RECT 1369.945 1022.530 1370.275 1022.545 ;
        RECT 1441.910 1022.530 1442.290 1022.540 ;
        RECT 1369.945 1022.230 1442.290 1022.530 ;
        RECT 1369.945 1022.215 1370.275 1022.230 ;
        RECT 1441.910 1022.220 1442.290 1022.230 ;
        RECT 1466.085 1021.850 1466.415 1021.865 ;
        RECT 1496.905 1021.850 1497.235 1021.865 ;
        RECT 1466.085 1021.550 1497.235 1021.850 ;
        RECT 1510.950 1021.850 1511.250 1022.910 ;
        RECT 1946.325 1022.910 1980.490 1023.210 ;
        RECT 1946.325 1022.895 1946.655 1022.910 ;
        RECT 1980.110 1022.900 1980.490 1022.910 ;
        RECT 1606.385 1022.530 1606.715 1022.545 ;
        RECT 1559.710 1022.230 1606.715 1022.530 ;
        RECT 1559.710 1021.850 1560.010 1022.230 ;
        RECT 1606.385 1022.215 1606.715 1022.230 ;
        RECT 1607.765 1022.530 1608.095 1022.545 ;
        RECT 1702.065 1022.530 1702.395 1022.545 ;
        RECT 1607.765 1022.230 1641.890 1022.530 ;
        RECT 1607.765 1022.215 1608.095 1022.230 ;
        RECT 1510.950 1021.550 1560.010 1021.850 ;
        RECT 1641.590 1021.850 1641.890 1022.230 ;
        RECT 1656.310 1022.230 1702.395 1022.530 ;
        RECT 1656.310 1021.850 1656.610 1022.230 ;
        RECT 1702.065 1022.215 1702.395 1022.230 ;
        RECT 1704.365 1022.530 1704.695 1022.545 ;
        RECT 1798.665 1022.530 1798.995 1022.545 ;
        RECT 1704.365 1022.230 1738.490 1022.530 ;
        RECT 1704.365 1022.215 1704.695 1022.230 ;
        RECT 1641.590 1021.550 1656.610 1021.850 ;
        RECT 1738.190 1021.850 1738.490 1022.230 ;
        RECT 1752.910 1022.230 1798.995 1022.530 ;
        RECT 1752.910 1021.850 1753.210 1022.230 ;
        RECT 1798.665 1022.215 1798.995 1022.230 ;
        RECT 1801.885 1022.530 1802.215 1022.545 ;
        RECT 1895.265 1022.530 1895.595 1022.545 ;
        RECT 1801.885 1022.230 1835.090 1022.530 ;
        RECT 1801.885 1022.215 1802.215 1022.230 ;
        RECT 1738.190 1021.550 1753.210 1021.850 ;
        RECT 1834.790 1021.850 1835.090 1022.230 ;
        RECT 1849.510 1022.230 1895.595 1022.530 ;
        RECT 1849.510 1021.850 1849.810 1022.230 ;
        RECT 1895.265 1022.215 1895.595 1022.230 ;
        RECT 2028.205 1022.530 2028.535 1022.545 ;
        RECT 2028.910 1022.530 2029.210 1023.590 ;
        RECT 2052.585 1023.575 2052.915 1023.590 ;
        RECT 2124.805 1023.210 2125.135 1023.225 ;
        RECT 2124.805 1022.910 2159.850 1023.210 ;
        RECT 2124.805 1022.895 2125.135 1022.910 ;
        RECT 2090.305 1022.530 2090.635 1022.545 ;
        RECT 2028.205 1022.230 2029.210 1022.530 ;
        RECT 2076.750 1022.230 2090.635 1022.530 ;
        RECT 2159.550 1022.530 2159.850 1022.910 ;
        RECT 2208.310 1022.910 2256.450 1023.210 ;
        RECT 2159.550 1022.230 2207.690 1022.530 ;
        RECT 2028.205 1022.215 2028.535 1022.230 ;
        RECT 1932.065 1021.850 1932.395 1021.865 ;
        RECT 1834.790 1021.550 1849.810 1021.850 ;
        RECT 1931.390 1021.550 1932.395 1021.850 ;
        RECT 1466.085 1021.535 1466.415 1021.550 ;
        RECT 1496.905 1021.535 1497.235 1021.550 ;
        RECT 1895.265 1020.490 1895.595 1020.505 ;
        RECT 1931.390 1020.490 1931.690 1021.550 ;
        RECT 1932.065 1021.535 1932.395 1021.550 ;
        RECT 2052.585 1021.850 2052.915 1021.865 ;
        RECT 2076.750 1021.850 2077.050 1022.230 ;
        RECT 2090.305 1022.215 2090.635 1022.230 ;
        RECT 2052.585 1021.550 2077.050 1021.850 ;
        RECT 2207.390 1021.850 2207.690 1022.230 ;
        RECT 2208.310 1021.850 2208.610 1022.910 ;
        RECT 2256.150 1022.530 2256.450 1022.910 ;
        RECT 2304.910 1022.910 2353.050 1023.210 ;
        RECT 2256.150 1022.230 2304.290 1022.530 ;
        RECT 2207.390 1021.550 2208.610 1021.850 ;
        RECT 2303.990 1021.850 2304.290 1022.230 ;
        RECT 2304.910 1021.850 2305.210 1022.910 ;
        RECT 2352.750 1022.530 2353.050 1022.910 ;
        RECT 2401.510 1022.910 2449.650 1023.210 ;
        RECT 2352.750 1022.230 2400.890 1022.530 ;
        RECT 2303.990 1021.550 2305.210 1021.850 ;
        RECT 2400.590 1021.850 2400.890 1022.230 ;
        RECT 2401.510 1021.850 2401.810 1022.910 ;
        RECT 2449.350 1022.530 2449.650 1022.910 ;
        RECT 2498.110 1022.910 2546.250 1023.210 ;
        RECT 2449.350 1022.230 2497.490 1022.530 ;
        RECT 2400.590 1021.550 2401.810 1021.850 ;
        RECT 2497.190 1021.850 2497.490 1022.230 ;
        RECT 2498.110 1021.850 2498.410 1022.910 ;
        RECT 2545.950 1022.530 2546.250 1022.910 ;
        RECT 2594.710 1022.910 2642.850 1023.210 ;
        RECT 2545.950 1022.230 2594.090 1022.530 ;
        RECT 2497.190 1021.550 2498.410 1021.850 ;
        RECT 2593.790 1021.850 2594.090 1022.230 ;
        RECT 2594.710 1021.850 2595.010 1022.910 ;
        RECT 2642.550 1022.530 2642.850 1022.910 ;
        RECT 2691.310 1022.910 2739.450 1023.210 ;
        RECT 2642.550 1022.230 2690.690 1022.530 ;
        RECT 2593.790 1021.550 2595.010 1021.850 ;
        RECT 2690.390 1021.850 2690.690 1022.230 ;
        RECT 2691.310 1021.850 2691.610 1022.910 ;
        RECT 2739.150 1022.530 2739.450 1022.910 ;
        RECT 2787.910 1022.910 2836.050 1023.210 ;
        RECT 2739.150 1022.230 2787.290 1022.530 ;
        RECT 2690.390 1021.550 2691.610 1021.850 ;
        RECT 2786.990 1021.850 2787.290 1022.230 ;
        RECT 2787.910 1021.850 2788.210 1022.910 ;
        RECT 2835.750 1022.530 2836.050 1022.910 ;
        RECT 2916.710 1022.530 2917.010 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2835.750 1022.230 2883.890 1022.530 ;
        RECT 2786.990 1021.550 2788.210 1021.850 ;
        RECT 2883.590 1021.850 2883.890 1022.230 ;
        RECT 2884.510 1022.230 2917.010 1022.530 ;
        RECT 2884.510 1021.850 2884.810 1022.230 ;
        RECT 2883.590 1021.550 2884.810 1021.850 ;
        RECT 2052.585 1021.535 2052.915 1021.550 ;
        RECT 1895.265 1020.190 1931.690 1020.490 ;
        RECT 1895.265 1020.175 1895.595 1020.190 ;
      LAYER via3 ;
        RECT 1234.020 2497.820 1234.340 2498.140 ;
        RECT 1234.020 1023.580 1234.340 1023.900 ;
        RECT 1980.140 1024.260 1980.460 1024.580 ;
        RECT 1441.940 1023.580 1442.260 1023.900 ;
        RECT 1441.940 1022.220 1442.260 1022.540 ;
        RECT 1980.140 1022.900 1980.460 1023.220 ;
      LAYER met4 ;
        RECT 1234.015 2497.815 1234.345 2498.145 ;
        RECT 1234.030 1023.905 1234.330 2497.815 ;
        RECT 1980.135 1024.255 1980.465 1024.585 ;
        RECT 1234.015 1023.575 1234.345 1023.905 ;
        RECT 1441.935 1023.575 1442.265 1023.905 ;
        RECT 1441.950 1022.545 1442.250 1023.575 ;
        RECT 1980.150 1023.225 1980.450 1024.255 ;
        RECT 1980.135 1022.895 1980.465 1023.225 ;
        RECT 1441.935 1022.215 1442.265 1022.545 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1798.670 1257.220 1798.990 1257.280 ;
        RECT 1811.550 1257.220 1811.870 1257.280 ;
        RECT 1798.670 1257.080 1811.870 1257.220 ;
        RECT 1798.670 1257.020 1798.990 1257.080 ;
        RECT 1811.550 1257.020 1811.870 1257.080 ;
        RECT 2090.310 1257.220 2090.630 1257.280 ;
        RECT 2124.810 1257.220 2125.130 1257.280 ;
        RECT 2090.310 1257.080 2125.130 1257.220 ;
        RECT 2090.310 1257.020 2090.630 1257.080 ;
        RECT 2124.810 1257.020 2125.130 1257.080 ;
        RECT 1690.570 1256.880 1690.890 1256.940 ;
        RECT 1704.370 1256.880 1704.690 1256.940 ;
        RECT 1690.570 1256.740 1704.690 1256.880 ;
        RECT 1690.570 1256.680 1690.890 1256.740 ;
        RECT 1704.370 1256.680 1704.690 1256.740 ;
        RECT 1895.270 1256.540 1895.590 1256.600 ;
        RECT 1930.230 1256.540 1930.550 1256.600 ;
        RECT 1895.270 1256.400 1930.550 1256.540 ;
        RECT 1895.270 1256.340 1895.590 1256.400 ;
        RECT 1930.230 1256.340 1930.550 1256.400 ;
        RECT 1932.070 1256.540 1932.390 1256.600 ;
        RECT 1956.450 1256.540 1956.770 1256.600 ;
        RECT 1932.070 1256.400 1956.770 1256.540 ;
        RECT 1932.070 1256.340 1932.390 1256.400 ;
        RECT 1956.450 1256.340 1956.770 1256.400 ;
        RECT 2042.010 1256.200 2042.330 1256.260 ;
        RECT 2069.610 1256.200 2069.930 1256.260 ;
        RECT 2042.010 1256.060 2069.930 1256.200 ;
        RECT 2042.010 1256.000 2042.330 1256.060 ;
        RECT 2069.610 1256.000 2069.930 1256.060 ;
      LAYER via ;
        RECT 1798.700 1257.020 1798.960 1257.280 ;
        RECT 1811.580 1257.020 1811.840 1257.280 ;
        RECT 2090.340 1257.020 2090.600 1257.280 ;
        RECT 2124.840 1257.020 2125.100 1257.280 ;
        RECT 1690.600 1256.680 1690.860 1256.940 ;
        RECT 1704.400 1256.680 1704.660 1256.940 ;
        RECT 1895.300 1256.340 1895.560 1256.600 ;
        RECT 1930.260 1256.340 1930.520 1256.600 ;
        RECT 1932.100 1256.340 1932.360 1256.600 ;
        RECT 1956.480 1256.340 1956.740 1256.600 ;
        RECT 2042.040 1256.000 2042.300 1256.260 ;
        RECT 2069.640 1256.000 2069.900 1256.260 ;
      LAYER met2 ;
        RECT 1252.210 2498.050 1252.490 2500.000 ;
        RECT 1253.590 2498.050 1253.870 2498.165 ;
        RECT 1252.210 2497.910 1253.870 2498.050 ;
        RECT 1252.210 2496.000 1252.490 2497.910 ;
        RECT 1253.590 2497.795 1253.870 2497.910 ;
        RECT 1956.470 1257.475 1956.750 1257.845 ;
        RECT 1993.730 1257.475 1994.010 1257.845 ;
        RECT 2124.830 1257.475 2125.110 1257.845 ;
        RECT 1798.700 1257.165 1798.960 1257.310 ;
        RECT 1811.580 1257.165 1811.840 1257.310 ;
        RECT 1690.590 1256.795 1690.870 1257.165 ;
        RECT 1704.390 1256.795 1704.670 1257.165 ;
        RECT 1798.690 1256.795 1798.970 1257.165 ;
        RECT 1811.570 1256.795 1811.850 1257.165 ;
        RECT 1895.290 1256.795 1895.570 1257.165 ;
        RECT 1690.600 1256.650 1690.860 1256.795 ;
        RECT 1704.400 1256.650 1704.660 1256.795 ;
        RECT 1895.360 1256.630 1895.500 1256.795 ;
        RECT 1895.300 1256.310 1895.560 1256.630 ;
        RECT 1930.250 1256.285 1930.530 1256.655 ;
        RECT 1956.540 1256.630 1956.680 1257.475 ;
        RECT 1993.800 1257.050 1993.940 1257.475 ;
        RECT 2124.900 1257.310 2125.040 1257.475 ;
        RECT 2090.340 1257.165 2090.600 1257.310 ;
        RECT 1994.650 1257.050 1994.930 1257.165 ;
        RECT 1993.800 1256.910 1994.930 1257.050 ;
        RECT 1994.650 1256.795 1994.930 1256.910 ;
        RECT 2090.330 1256.795 2090.610 1257.165 ;
        RECT 2124.840 1256.990 2125.100 1257.310 ;
        RECT 1932.100 1256.485 1932.360 1256.630 ;
        RECT 1932.090 1256.115 1932.370 1256.485 ;
        RECT 1956.480 1256.310 1956.740 1256.630 ;
        RECT 2042.030 1256.115 2042.310 1256.485 ;
        RECT 2069.630 1256.115 2069.910 1256.485 ;
        RECT 2042.040 1255.970 2042.300 1256.115 ;
        RECT 2069.640 1255.970 2069.900 1256.115 ;
      LAYER via2 ;
        RECT 1253.590 2497.840 1253.870 2498.120 ;
        RECT 1956.470 1257.520 1956.750 1257.800 ;
        RECT 1993.730 1257.520 1994.010 1257.800 ;
        RECT 2124.830 1257.520 2125.110 1257.800 ;
        RECT 1690.590 1256.840 1690.870 1257.120 ;
        RECT 1704.390 1256.840 1704.670 1257.120 ;
        RECT 1798.690 1256.840 1798.970 1257.120 ;
        RECT 1811.570 1256.840 1811.850 1257.120 ;
        RECT 1895.290 1256.840 1895.570 1257.120 ;
        RECT 1994.650 1256.840 1994.930 1257.120 ;
        RECT 2090.330 1256.840 2090.610 1257.120 ;
        RECT 1930.250 1256.330 1930.530 1256.610 ;
        RECT 1932.090 1256.160 1932.370 1256.440 ;
        RECT 2042.030 1256.160 2042.310 1256.440 ;
        RECT 2069.630 1256.160 2069.910 1256.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1260.460 2924.800 1261.660 ;
=======
        RECT 1253.565 2498.130 1253.895 2498.145 ;
        RECT 1255.150 2498.130 1255.530 2498.140 ;
        RECT 1253.565 2497.830 1255.530 2498.130 ;
        RECT 1253.565 2497.815 1253.895 2497.830 ;
        RECT 1255.150 2497.820 1255.530 2497.830 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2916.710 1260.910 2924.800 1261.210 ;
        RECT 1442.830 1257.810 1443.210 1257.820 ;
        RECT 1956.445 1257.810 1956.775 1257.825 ;
        RECT 1993.705 1257.810 1994.035 1257.825 ;
        RECT 1442.830 1257.510 1562.770 1257.810 ;
        RECT 1442.830 1257.500 1443.210 1257.510 ;
        RECT 1562.470 1257.130 1562.770 1257.510 ;
        RECT 1956.445 1257.510 1994.035 1257.810 ;
        RECT 1956.445 1257.495 1956.775 1257.510 ;
        RECT 1993.705 1257.495 1994.035 1257.510 ;
        RECT 2124.805 1257.810 2125.135 1257.825 ;
        RECT 2124.805 1257.510 2159.850 1257.810 ;
        RECT 2124.805 1257.495 2125.135 1257.510 ;
        RECT 1690.565 1257.130 1690.895 1257.145 ;
        RECT 1369.270 1256.830 1442.250 1257.130 ;
        RECT 1562.470 1256.830 1606.930 1257.130 ;
        RECT 1255.150 1256.450 1255.530 1256.460 ;
        RECT 1369.270 1256.450 1369.570 1256.830 ;
        RECT 1441.950 1256.460 1442.250 1256.830 ;
        RECT 1255.150 1256.150 1365.890 1256.450 ;
        RECT 1255.150 1256.140 1255.530 1256.150 ;
        RECT 1365.590 1255.940 1365.890 1256.150 ;
        RECT 1366.510 1256.150 1369.570 1256.450 ;
        RECT 1366.510 1255.940 1366.810 1256.150 ;
        RECT 1441.910 1256.140 1442.290 1256.460 ;
        RECT 1606.630 1256.450 1606.930 1256.830 ;
        RECT 1656.310 1256.830 1690.895 1257.130 ;
        RECT 1656.310 1256.450 1656.610 1256.830 ;
        RECT 1690.565 1256.815 1690.895 1256.830 ;
        RECT 1704.365 1257.130 1704.695 1257.145 ;
        RECT 1798.665 1257.130 1798.995 1257.145 ;
        RECT 1704.365 1256.830 1738.490 1257.130 ;
        RECT 1704.365 1256.815 1704.695 1256.830 ;
        RECT 1606.630 1256.150 1656.610 1256.450 ;
        RECT 1738.190 1256.450 1738.490 1256.830 ;
        RECT 1752.910 1256.830 1798.995 1257.130 ;
        RECT 1752.910 1256.450 1753.210 1256.830 ;
        RECT 1798.665 1256.815 1798.995 1256.830 ;
        RECT 1811.545 1257.130 1811.875 1257.145 ;
        RECT 1895.265 1257.130 1895.595 1257.145 ;
        RECT 1811.545 1256.830 1835.090 1257.130 ;
        RECT 1811.545 1256.815 1811.875 1256.830 ;
        RECT 1738.190 1256.150 1753.210 1256.450 ;
        RECT 1834.790 1256.450 1835.090 1256.830 ;
        RECT 1849.510 1256.830 1895.595 1257.130 ;
        RECT 1849.510 1256.450 1849.810 1256.830 ;
        RECT 1895.265 1256.815 1895.595 1256.830 ;
        RECT 1994.625 1257.130 1994.955 1257.145 ;
        RECT 2090.305 1257.130 2090.635 1257.145 ;
        RECT 1994.625 1256.830 2021.850 1257.130 ;
        RECT 1994.625 1256.815 1994.955 1256.830 ;
        RECT 1834.790 1256.150 1849.810 1256.450 ;
        RECT 1930.225 1256.620 1930.555 1256.635 ;
        RECT 1930.225 1256.450 1931.690 1256.620 ;
        RECT 1932.065 1256.450 1932.395 1256.465 ;
        RECT 1930.225 1256.320 1932.395 1256.450 ;
        RECT 1930.225 1256.305 1930.555 1256.320 ;
        RECT 1931.390 1256.150 1932.395 1256.320 ;
        RECT 2021.550 1256.450 2021.850 1256.830 ;
        RECT 2076.750 1256.830 2090.635 1257.130 ;
        RECT 2159.550 1257.130 2159.850 1257.510 ;
        RECT 2208.310 1257.510 2256.450 1257.810 ;
        RECT 2159.550 1256.830 2207.690 1257.130 ;
        RECT 2042.005 1256.450 2042.335 1256.465 ;
        RECT 2021.550 1256.150 2042.335 1256.450 ;
        RECT 1932.065 1256.135 1932.395 1256.150 ;
        RECT 2042.005 1256.135 2042.335 1256.150 ;
        RECT 2069.605 1256.450 2069.935 1256.465 ;
        RECT 2076.750 1256.450 2077.050 1256.830 ;
        RECT 2090.305 1256.815 2090.635 1256.830 ;
        RECT 2069.605 1256.150 2077.050 1256.450 ;
        RECT 2207.390 1256.450 2207.690 1256.830 ;
        RECT 2208.310 1256.450 2208.610 1257.510 ;
        RECT 2256.150 1257.130 2256.450 1257.510 ;
        RECT 2304.910 1257.510 2353.050 1257.810 ;
        RECT 2256.150 1256.830 2304.290 1257.130 ;
        RECT 2207.390 1256.150 2208.610 1256.450 ;
        RECT 2303.990 1256.450 2304.290 1256.830 ;
        RECT 2304.910 1256.450 2305.210 1257.510 ;
        RECT 2352.750 1257.130 2353.050 1257.510 ;
        RECT 2401.510 1257.510 2449.650 1257.810 ;
        RECT 2352.750 1256.830 2400.890 1257.130 ;
        RECT 2303.990 1256.150 2305.210 1256.450 ;
        RECT 2400.590 1256.450 2400.890 1256.830 ;
        RECT 2401.510 1256.450 2401.810 1257.510 ;
        RECT 2449.350 1257.130 2449.650 1257.510 ;
        RECT 2498.110 1257.510 2546.250 1257.810 ;
        RECT 2449.350 1256.830 2497.490 1257.130 ;
        RECT 2400.590 1256.150 2401.810 1256.450 ;
        RECT 2497.190 1256.450 2497.490 1256.830 ;
        RECT 2498.110 1256.450 2498.410 1257.510 ;
        RECT 2545.950 1257.130 2546.250 1257.510 ;
        RECT 2594.710 1257.510 2642.850 1257.810 ;
        RECT 2545.950 1256.830 2594.090 1257.130 ;
        RECT 2497.190 1256.150 2498.410 1256.450 ;
        RECT 2593.790 1256.450 2594.090 1256.830 ;
        RECT 2594.710 1256.450 2595.010 1257.510 ;
        RECT 2642.550 1257.130 2642.850 1257.510 ;
        RECT 2691.310 1257.510 2739.450 1257.810 ;
        RECT 2642.550 1256.830 2690.690 1257.130 ;
        RECT 2593.790 1256.150 2595.010 1256.450 ;
        RECT 2690.390 1256.450 2690.690 1256.830 ;
        RECT 2691.310 1256.450 2691.610 1257.510 ;
        RECT 2739.150 1257.130 2739.450 1257.510 ;
        RECT 2787.910 1257.510 2836.050 1257.810 ;
        RECT 2739.150 1256.830 2787.290 1257.130 ;
        RECT 2690.390 1256.150 2691.610 1256.450 ;
        RECT 2786.990 1256.450 2787.290 1256.830 ;
        RECT 2787.910 1256.450 2788.210 1257.510 ;
        RECT 2835.750 1257.130 2836.050 1257.510 ;
        RECT 2916.710 1257.130 2917.010 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2835.750 1256.830 2883.890 1257.130 ;
        RECT 2786.990 1256.150 2788.210 1256.450 ;
        RECT 2883.590 1256.450 2883.890 1256.830 ;
        RECT 2884.510 1256.830 2917.010 1257.130 ;
        RECT 2884.510 1256.450 2884.810 1256.830 ;
        RECT 2883.590 1256.150 2884.810 1256.450 ;
        RECT 2069.605 1256.135 2069.935 1256.150 ;
        RECT 1365.590 1255.640 1366.810 1255.940 ;
      LAYER via3 ;
        RECT 1255.180 2497.820 1255.500 2498.140 ;
        RECT 1442.860 1257.500 1443.180 1257.820 ;
        RECT 1255.180 1256.140 1255.500 1256.460 ;
        RECT 1441.940 1256.140 1442.260 1256.460 ;
      LAYER met4 ;
        RECT 1255.175 2497.815 1255.505 2498.145 ;
        RECT 1255.190 1256.465 1255.490 2497.815 ;
        RECT 1442.855 1257.495 1443.185 1257.825 ;
        RECT 1255.175 1256.135 1255.505 1256.465 ;
        RECT 1441.935 1256.450 1442.265 1256.465 ;
        RECT 1442.870 1256.450 1443.170 1257.495 ;
        RECT 1441.935 1256.150 1443.170 1256.450 ;
        RECT 1441.935 1256.135 1442.265 1256.150 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1365.810 1491.820 1366.130 1491.880 ;
        RECT 1369.950 1491.820 1370.270 1491.880 ;
        RECT 1365.810 1491.680 1370.270 1491.820 ;
        RECT 1365.810 1491.620 1366.130 1491.680 ;
        RECT 1369.950 1491.620 1370.270 1491.680 ;
        RECT 1702.070 1491.820 1702.390 1491.880 ;
        RECT 1704.370 1491.820 1704.690 1491.880 ;
        RECT 1702.070 1491.680 1704.690 1491.820 ;
        RECT 1702.070 1491.620 1702.390 1491.680 ;
        RECT 1704.370 1491.620 1704.690 1491.680 ;
        RECT 1798.670 1491.820 1798.990 1491.880 ;
        RECT 1801.890 1491.820 1802.210 1491.880 ;
        RECT 1798.670 1491.680 1802.210 1491.820 ;
        RECT 1798.670 1491.620 1798.990 1491.680 ;
        RECT 1801.890 1491.620 1802.210 1491.680 ;
        RECT 2090.310 1491.820 2090.630 1491.880 ;
        RECT 2124.810 1491.820 2125.130 1491.880 ;
        RECT 2090.310 1491.680 2125.130 1491.820 ;
        RECT 2090.310 1491.620 2090.630 1491.680 ;
        RECT 2124.810 1491.620 2125.130 1491.680 ;
        RECT 1606.390 1491.480 1606.710 1491.540 ;
        RECT 1607.770 1491.480 1608.090 1491.540 ;
        RECT 1606.390 1491.340 1608.090 1491.480 ;
        RECT 1606.390 1491.280 1606.710 1491.340 ;
        RECT 1607.770 1491.280 1608.090 1491.340 ;
        RECT 1932.070 1491.140 1932.390 1491.200 ;
        RECT 1946.330 1491.140 1946.650 1491.200 ;
        RECT 1932.070 1491.000 1946.650 1491.140 ;
        RECT 1932.070 1490.940 1932.390 1491.000 ;
        RECT 1946.330 1490.940 1946.650 1491.000 ;
      LAYER via ;
        RECT 1365.840 1491.620 1366.100 1491.880 ;
        RECT 1369.980 1491.620 1370.240 1491.880 ;
        RECT 1702.100 1491.620 1702.360 1491.880 ;
        RECT 1704.400 1491.620 1704.660 1491.880 ;
        RECT 1798.700 1491.620 1798.960 1491.880 ;
        RECT 1801.920 1491.620 1802.180 1491.880 ;
        RECT 2090.340 1491.620 2090.600 1491.880 ;
        RECT 2124.840 1491.620 2125.100 1491.880 ;
        RECT 1606.420 1491.280 1606.680 1491.540 ;
        RECT 1607.800 1491.280 1608.060 1491.540 ;
        RECT 1932.100 1490.940 1932.360 1491.200 ;
        RECT 1946.360 1490.940 1946.620 1491.200 ;
      LAYER met2 ;
        RECT 1271.990 2498.050 1272.270 2500.000 ;
        RECT 1273.830 2498.050 1274.110 2498.165 ;
        RECT 1271.990 2497.910 1274.110 2498.050 ;
        RECT 1271.990 2496.000 1272.270 2497.910 ;
        RECT 1273.830 2497.795 1274.110 2497.910 ;
        RECT 2028.230 1493.435 2028.510 1493.805 ;
        RECT 1483.130 1492.755 1483.410 1493.125 ;
        RECT 1365.840 1491.765 1366.100 1491.910 ;
        RECT 1369.980 1491.765 1370.240 1491.910 ;
        RECT 1365.830 1491.395 1366.110 1491.765 ;
        RECT 1369.970 1491.395 1370.250 1491.765 ;
        RECT 1483.200 1491.085 1483.340 1492.755 ;
        RECT 1946.350 1492.075 1946.630 1492.445 ;
        RECT 1702.100 1491.765 1702.360 1491.910 ;
        RECT 1704.400 1491.765 1704.660 1491.910 ;
        RECT 1798.700 1491.765 1798.960 1491.910 ;
        RECT 1801.920 1491.765 1802.180 1491.910 ;
        RECT 1497.850 1491.395 1498.130 1491.765 ;
        RECT 1606.410 1491.395 1606.690 1491.765 ;
        RECT 1607.790 1491.395 1608.070 1491.765 ;
        RECT 1702.090 1491.395 1702.370 1491.765 ;
        RECT 1704.390 1491.395 1704.670 1491.765 ;
        RECT 1798.690 1491.395 1798.970 1491.765 ;
        RECT 1801.910 1491.395 1802.190 1491.765 ;
        RECT 1895.290 1491.395 1895.570 1491.765 ;
        RECT 1483.130 1490.715 1483.410 1491.085 ;
        RECT 1496.930 1490.970 1497.210 1491.085 ;
        RECT 1497.920 1490.970 1498.060 1491.395 ;
        RECT 1606.420 1491.250 1606.680 1491.395 ;
        RECT 1607.800 1491.250 1608.060 1491.395 ;
        RECT 1496.930 1490.830 1498.060 1490.970 ;
        RECT 1496.930 1490.715 1497.210 1490.830 ;
        RECT 1895.360 1489.725 1895.500 1491.395 ;
        RECT 1946.420 1491.230 1946.560 1492.075 ;
        RECT 2028.300 1491.765 2028.440 1493.435 ;
        RECT 2052.610 1492.755 2052.890 1493.125 ;
        RECT 2028.230 1491.395 2028.510 1491.765 ;
        RECT 1932.100 1491.085 1932.360 1491.230 ;
        RECT 1932.090 1490.715 1932.370 1491.085 ;
        RECT 1946.360 1490.910 1946.620 1491.230 ;
        RECT 2052.680 1491.085 2052.820 1492.755 ;
        RECT 2124.830 1492.075 2125.110 1492.445 ;
        RECT 2124.900 1491.910 2125.040 1492.075 ;
        RECT 2090.340 1491.765 2090.600 1491.910 ;
        RECT 2090.330 1491.395 2090.610 1491.765 ;
        RECT 2124.840 1491.590 2125.100 1491.910 ;
        RECT 2052.610 1490.715 2052.890 1491.085 ;
        RECT 1895.290 1489.355 1895.570 1489.725 ;
      LAYER via2 ;
        RECT 1273.830 2497.840 1274.110 2498.120 ;
        RECT 2028.230 1493.480 2028.510 1493.760 ;
        RECT 1483.130 1492.800 1483.410 1493.080 ;
        RECT 1365.830 1491.440 1366.110 1491.720 ;
        RECT 1369.970 1491.440 1370.250 1491.720 ;
        RECT 1946.350 1492.120 1946.630 1492.400 ;
        RECT 1497.850 1491.440 1498.130 1491.720 ;
        RECT 1606.410 1491.440 1606.690 1491.720 ;
        RECT 1607.790 1491.440 1608.070 1491.720 ;
        RECT 1702.090 1491.440 1702.370 1491.720 ;
        RECT 1704.390 1491.440 1704.670 1491.720 ;
        RECT 1798.690 1491.440 1798.970 1491.720 ;
        RECT 1801.910 1491.440 1802.190 1491.720 ;
        RECT 1895.290 1491.440 1895.570 1491.720 ;
        RECT 1483.130 1490.760 1483.410 1491.040 ;
        RECT 1496.930 1490.760 1497.210 1491.040 ;
        RECT 2052.610 1492.800 2052.890 1493.080 ;
        RECT 2028.230 1491.440 2028.510 1491.720 ;
        RECT 1932.090 1490.760 1932.370 1491.040 ;
        RECT 2124.830 1492.120 2125.110 1492.400 ;
        RECT 2090.330 1491.440 2090.610 1491.720 ;
        RECT 2052.610 1490.760 2052.890 1491.040 ;
        RECT 1895.290 1489.400 1895.570 1489.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1495.060 2924.800 1496.260 ;
=======
        RECT 1273.805 2498.130 1274.135 2498.145 ;
        RECT 1275.390 2498.130 1275.770 2498.140 ;
        RECT 1273.805 2497.830 1275.770 2498.130 ;
        RECT 1273.805 2497.815 1274.135 2497.830 ;
        RECT 1275.390 2497.820 1275.770 2497.830 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2916.710 1495.510 2924.800 1495.810 ;
        RECT 1980.110 1493.770 1980.490 1493.780 ;
        RECT 2028.205 1493.770 2028.535 1493.785 ;
        RECT 1980.110 1493.470 2028.535 1493.770 ;
        RECT 1980.110 1493.460 1980.490 1493.470 ;
        RECT 2028.205 1493.455 2028.535 1493.470 ;
        RECT 1435.470 1493.090 1435.850 1493.100 ;
        RECT 1483.105 1493.090 1483.435 1493.105 ;
        RECT 2052.585 1493.090 2052.915 1493.105 ;
        RECT 1435.470 1492.790 1483.435 1493.090 ;
        RECT 1435.470 1492.780 1435.850 1492.790 ;
        RECT 1483.105 1492.775 1483.435 1492.790 ;
        RECT 2028.910 1492.790 2052.915 1493.090 ;
        RECT 1275.390 1492.410 1275.770 1492.420 ;
        RECT 1946.325 1492.410 1946.655 1492.425 ;
        RECT 1980.110 1492.410 1980.490 1492.420 ;
        RECT 1275.390 1492.110 1296.890 1492.410 ;
        RECT 1275.390 1492.100 1275.770 1492.110 ;
        RECT 1296.590 1491.730 1296.890 1492.110 ;
        RECT 1544.990 1492.110 1546.210 1492.410 ;
        RECT 1365.805 1491.730 1366.135 1491.745 ;
        RECT 1296.590 1491.430 1321.730 1491.730 ;
        RECT 1321.430 1491.050 1321.730 1491.430 ;
        RECT 1345.350 1491.430 1366.135 1491.730 ;
        RECT 1345.350 1491.050 1345.650 1491.430 ;
        RECT 1365.805 1491.415 1366.135 1491.430 ;
        RECT 1369.945 1491.730 1370.275 1491.745 ;
        RECT 1435.470 1491.730 1435.850 1491.740 ;
        RECT 1369.945 1491.430 1435.850 1491.730 ;
        RECT 1369.945 1491.415 1370.275 1491.430 ;
        RECT 1435.470 1491.420 1435.850 1491.430 ;
        RECT 1497.825 1491.730 1498.155 1491.745 ;
        RECT 1544.990 1491.730 1545.290 1492.110 ;
        RECT 1497.825 1491.430 1545.290 1491.730 ;
        RECT 1545.910 1491.730 1546.210 1492.110 ;
        RECT 1946.325 1492.110 1980.490 1492.410 ;
        RECT 1946.325 1492.095 1946.655 1492.110 ;
        RECT 1980.110 1492.100 1980.490 1492.110 ;
        RECT 1606.385 1491.730 1606.715 1491.745 ;
        RECT 1545.910 1491.430 1606.715 1491.730 ;
        RECT 1497.825 1491.415 1498.155 1491.430 ;
        RECT 1606.385 1491.415 1606.715 1491.430 ;
        RECT 1607.765 1491.730 1608.095 1491.745 ;
        RECT 1702.065 1491.730 1702.395 1491.745 ;
        RECT 1607.765 1491.430 1641.890 1491.730 ;
        RECT 1607.765 1491.415 1608.095 1491.430 ;
        RECT 1321.430 1490.750 1345.650 1491.050 ;
        RECT 1483.105 1491.050 1483.435 1491.065 ;
        RECT 1496.905 1491.050 1497.235 1491.065 ;
        RECT 1483.105 1490.750 1497.235 1491.050 ;
        RECT 1641.590 1491.050 1641.890 1491.430 ;
        RECT 1656.310 1491.430 1702.395 1491.730 ;
        RECT 1656.310 1491.050 1656.610 1491.430 ;
        RECT 1702.065 1491.415 1702.395 1491.430 ;
        RECT 1704.365 1491.730 1704.695 1491.745 ;
        RECT 1798.665 1491.730 1798.995 1491.745 ;
        RECT 1704.365 1491.430 1738.490 1491.730 ;
        RECT 1704.365 1491.415 1704.695 1491.430 ;
        RECT 1641.590 1490.750 1656.610 1491.050 ;
        RECT 1738.190 1491.050 1738.490 1491.430 ;
        RECT 1752.910 1491.430 1798.995 1491.730 ;
        RECT 1752.910 1491.050 1753.210 1491.430 ;
        RECT 1798.665 1491.415 1798.995 1491.430 ;
        RECT 1801.885 1491.730 1802.215 1491.745 ;
        RECT 1895.265 1491.730 1895.595 1491.745 ;
        RECT 1801.885 1491.430 1835.090 1491.730 ;
        RECT 1801.885 1491.415 1802.215 1491.430 ;
        RECT 1738.190 1490.750 1753.210 1491.050 ;
        RECT 1834.790 1491.050 1835.090 1491.430 ;
        RECT 1849.510 1491.430 1895.595 1491.730 ;
        RECT 1849.510 1491.050 1849.810 1491.430 ;
        RECT 1895.265 1491.415 1895.595 1491.430 ;
        RECT 2028.205 1491.730 2028.535 1491.745 ;
        RECT 2028.910 1491.730 2029.210 1492.790 ;
        RECT 2052.585 1492.775 2052.915 1492.790 ;
        RECT 2124.805 1492.410 2125.135 1492.425 ;
        RECT 2124.805 1492.110 2159.850 1492.410 ;
        RECT 2124.805 1492.095 2125.135 1492.110 ;
        RECT 2090.305 1491.730 2090.635 1491.745 ;
        RECT 2028.205 1491.430 2029.210 1491.730 ;
        RECT 2076.750 1491.430 2090.635 1491.730 ;
        RECT 2159.550 1491.730 2159.850 1492.110 ;
        RECT 2208.310 1492.110 2256.450 1492.410 ;
        RECT 2159.550 1491.430 2207.690 1491.730 ;
        RECT 2028.205 1491.415 2028.535 1491.430 ;
        RECT 1932.065 1491.050 1932.395 1491.065 ;
        RECT 1834.790 1490.750 1849.810 1491.050 ;
        RECT 1931.390 1490.750 1932.395 1491.050 ;
        RECT 1483.105 1490.735 1483.435 1490.750 ;
        RECT 1496.905 1490.735 1497.235 1490.750 ;
        RECT 1895.265 1489.690 1895.595 1489.705 ;
        RECT 1931.390 1489.690 1931.690 1490.750 ;
        RECT 1932.065 1490.735 1932.395 1490.750 ;
        RECT 2052.585 1491.050 2052.915 1491.065 ;
        RECT 2076.750 1491.050 2077.050 1491.430 ;
        RECT 2090.305 1491.415 2090.635 1491.430 ;
        RECT 2052.585 1490.750 2077.050 1491.050 ;
        RECT 2207.390 1491.050 2207.690 1491.430 ;
        RECT 2208.310 1491.050 2208.610 1492.110 ;
        RECT 2256.150 1491.730 2256.450 1492.110 ;
        RECT 2304.910 1492.110 2353.050 1492.410 ;
        RECT 2256.150 1491.430 2304.290 1491.730 ;
        RECT 2207.390 1490.750 2208.610 1491.050 ;
        RECT 2303.990 1491.050 2304.290 1491.430 ;
        RECT 2304.910 1491.050 2305.210 1492.110 ;
        RECT 2352.750 1491.730 2353.050 1492.110 ;
        RECT 2401.510 1492.110 2449.650 1492.410 ;
        RECT 2352.750 1491.430 2400.890 1491.730 ;
        RECT 2303.990 1490.750 2305.210 1491.050 ;
        RECT 2400.590 1491.050 2400.890 1491.430 ;
        RECT 2401.510 1491.050 2401.810 1492.110 ;
        RECT 2449.350 1491.730 2449.650 1492.110 ;
        RECT 2498.110 1492.110 2546.250 1492.410 ;
        RECT 2449.350 1491.430 2497.490 1491.730 ;
        RECT 2400.590 1490.750 2401.810 1491.050 ;
        RECT 2497.190 1491.050 2497.490 1491.430 ;
        RECT 2498.110 1491.050 2498.410 1492.110 ;
        RECT 2545.950 1491.730 2546.250 1492.110 ;
        RECT 2594.710 1492.110 2642.850 1492.410 ;
        RECT 2545.950 1491.430 2594.090 1491.730 ;
        RECT 2497.190 1490.750 2498.410 1491.050 ;
        RECT 2593.790 1491.050 2594.090 1491.430 ;
        RECT 2594.710 1491.050 2595.010 1492.110 ;
        RECT 2642.550 1491.730 2642.850 1492.110 ;
        RECT 2691.310 1492.110 2739.450 1492.410 ;
        RECT 2642.550 1491.430 2690.690 1491.730 ;
        RECT 2593.790 1490.750 2595.010 1491.050 ;
        RECT 2690.390 1491.050 2690.690 1491.430 ;
        RECT 2691.310 1491.050 2691.610 1492.110 ;
        RECT 2739.150 1491.730 2739.450 1492.110 ;
        RECT 2787.910 1492.110 2836.050 1492.410 ;
        RECT 2739.150 1491.430 2787.290 1491.730 ;
        RECT 2690.390 1490.750 2691.610 1491.050 ;
        RECT 2786.990 1491.050 2787.290 1491.430 ;
        RECT 2787.910 1491.050 2788.210 1492.110 ;
        RECT 2835.750 1491.730 2836.050 1492.110 ;
        RECT 2916.710 1491.730 2917.010 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2835.750 1491.430 2883.890 1491.730 ;
        RECT 2786.990 1490.750 2788.210 1491.050 ;
        RECT 2883.590 1491.050 2883.890 1491.430 ;
        RECT 2884.510 1491.430 2917.010 1491.730 ;
        RECT 2884.510 1491.050 2884.810 1491.430 ;
        RECT 2883.590 1490.750 2884.810 1491.050 ;
        RECT 2052.585 1490.735 2052.915 1490.750 ;
        RECT 1895.265 1489.390 1931.690 1489.690 ;
        RECT 1895.265 1489.375 1895.595 1489.390 ;
      LAYER via3 ;
        RECT 1275.420 2497.820 1275.740 2498.140 ;
        RECT 1980.140 1493.460 1980.460 1493.780 ;
        RECT 1435.500 1492.780 1435.820 1493.100 ;
        RECT 1275.420 1492.100 1275.740 1492.420 ;
        RECT 1435.500 1491.420 1435.820 1491.740 ;
        RECT 1980.140 1492.100 1980.460 1492.420 ;
      LAYER met4 ;
        RECT 1275.415 2497.815 1275.745 2498.145 ;
        RECT 1275.430 1492.425 1275.730 2497.815 ;
        RECT 1980.135 1493.455 1980.465 1493.785 ;
        RECT 1435.495 1492.775 1435.825 1493.105 ;
        RECT 1275.415 1492.095 1275.745 1492.425 ;
        RECT 1435.510 1491.745 1435.810 1492.775 ;
        RECT 1980.150 1492.425 1980.450 1493.455 ;
        RECT 1980.135 1492.095 1980.465 1492.425 ;
        RECT 1435.495 1491.415 1435.825 1491.745 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1293.130 2496.320 1293.450 2496.580 ;
        RECT 1293.220 2495.500 1293.360 2496.320 ;
        RECT 2901.290 2495.500 2901.610 2495.560 ;
        RECT 1293.220 2495.360 2901.610 2495.500 ;
        RECT 2901.290 2495.300 2901.610 2495.360 ;
      LAYER via ;
        RECT 1293.160 2496.320 1293.420 2496.580 ;
        RECT 2901.320 2495.300 2901.580 2495.560 ;
      LAYER met2 ;
        RECT 1291.770 2496.690 1292.050 2500.000 ;
        RECT 1291.770 2496.610 1293.360 2496.690 ;
        RECT 1291.770 2496.550 1293.420 2496.610 ;
        RECT 1291.770 2496.000 1292.050 2496.550 ;
        RECT 1293.160 2496.290 1293.420 2496.550 ;
        RECT 2901.320 2495.270 2901.580 2495.590 ;
        RECT 2901.380 1730.445 2901.520 2495.270 ;
        RECT 2901.310 1730.075 2901.590 1730.445 ;
      LAYER via2 ;
        RECT 2901.310 1730.120 2901.590 1730.400 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1729.660 2924.800 1730.860 ;
=======
        RECT 2901.285 1730.410 2901.615 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2901.285 1730.110 2924.800 1730.410 ;
        RECT 2901.285 1730.095 2901.615 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1311.530 2515.560 1311.850 2515.620 ;
        RECT 1950.010 2515.560 1950.330 2515.620 ;
        RECT 1311.530 2515.420 1950.330 2515.560 ;
        RECT 1311.530 2515.360 1311.850 2515.420 ;
        RECT 1950.010 2515.360 1950.330 2515.420 ;
        RECT 1950.010 1966.460 1950.330 1966.520 ;
        RECT 2898.070 1966.460 2898.390 1966.520 ;
        RECT 1950.010 1966.320 2898.390 1966.460 ;
        RECT 1950.010 1966.260 1950.330 1966.320 ;
        RECT 2898.070 1966.260 2898.390 1966.320 ;
      LAYER via ;
        RECT 1311.560 2515.360 1311.820 2515.620 ;
        RECT 1950.040 2515.360 1950.300 2515.620 ;
        RECT 1950.040 1966.260 1950.300 1966.520 ;
        RECT 2898.100 1966.260 2898.360 1966.520 ;
      LAYER met2 ;
        RECT 1311.560 2515.330 1311.820 2515.650 ;
        RECT 1950.040 2515.330 1950.300 2515.650 ;
        RECT 1311.620 2500.000 1311.760 2515.330 ;
        RECT 1311.550 2496.000 1311.830 2500.000 ;
        RECT 1950.100 1966.550 1950.240 2515.330 ;
        RECT 1950.040 1966.230 1950.300 1966.550 ;
        RECT 2898.100 1966.230 2898.360 1966.550 ;
        RECT 2898.160 1965.045 2898.300 1966.230 ;
        RECT 2898.090 1964.675 2898.370 1965.045 ;
      LAYER via2 ;
        RECT 2898.090 1964.720 2898.370 1965.000 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1964.260 2924.800 1965.460 ;
=======
        RECT 2898.065 1965.010 2898.395 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2898.065 1964.710 2924.800 1965.010 ;
        RECT 2898.065 1964.695 2898.395 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1932.145 2514.385 1932.315 2516.595 ;
      LAYER mcon ;
        RECT 1932.145 2516.425 1932.315 2516.595 ;
      LAYER met1 ;
        RECT 1331.770 2516.580 1332.090 2516.640 ;
        RECT 1932.085 2516.580 1932.375 2516.625 ;
        RECT 1331.770 2516.440 1932.375 2516.580 ;
        RECT 1331.770 2516.380 1332.090 2516.440 ;
        RECT 1932.085 2516.395 1932.375 2516.440 ;
        RECT 1932.085 2514.540 1932.375 2514.585 ;
        RECT 1951.850 2514.540 1952.170 2514.600 ;
        RECT 1932.085 2514.400 1952.170 2514.540 ;
        RECT 1932.085 2514.355 1932.375 2514.400 ;
        RECT 1951.850 2514.340 1952.170 2514.400 ;
        RECT 1951.850 2201.060 1952.170 2201.120 ;
        RECT 2898.070 2201.060 2898.390 2201.120 ;
        RECT 1951.850 2200.920 2898.390 2201.060 ;
        RECT 1951.850 2200.860 1952.170 2200.920 ;
        RECT 2898.070 2200.860 2898.390 2200.920 ;
      LAYER via ;
        RECT 1331.800 2516.380 1332.060 2516.640 ;
        RECT 1951.880 2514.340 1952.140 2514.600 ;
        RECT 1951.880 2200.860 1952.140 2201.120 ;
        RECT 2898.100 2200.860 2898.360 2201.120 ;
      LAYER met2 ;
        RECT 1331.800 2516.350 1332.060 2516.670 ;
        RECT 1331.860 2500.000 1332.000 2516.350 ;
        RECT 1951.880 2514.310 1952.140 2514.630 ;
        RECT 1331.790 2496.000 1332.070 2500.000 ;
        RECT 1951.940 2201.150 1952.080 2514.310 ;
        RECT 1951.880 2200.830 1952.140 2201.150 ;
        RECT 2898.100 2200.830 2898.360 2201.150 ;
        RECT 2898.160 2199.645 2898.300 2200.830 ;
        RECT 2898.090 2199.275 2898.370 2199.645 ;
      LAYER via2 ;
        RECT 2898.090 2199.320 2898.370 2199.600 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2198.860 2924.800 2200.060 ;
=======
        RECT 2898.065 2199.610 2898.395 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2898.065 2199.310 2924.800 2199.610 ;
        RECT 2898.065 2199.295 2898.395 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1798.670 201.180 1798.990 201.240 ;
        RECT 1811.550 201.180 1811.870 201.240 ;
        RECT 1798.670 201.040 1811.870 201.180 ;
        RECT 1798.670 200.980 1798.990 201.040 ;
        RECT 1811.550 200.980 1811.870 201.040 ;
        RECT 2090.310 201.180 2090.630 201.240 ;
        RECT 2124.810 201.180 2125.130 201.240 ;
        RECT 2090.310 201.040 2125.130 201.180 ;
        RECT 2090.310 200.980 2090.630 201.040 ;
        RECT 2124.810 200.980 2125.130 201.040 ;
        RECT 1606.390 200.840 1606.710 200.900 ;
        RECT 1607.770 200.840 1608.090 200.900 ;
        RECT 1606.390 200.700 1608.090 200.840 ;
        RECT 1606.390 200.640 1606.710 200.700 ;
        RECT 1607.770 200.640 1608.090 200.700 ;
        RECT 1702.070 200.840 1702.390 200.900 ;
        RECT 1714.490 200.840 1714.810 200.900 ;
        RECT 1702.070 200.700 1714.810 200.840 ;
        RECT 1702.070 200.640 1702.390 200.700 ;
        RECT 1714.490 200.640 1714.810 200.700 ;
        RECT 1932.070 200.500 1932.390 200.560 ;
        RECT 1946.330 200.500 1946.650 200.560 ;
        RECT 1932.070 200.360 1946.650 200.500 ;
        RECT 1932.070 200.300 1932.390 200.360 ;
        RECT 1946.330 200.300 1946.650 200.360 ;
      LAYER via ;
        RECT 1798.700 200.980 1798.960 201.240 ;
        RECT 1811.580 200.980 1811.840 201.240 ;
        RECT 2090.340 200.980 2090.600 201.240 ;
        RECT 2124.840 200.980 2125.100 201.240 ;
        RECT 1606.420 200.640 1606.680 200.900 ;
        RECT 1607.800 200.640 1608.060 200.900 ;
        RECT 1702.100 200.640 1702.360 200.900 ;
        RECT 1714.520 200.640 1714.780 200.900 ;
        RECT 1932.100 200.300 1932.360 200.560 ;
        RECT 1946.360 200.300 1946.620 200.560 ;
      LAYER met2 ;
        RECT 1159.750 2498.050 1160.030 2500.000 ;
        RECT 1161.590 2498.050 1161.870 2498.165 ;
        RECT 1159.750 2497.910 1161.870 2498.050 ;
        RECT 1159.750 2496.000 1160.030 2497.910 ;
        RECT 1161.590 2497.795 1161.870 2497.910 ;
        RECT 1200.230 217.755 1200.510 218.125 ;
        RECT 1200.300 201.125 1200.440 217.755 ;
        RECT 2028.230 202.795 2028.510 203.165 ;
        RECT 1532.350 201.435 1532.630 201.805 ;
        RECT 1946.350 201.435 1946.630 201.805 ;
        RECT 1532.420 201.125 1532.560 201.435 ;
        RECT 1798.700 201.125 1798.960 201.270 ;
        RECT 1811.580 201.125 1811.840 201.270 ;
        RECT 1200.230 200.755 1200.510 201.125 ;
        RECT 1297.290 200.755 1297.570 201.125 ;
        RECT 1393.430 200.755 1393.710 201.125 ;
        RECT 1532.350 200.755 1532.630 201.125 ;
        RECT 1606.410 200.755 1606.690 201.125 ;
        RECT 1607.790 200.755 1608.070 201.125 ;
        RECT 1702.090 200.755 1702.370 201.125 ;
        RECT 1714.510 200.755 1714.790 201.125 ;
        RECT 1798.690 200.755 1798.970 201.125 ;
        RECT 1811.570 200.755 1811.850 201.125 ;
        RECT 1895.290 200.755 1895.570 201.125 ;
        RECT 1297.360 200.445 1297.500 200.755 ;
        RECT 1297.290 200.075 1297.570 200.445 ;
        RECT 1393.500 199.085 1393.640 200.755 ;
        RECT 1606.420 200.610 1606.680 200.755 ;
        RECT 1607.800 200.610 1608.060 200.755 ;
        RECT 1702.100 200.610 1702.360 200.755 ;
        RECT 1714.520 200.610 1714.780 200.755 ;
        RECT 1895.360 199.085 1895.500 200.755 ;
        RECT 1946.420 200.590 1946.560 201.435 ;
        RECT 2028.300 201.125 2028.440 202.795 ;
        RECT 2052.610 202.115 2052.890 202.485 ;
        RECT 2028.230 200.755 2028.510 201.125 ;
        RECT 1932.100 200.445 1932.360 200.590 ;
        RECT 1932.090 200.075 1932.370 200.445 ;
        RECT 1946.360 200.270 1946.620 200.590 ;
        RECT 2052.680 200.445 2052.820 202.115 ;
        RECT 2124.830 201.435 2125.110 201.805 ;
        RECT 2124.900 201.270 2125.040 201.435 ;
        RECT 2090.340 201.125 2090.600 201.270 ;
        RECT 2090.330 200.755 2090.610 201.125 ;
        RECT 2124.840 200.950 2125.100 201.270 ;
        RECT 2052.610 200.075 2052.890 200.445 ;
        RECT 1393.430 198.715 1393.710 199.085 ;
        RECT 1895.290 198.715 1895.570 199.085 ;
      LAYER via2 ;
        RECT 1161.590 2497.840 1161.870 2498.120 ;
        RECT 1200.230 217.800 1200.510 218.080 ;
        RECT 2028.230 202.840 2028.510 203.120 ;
        RECT 1532.350 201.480 1532.630 201.760 ;
        RECT 1946.350 201.480 1946.630 201.760 ;
        RECT 1200.230 200.800 1200.510 201.080 ;
        RECT 1297.290 200.800 1297.570 201.080 ;
        RECT 1393.430 200.800 1393.710 201.080 ;
        RECT 1532.350 200.800 1532.630 201.080 ;
        RECT 1606.410 200.800 1606.690 201.080 ;
        RECT 1607.790 200.800 1608.070 201.080 ;
        RECT 1702.090 200.800 1702.370 201.080 ;
        RECT 1714.510 200.800 1714.790 201.080 ;
        RECT 1798.690 200.800 1798.970 201.080 ;
        RECT 1811.570 200.800 1811.850 201.080 ;
        RECT 1895.290 200.800 1895.570 201.080 ;
        RECT 1297.290 200.120 1297.570 200.400 ;
        RECT 2052.610 202.160 2052.890 202.440 ;
        RECT 2028.230 200.800 2028.510 201.080 ;
        RECT 1932.090 200.120 1932.370 200.400 ;
        RECT 2124.830 201.480 2125.110 201.760 ;
        RECT 2090.330 200.800 2090.610 201.080 ;
        RECT 2052.610 200.120 2052.890 200.400 ;
        RECT 1393.430 198.760 1393.710 199.040 ;
        RECT 1895.290 198.760 1895.570 199.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 204.420 2924.800 205.620 ;
=======
        RECT 1161.565 2498.130 1161.895 2498.145 ;
        RECT 1164.990 2498.130 1165.370 2498.140 ;
        RECT 1161.565 2497.830 1165.370 2498.130 ;
        RECT 1161.565 2497.815 1161.895 2497.830 ;
        RECT 1164.990 2497.820 1165.370 2497.830 ;
        RECT 1164.990 218.090 1165.370 218.100 ;
        RECT 1200.205 218.090 1200.535 218.105 ;
        RECT 1164.990 217.790 1200.535 218.090 ;
        RECT 1164.990 217.780 1165.370 217.790 ;
        RECT 1200.205 217.775 1200.535 217.790 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2916.710 204.870 2924.800 205.170 ;
        RECT 1980.110 203.130 1980.490 203.140 ;
        RECT 2028.205 203.130 2028.535 203.145 ;
        RECT 1980.110 202.830 2028.535 203.130 ;
        RECT 1980.110 202.820 1980.490 202.830 ;
        RECT 2028.205 202.815 2028.535 202.830 ;
        RECT 2052.585 202.450 2052.915 202.465 ;
        RECT 2028.910 202.150 2052.915 202.450 ;
        RECT 1248.710 201.770 1249.090 201.780 ;
        RECT 1532.325 201.770 1532.655 201.785 ;
        RECT 1248.710 201.470 1249.970 201.770 ;
        RECT 1248.710 201.460 1249.090 201.470 ;
        RECT 1200.205 201.090 1200.535 201.105 ;
        RECT 1249.670 201.090 1249.970 201.470 ;
        RECT 1441.030 201.470 1442.250 201.770 ;
        RECT 1297.265 201.090 1297.595 201.105 ;
        RECT 1200.205 200.790 1201.210 201.090 ;
        RECT 1249.670 200.790 1297.595 201.090 ;
        RECT 1200.205 200.775 1200.535 200.790 ;
        RECT 1200.910 200.410 1201.210 200.790 ;
        RECT 1297.265 200.775 1297.595 200.790 ;
        RECT 1393.405 201.090 1393.735 201.105 ;
        RECT 1441.030 201.090 1441.330 201.470 ;
        RECT 1393.405 200.790 1441.330 201.090 ;
        RECT 1441.950 201.090 1442.250 201.470 ;
        RECT 1459.430 201.470 1532.655 201.770 ;
        RECT 1459.430 201.090 1459.730 201.470 ;
        RECT 1532.325 201.455 1532.655 201.470 ;
        RECT 1946.325 201.770 1946.655 201.785 ;
        RECT 1980.110 201.770 1980.490 201.780 ;
        RECT 1946.325 201.470 1980.490 201.770 ;
        RECT 1946.325 201.455 1946.655 201.470 ;
        RECT 1980.110 201.460 1980.490 201.470 ;
        RECT 1441.950 200.790 1459.730 201.090 ;
        RECT 1532.325 201.090 1532.655 201.105 ;
        RECT 1606.385 201.090 1606.715 201.105 ;
        RECT 1532.325 200.790 1606.715 201.090 ;
        RECT 1393.405 200.775 1393.735 200.790 ;
        RECT 1532.325 200.775 1532.655 200.790 ;
        RECT 1606.385 200.775 1606.715 200.790 ;
        RECT 1607.765 201.090 1608.095 201.105 ;
        RECT 1702.065 201.090 1702.395 201.105 ;
        RECT 1607.765 200.790 1641.890 201.090 ;
        RECT 1607.765 200.775 1608.095 200.790 ;
        RECT 1248.710 200.410 1249.090 200.420 ;
        RECT 1200.910 200.110 1249.090 200.410 ;
        RECT 1248.710 200.100 1249.090 200.110 ;
        RECT 1297.265 200.410 1297.595 200.425 ;
        RECT 1345.310 200.410 1345.690 200.420 ;
        RECT 1297.265 200.110 1345.690 200.410 ;
        RECT 1641.590 200.410 1641.890 200.790 ;
        RECT 1656.310 200.790 1702.395 201.090 ;
        RECT 1656.310 200.410 1656.610 200.790 ;
        RECT 1702.065 200.775 1702.395 200.790 ;
        RECT 1714.485 201.090 1714.815 201.105 ;
        RECT 1798.665 201.090 1798.995 201.105 ;
        RECT 1714.485 200.790 1738.490 201.090 ;
        RECT 1714.485 200.775 1714.815 200.790 ;
        RECT 1641.590 200.110 1656.610 200.410 ;
        RECT 1738.190 200.410 1738.490 200.790 ;
        RECT 1752.910 200.790 1798.995 201.090 ;
        RECT 1752.910 200.410 1753.210 200.790 ;
        RECT 1798.665 200.775 1798.995 200.790 ;
        RECT 1811.545 201.090 1811.875 201.105 ;
        RECT 1895.265 201.090 1895.595 201.105 ;
        RECT 1811.545 200.790 1835.090 201.090 ;
        RECT 1811.545 200.775 1811.875 200.790 ;
        RECT 1738.190 200.110 1753.210 200.410 ;
        RECT 1834.790 200.410 1835.090 200.790 ;
        RECT 1849.510 200.790 1895.595 201.090 ;
        RECT 1849.510 200.410 1849.810 200.790 ;
        RECT 1895.265 200.775 1895.595 200.790 ;
        RECT 2028.205 201.090 2028.535 201.105 ;
        RECT 2028.910 201.090 2029.210 202.150 ;
        RECT 2052.585 202.135 2052.915 202.150 ;
        RECT 2124.805 201.770 2125.135 201.785 ;
        RECT 2124.805 201.470 2159.850 201.770 ;
        RECT 2124.805 201.455 2125.135 201.470 ;
        RECT 2090.305 201.090 2090.635 201.105 ;
        RECT 2028.205 200.790 2029.210 201.090 ;
        RECT 2076.750 200.790 2090.635 201.090 ;
        RECT 2159.550 201.090 2159.850 201.470 ;
        RECT 2208.310 201.470 2256.450 201.770 ;
        RECT 2159.550 200.790 2207.690 201.090 ;
        RECT 2028.205 200.775 2028.535 200.790 ;
        RECT 1932.065 200.410 1932.395 200.425 ;
        RECT 1834.790 200.110 1849.810 200.410 ;
        RECT 1931.390 200.110 1932.395 200.410 ;
        RECT 1297.265 200.095 1297.595 200.110 ;
        RECT 1345.310 200.100 1345.690 200.110 ;
        RECT 1345.310 199.050 1345.690 199.060 ;
        RECT 1393.405 199.050 1393.735 199.065 ;
        RECT 1345.310 198.750 1393.735 199.050 ;
        RECT 1345.310 198.740 1345.690 198.750 ;
        RECT 1393.405 198.735 1393.735 198.750 ;
        RECT 1895.265 199.050 1895.595 199.065 ;
        RECT 1931.390 199.050 1931.690 200.110 ;
        RECT 1932.065 200.095 1932.395 200.110 ;
        RECT 2052.585 200.410 2052.915 200.425 ;
        RECT 2076.750 200.410 2077.050 200.790 ;
        RECT 2090.305 200.775 2090.635 200.790 ;
        RECT 2052.585 200.110 2077.050 200.410 ;
        RECT 2207.390 200.410 2207.690 200.790 ;
        RECT 2208.310 200.410 2208.610 201.470 ;
        RECT 2256.150 201.090 2256.450 201.470 ;
        RECT 2304.910 201.470 2353.050 201.770 ;
        RECT 2256.150 200.790 2304.290 201.090 ;
        RECT 2207.390 200.110 2208.610 200.410 ;
        RECT 2303.990 200.410 2304.290 200.790 ;
        RECT 2304.910 200.410 2305.210 201.470 ;
        RECT 2352.750 201.090 2353.050 201.470 ;
        RECT 2401.510 201.470 2449.650 201.770 ;
        RECT 2352.750 200.790 2400.890 201.090 ;
        RECT 2303.990 200.110 2305.210 200.410 ;
        RECT 2400.590 200.410 2400.890 200.790 ;
        RECT 2401.510 200.410 2401.810 201.470 ;
        RECT 2449.350 201.090 2449.650 201.470 ;
        RECT 2498.110 201.470 2546.250 201.770 ;
        RECT 2449.350 200.790 2497.490 201.090 ;
        RECT 2400.590 200.110 2401.810 200.410 ;
        RECT 2497.190 200.410 2497.490 200.790 ;
        RECT 2498.110 200.410 2498.410 201.470 ;
        RECT 2545.950 201.090 2546.250 201.470 ;
        RECT 2594.710 201.470 2642.850 201.770 ;
        RECT 2545.950 200.790 2594.090 201.090 ;
        RECT 2497.190 200.110 2498.410 200.410 ;
        RECT 2593.790 200.410 2594.090 200.790 ;
        RECT 2594.710 200.410 2595.010 201.470 ;
        RECT 2642.550 201.090 2642.850 201.470 ;
        RECT 2691.310 201.470 2739.450 201.770 ;
        RECT 2642.550 200.790 2690.690 201.090 ;
        RECT 2593.790 200.110 2595.010 200.410 ;
        RECT 2690.390 200.410 2690.690 200.790 ;
        RECT 2691.310 200.410 2691.610 201.470 ;
        RECT 2739.150 201.090 2739.450 201.470 ;
        RECT 2787.910 201.470 2836.050 201.770 ;
        RECT 2739.150 200.790 2787.290 201.090 ;
        RECT 2690.390 200.110 2691.610 200.410 ;
        RECT 2786.990 200.410 2787.290 200.790 ;
        RECT 2787.910 200.410 2788.210 201.470 ;
        RECT 2835.750 201.090 2836.050 201.470 ;
        RECT 2916.710 201.090 2917.010 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2835.750 200.790 2883.890 201.090 ;
        RECT 2786.990 200.110 2788.210 200.410 ;
        RECT 2883.590 200.410 2883.890 200.790 ;
        RECT 2884.510 200.790 2917.010 201.090 ;
        RECT 2884.510 200.410 2884.810 200.790 ;
        RECT 2883.590 200.110 2884.810 200.410 ;
        RECT 2052.585 200.095 2052.915 200.110 ;
        RECT 1895.265 198.750 1931.690 199.050 ;
        RECT 1895.265 198.735 1895.595 198.750 ;
      LAYER via3 ;
        RECT 1165.020 2497.820 1165.340 2498.140 ;
        RECT 1165.020 217.780 1165.340 218.100 ;
        RECT 1980.140 202.820 1980.460 203.140 ;
        RECT 1248.740 201.460 1249.060 201.780 ;
        RECT 1980.140 201.460 1980.460 201.780 ;
        RECT 1248.740 200.100 1249.060 200.420 ;
        RECT 1345.340 200.100 1345.660 200.420 ;
        RECT 1345.340 198.740 1345.660 199.060 ;
      LAYER met4 ;
        RECT 1165.015 2497.815 1165.345 2498.145 ;
        RECT 1165.030 218.105 1165.330 2497.815 ;
        RECT 1165.015 217.775 1165.345 218.105 ;
        RECT 1980.135 202.815 1980.465 203.145 ;
        RECT 1980.150 201.785 1980.450 202.815 ;
        RECT 1248.735 201.455 1249.065 201.785 ;
        RECT 1980.135 201.455 1980.465 201.785 ;
        RECT 1248.750 200.425 1249.050 201.455 ;
        RECT 1248.735 200.095 1249.065 200.425 ;
        RECT 1345.335 200.095 1345.665 200.425 ;
        RECT 1345.350 199.065 1345.650 200.095 ;
        RECT 1345.335 198.735 1345.665 199.065 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1352.470 2546.840 1352.790 2546.900 ;
        RECT 2900.830 2546.840 2901.150 2546.900 ;
        RECT 1352.470 2546.700 2901.150 2546.840 ;
        RECT 1352.470 2546.640 1352.790 2546.700 ;
        RECT 2900.830 2546.640 2901.150 2546.700 ;
        RECT 1352.470 2518.280 1352.790 2518.340 ;
        RECT 1357.990 2518.280 1358.310 2518.340 ;
        RECT 1352.470 2518.140 1358.310 2518.280 ;
        RECT 1352.470 2518.080 1352.790 2518.140 ;
        RECT 1357.990 2518.080 1358.310 2518.140 ;
      LAYER via ;
        RECT 1352.500 2546.640 1352.760 2546.900 ;
        RECT 2900.860 2546.640 2901.120 2546.900 ;
        RECT 1352.500 2518.080 1352.760 2518.340 ;
        RECT 1358.020 2518.080 1358.280 2518.340 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.930 2901.060 2551.515 ;
        RECT 1352.500 2546.610 1352.760 2546.930 ;
        RECT 2900.860 2546.610 2901.120 2546.930 ;
        RECT 1352.560 2518.370 1352.700 2546.610 ;
        RECT 1352.500 2518.050 1352.760 2518.370 ;
        RECT 1358.020 2518.050 1358.280 2518.370 ;
        RECT 1358.080 2500.000 1358.220 2518.050 ;
        RECT 1358.010 2496.000 1358.290 2500.000 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2551.100 2924.800 2552.300 ;
=======
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1379.610 2781.100 1379.930 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 1379.610 2780.960 2901.150 2781.100 ;
        RECT 1379.610 2780.900 1379.930 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 1379.640 2780.900 1379.900 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 1379.640 2780.870 1379.900 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 1377.790 2499.410 1378.070 2500.000 ;
        RECT 1379.700 2499.410 1379.840 2780.870 ;
        RECT 1377.790 2499.270 1379.840 2499.410 ;
        RECT 1377.790 2496.000 1378.070 2499.270 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2785.700 2924.800 2786.900 ;
=======
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1400.310 3015.700 1400.630 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 1400.310 3015.560 2901.150 3015.700 ;
        RECT 1400.310 3015.500 1400.630 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 1400.340 3015.500 1400.600 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 1400.340 3015.470 1400.600 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 1397.570 2498.730 1397.850 2500.000 ;
        RECT 1400.400 2499.410 1400.540 3015.470 ;
        RECT 1399.940 2499.270 1400.540 2499.410 ;
        RECT 1399.940 2498.730 1400.080 2499.270 ;
        RECT 1397.570 2498.590 1400.080 2498.730 ;
        RECT 1397.570 2496.000 1397.850 2498.590 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3020.300 2924.800 3021.500 ;
=======
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1420.550 3250.300 1420.870 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1420.550 3250.160 2901.150 3250.300 ;
        RECT 1420.550 3250.100 1420.870 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 1420.580 3250.100 1420.840 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1420.580 3250.070 1420.840 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1420.640 2500.090 1420.780 3250.070 ;
        RECT 1417.350 2499.410 1417.630 2500.000 ;
        RECT 1419.720 2499.950 1420.780 2500.090 ;
        RECT 1419.720 2499.410 1419.860 2499.950 ;
        RECT 1417.350 2499.270 1419.860 2499.410 ;
        RECT 1417.350 2496.000 1417.630 2499.270 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3254.900 2924.800 3256.100 ;
=======
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1441.710 3484.900 1442.030 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1441.710 3484.760 2901.150 3484.900 ;
        RECT 1441.710 3484.700 1442.030 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 1437.110 2514.880 1437.430 2514.940 ;
        RECT 1441.710 2514.880 1442.030 2514.940 ;
        RECT 1437.110 2514.740 1442.030 2514.880 ;
        RECT 1437.110 2514.680 1437.430 2514.740 ;
        RECT 1441.710 2514.680 1442.030 2514.740 ;
      LAYER via ;
        RECT 1441.740 3484.700 1442.000 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 1437.140 2514.680 1437.400 2514.940 ;
        RECT 1441.740 2514.680 1442.000 2514.940 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1441.740 3484.670 1442.000 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1441.800 2514.970 1441.940 3484.670 ;
        RECT 1437.140 2514.650 1437.400 2514.970 ;
        RECT 1441.740 2514.650 1442.000 2514.970 ;
        RECT 1437.200 2500.000 1437.340 2514.650 ;
        RECT 1437.130 2496.000 1437.410 2500.000 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3489.500 2924.800 3490.700 ;
=======
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1462.410 3502.580 1462.730 3502.640 ;
        RECT 2635.870 3502.580 2636.190 3502.640 ;
        RECT 1462.410 3502.440 2636.190 3502.580 ;
        RECT 1462.410 3502.380 1462.730 3502.440 ;
        RECT 2635.870 3502.380 2636.190 3502.440 ;
        RECT 1457.350 2514.880 1457.670 2514.940 ;
        RECT 1462.410 2514.880 1462.730 2514.940 ;
        RECT 1457.350 2514.740 1462.730 2514.880 ;
        RECT 1457.350 2514.680 1457.670 2514.740 ;
        RECT 1462.410 2514.680 1462.730 2514.740 ;
      LAYER via ;
        RECT 1462.440 3502.380 1462.700 3502.640 ;
        RECT 2635.900 3502.380 2636.160 3502.640 ;
        RECT 1457.380 2514.680 1457.640 2514.940 ;
        RECT 1462.440 2514.680 1462.700 2514.940 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2635.750 3519.700 2636.310 3524.800 ;
=======
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3502.670 2636.100 3517.600 ;
        RECT 1462.440 3502.350 1462.700 3502.670 ;
        RECT 2635.900 3502.350 2636.160 3502.670 ;
        RECT 1462.500 2514.970 1462.640 3502.350 ;
        RECT 1457.380 2514.650 1457.640 2514.970 ;
        RECT 1462.440 2514.650 1462.700 2514.970 ;
        RECT 1457.440 2500.000 1457.580 2514.650 ;
        RECT 1457.370 2496.000 1457.650 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1483.110 3504.280 1483.430 3504.340 ;
        RECT 2311.570 3504.280 2311.890 3504.340 ;
        RECT 1483.110 3504.140 2311.890 3504.280 ;
        RECT 1483.110 3504.080 1483.430 3504.140 ;
        RECT 2311.570 3504.080 2311.890 3504.140 ;
        RECT 1477.130 2514.880 1477.450 2514.940 ;
        RECT 1483.110 2514.880 1483.430 2514.940 ;
        RECT 1477.130 2514.740 1483.430 2514.880 ;
        RECT 1477.130 2514.680 1477.450 2514.740 ;
        RECT 1483.110 2514.680 1483.430 2514.740 ;
      LAYER via ;
        RECT 1483.140 3504.080 1483.400 3504.340 ;
        RECT 2311.600 3504.080 2311.860 3504.340 ;
        RECT 1477.160 2514.680 1477.420 2514.940 ;
        RECT 1483.140 2514.680 1483.400 2514.940 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2311.450 3519.700 2312.010 3524.800 ;
=======
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3504.370 2311.800 3517.600 ;
        RECT 1483.140 3504.050 1483.400 3504.370 ;
        RECT 2311.600 3504.050 2311.860 3504.370 ;
        RECT 1483.200 2514.970 1483.340 3504.050 ;
        RECT 1477.160 2514.650 1477.420 2514.970 ;
        RECT 1483.140 2514.650 1483.400 2514.970 ;
        RECT 1477.220 2500.000 1477.360 2514.650 ;
        RECT 1477.150 2496.000 1477.430 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1496.910 3500.880 1497.230 3500.940 ;
        RECT 1987.270 3500.880 1987.590 3500.940 ;
        RECT 1496.910 3500.740 1987.590 3500.880 ;
        RECT 1496.910 3500.680 1497.230 3500.740 ;
        RECT 1987.270 3500.680 1987.590 3500.740 ;
      LAYER via ;
        RECT 1496.940 3500.680 1497.200 3500.940 ;
        RECT 1987.300 3500.680 1987.560 3500.940 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1987.150 3519.700 1987.710 3524.800 ;
=======
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3500.970 1987.500 3517.600 ;
        RECT 1496.940 3500.650 1497.200 3500.970 ;
        RECT 1987.300 3500.650 1987.560 3500.970 ;
        RECT 1497.000 2500.000 1497.140 3500.650 ;
        RECT 1496.930 2496.000 1497.210 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1517.610 3498.840 1517.930 3498.900 ;
        RECT 1662.510 3498.840 1662.830 3498.900 ;
        RECT 1517.610 3498.700 1662.830 3498.840 ;
        RECT 1517.610 3498.640 1517.930 3498.700 ;
        RECT 1662.510 3498.640 1662.830 3498.700 ;
      LAYER via ;
        RECT 1517.640 3498.640 1517.900 3498.900 ;
        RECT 1662.540 3498.640 1662.800 3498.900 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1662.390 3519.700 1662.950 3524.800 ;
=======
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3498.930 1662.740 3517.600 ;
        RECT 1517.640 3498.610 1517.900 3498.930 ;
        RECT 1662.540 3498.610 1662.800 3498.930 ;
        RECT 1516.710 2499.410 1516.990 2500.000 ;
        RECT 1517.700 2499.410 1517.840 3498.610 ;
        RECT 1516.710 2499.270 1517.840 2499.410 ;
        RECT 1516.710 2496.000 1516.990 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1524.125 3499.195 1524.295 3499.535 ;
        RECT 1524.125 3499.025 1525.675 3499.195 ;
      LAYER mcon ;
        RECT 1524.125 3499.365 1524.295 3499.535 ;
        RECT 1525.505 3499.025 1525.675 3499.195 ;
      LAYER met1 ;
        RECT 1524.065 3499.520 1524.355 3499.565 ;
        RECT 1500.220 3499.380 1524.355 3499.520 ;
        RECT 1338.210 3499.180 1338.530 3499.240 ;
        RECT 1500.220 3499.180 1500.360 3499.380 ;
        RECT 1524.065 3499.335 1524.355 3499.380 ;
        RECT 1338.210 3499.040 1500.360 3499.180 ;
        RECT 1525.445 3499.180 1525.735 3499.225 ;
        RECT 1528.190 3499.180 1528.510 3499.240 ;
        RECT 1525.445 3499.040 1528.510 3499.180 ;
        RECT 1338.210 3498.980 1338.530 3499.040 ;
        RECT 1525.445 3498.995 1525.735 3499.040 ;
        RECT 1528.190 3498.980 1528.510 3499.040 ;
        RECT 1528.190 2518.280 1528.510 2518.340 ;
        RECT 1534.630 2518.280 1534.950 2518.340 ;
        RECT 1528.190 2518.140 1534.950 2518.280 ;
        RECT 1528.190 2518.080 1528.510 2518.140 ;
        RECT 1534.630 2518.080 1534.950 2518.140 ;
      LAYER via ;
        RECT 1338.240 3498.980 1338.500 3499.240 ;
        RECT 1528.220 3498.980 1528.480 3499.240 ;
        RECT 1528.220 2518.080 1528.480 2518.340 ;
        RECT 1534.660 2518.080 1534.920 2518.340 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1338.090 3519.700 1338.650 3524.800 ;
=======
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3499.270 1338.440 3517.600 ;
        RECT 1338.240 3498.950 1338.500 3499.270 ;
        RECT 1528.220 3498.950 1528.480 3499.270 ;
        RECT 1528.280 2518.370 1528.420 3498.950 ;
        RECT 1528.220 2518.050 1528.480 2518.370 ;
        RECT 1534.660 2518.050 1534.920 2518.370 ;
        RECT 1534.720 2499.410 1534.860 2518.050 ;
        RECT 1536.490 2499.410 1536.770 2500.000 ;
        RECT 1534.720 2499.270 1536.770 2499.410 ;
        RECT 1536.490 2496.000 1536.770 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2090.310 435.780 2090.630 435.840 ;
        RECT 2124.810 435.780 2125.130 435.840 ;
        RECT 2090.310 435.640 2125.130 435.780 ;
        RECT 2090.310 435.580 2090.630 435.640 ;
        RECT 2124.810 435.580 2125.130 435.640 ;
        RECT 1895.270 435.440 1895.590 435.500 ;
        RECT 1930.230 435.440 1930.550 435.500 ;
        RECT 1895.270 435.300 1930.550 435.440 ;
        RECT 1895.270 435.240 1895.590 435.300 ;
        RECT 1930.230 435.240 1930.550 435.300 ;
        RECT 1932.070 435.100 1932.390 435.160 ;
        RECT 1956.450 435.100 1956.770 435.160 ;
        RECT 1932.070 434.960 1956.770 435.100 ;
        RECT 1932.070 434.900 1932.390 434.960 ;
        RECT 1956.450 434.900 1956.770 434.960 ;
        RECT 2042.010 434.760 2042.330 434.820 ;
        RECT 2069.610 434.760 2069.930 434.820 ;
        RECT 2042.010 434.620 2069.930 434.760 ;
        RECT 2042.010 434.560 2042.330 434.620 ;
        RECT 2069.610 434.560 2069.930 434.620 ;
      LAYER via ;
        RECT 2090.340 435.580 2090.600 435.840 ;
        RECT 2124.840 435.580 2125.100 435.840 ;
        RECT 1895.300 435.240 1895.560 435.500 ;
        RECT 1930.260 435.240 1930.520 435.500 ;
        RECT 1932.100 434.900 1932.360 435.160 ;
        RECT 1956.480 434.900 1956.740 435.160 ;
        RECT 2042.040 434.560 2042.300 434.820 ;
        RECT 2069.640 434.560 2069.900 434.820 ;
      LAYER met2 ;
        RECT 1178.150 2498.050 1178.430 2498.165 ;
        RECT 1179.530 2498.050 1179.810 2500.000 ;
        RECT 1178.150 2497.910 1179.810 2498.050 ;
        RECT 1178.150 2497.795 1178.430 2497.910 ;
        RECT 1179.530 2496.000 1179.810 2497.910 ;
        RECT 1255.890 436.715 1256.170 437.085 ;
        RECT 1255.960 436.405 1256.100 436.715 ;
        RECT 1255.890 436.035 1256.170 436.405 ;
        RECT 1956.470 436.035 1956.750 436.405 ;
        RECT 1993.730 436.035 1994.010 436.405 ;
        RECT 2124.830 436.035 2125.110 436.405 ;
        RECT 1895.290 435.355 1895.570 435.725 ;
        RECT 1895.300 435.210 1895.560 435.355 ;
        RECT 1930.260 435.215 1930.520 435.530 ;
        RECT 1930.250 434.845 1930.530 435.215 ;
        RECT 1956.540 435.190 1956.680 436.035 ;
        RECT 1993.800 435.610 1993.940 436.035 ;
        RECT 2124.900 435.870 2125.040 436.035 ;
        RECT 2090.340 435.725 2090.600 435.870 ;
        RECT 1994.650 435.610 1994.930 435.725 ;
        RECT 1993.800 435.470 1994.930 435.610 ;
        RECT 1994.650 435.355 1994.930 435.470 ;
        RECT 2090.330 435.355 2090.610 435.725 ;
        RECT 2124.840 435.550 2125.100 435.870 ;
        RECT 1932.100 435.045 1932.360 435.190 ;
        RECT 1932.090 434.675 1932.370 435.045 ;
        RECT 1956.480 434.870 1956.740 435.190 ;
        RECT 2042.030 434.675 2042.310 435.045 ;
        RECT 2069.630 434.675 2069.910 435.045 ;
        RECT 2042.040 434.530 2042.300 434.675 ;
        RECT 2069.640 434.530 2069.900 434.675 ;
      LAYER via2 ;
        RECT 1178.150 2497.840 1178.430 2498.120 ;
        RECT 1255.890 436.760 1256.170 437.040 ;
        RECT 1255.890 436.080 1256.170 436.360 ;
        RECT 1956.470 436.080 1956.750 436.360 ;
        RECT 1993.730 436.080 1994.010 436.360 ;
        RECT 2124.830 436.080 2125.110 436.360 ;
        RECT 1895.290 435.400 1895.570 435.680 ;
        RECT 1994.650 435.400 1994.930 435.680 ;
        RECT 2090.330 435.400 2090.610 435.680 ;
        RECT 1930.250 434.890 1930.530 435.170 ;
        RECT 1932.090 434.720 1932.370 435.000 ;
        RECT 2042.030 434.720 2042.310 435.000 ;
        RECT 2069.630 434.720 2069.910 435.000 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 439.020 2924.800 440.220 ;
=======
        RECT 1178.125 2498.140 1178.455 2498.145 ;
        RECT 1177.870 2498.130 1178.455 2498.140 ;
        RECT 1177.670 2497.830 1178.455 2498.130 ;
        RECT 1177.870 2497.820 1178.455 2497.830 ;
        RECT 1178.125 2497.815 1178.455 2497.820 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2916.710 439.470 2924.800 439.770 ;
        RECT 1177.870 437.050 1178.250 437.060 ;
        RECT 1255.865 437.050 1256.195 437.065 ;
        RECT 1177.870 436.750 1231.570 437.050 ;
        RECT 1177.870 436.740 1178.250 436.750 ;
        RECT 1231.270 436.370 1231.570 436.750 ;
        RECT 1255.865 436.750 1269.290 437.050 ;
        RECT 1255.865 436.735 1256.195 436.750 ;
        RECT 1255.865 436.370 1256.195 436.385 ;
        RECT 1231.270 436.070 1256.195 436.370 ;
        RECT 1268.990 436.370 1269.290 436.750 ;
        RECT 1738.150 436.370 1738.530 436.380 ;
        RECT 1834.750 436.370 1835.130 436.380 ;
        RECT 1268.990 436.070 1366.810 436.370 ;
        RECT 1255.865 436.055 1256.195 436.070 ;
        RECT 1366.510 435.690 1366.810 436.070 ;
        RECT 1463.110 436.070 1511.250 436.370 ;
        RECT 1463.110 435.690 1463.410 436.070 ;
        RECT 1366.510 435.390 1463.410 435.690 ;
        RECT 1510.950 435.010 1511.250 436.070 ;
        RECT 1617.670 436.070 1641.890 436.370 ;
        RECT 1617.670 435.690 1617.970 436.070 ;
        RECT 1559.710 435.390 1617.970 435.690 ;
        RECT 1559.710 435.010 1560.010 435.390 ;
        RECT 1510.950 434.710 1560.010 435.010 ;
        RECT 1641.590 435.010 1641.890 436.070 ;
        RECT 1703.230 436.070 1738.530 436.370 ;
        RECT 1703.230 435.690 1703.530 436.070 ;
        RECT 1738.150 436.060 1738.530 436.070 ;
        RECT 1799.830 436.070 1835.130 436.370 ;
        RECT 1799.830 435.690 1800.130 436.070 ;
        RECT 1834.750 436.060 1835.130 436.070 ;
        RECT 1956.445 436.370 1956.775 436.385 ;
        RECT 1993.705 436.370 1994.035 436.385 ;
        RECT 1956.445 436.070 1994.035 436.370 ;
        RECT 1956.445 436.055 1956.775 436.070 ;
        RECT 1993.705 436.055 1994.035 436.070 ;
        RECT 2124.805 436.370 2125.135 436.385 ;
        RECT 2124.805 436.070 2159.850 436.370 ;
        RECT 2124.805 436.055 2125.135 436.070 ;
        RECT 1895.265 435.690 1895.595 435.705 ;
        RECT 1656.310 435.390 1703.530 435.690 ;
        RECT 1752.910 435.390 1800.130 435.690 ;
        RECT 1849.510 435.390 1895.595 435.690 ;
        RECT 1656.310 435.010 1656.610 435.390 ;
        RECT 1641.590 434.710 1656.610 435.010 ;
        RECT 1738.150 435.010 1738.530 435.020 ;
        RECT 1752.910 435.010 1753.210 435.390 ;
        RECT 1738.150 434.710 1753.210 435.010 ;
        RECT 1834.750 435.010 1835.130 435.020 ;
        RECT 1849.510 435.010 1849.810 435.390 ;
        RECT 1895.265 435.375 1895.595 435.390 ;
        RECT 1994.625 435.690 1994.955 435.705 ;
        RECT 2090.305 435.690 2090.635 435.705 ;
        RECT 1994.625 435.390 2021.850 435.690 ;
        RECT 1994.625 435.375 1994.955 435.390 ;
        RECT 1834.750 434.710 1849.810 435.010 ;
        RECT 1930.225 435.180 1930.555 435.195 ;
        RECT 1930.225 435.010 1931.690 435.180 ;
        RECT 1932.065 435.010 1932.395 435.025 ;
        RECT 1930.225 434.880 1932.395 435.010 ;
        RECT 1930.225 434.865 1930.555 434.880 ;
        RECT 1931.390 434.710 1932.395 434.880 ;
        RECT 2021.550 435.010 2021.850 435.390 ;
        RECT 2076.750 435.390 2090.635 435.690 ;
        RECT 2159.550 435.690 2159.850 436.070 ;
        RECT 2208.310 436.070 2256.450 436.370 ;
        RECT 2159.550 435.390 2207.690 435.690 ;
        RECT 2042.005 435.010 2042.335 435.025 ;
        RECT 2021.550 434.710 2042.335 435.010 ;
        RECT 1738.150 434.700 1738.530 434.710 ;
        RECT 1834.750 434.700 1835.130 434.710 ;
        RECT 1932.065 434.695 1932.395 434.710 ;
        RECT 2042.005 434.695 2042.335 434.710 ;
        RECT 2069.605 435.010 2069.935 435.025 ;
        RECT 2076.750 435.010 2077.050 435.390 ;
        RECT 2090.305 435.375 2090.635 435.390 ;
        RECT 2069.605 434.710 2077.050 435.010 ;
        RECT 2207.390 435.010 2207.690 435.390 ;
        RECT 2208.310 435.010 2208.610 436.070 ;
        RECT 2256.150 435.690 2256.450 436.070 ;
        RECT 2304.910 436.070 2353.050 436.370 ;
        RECT 2256.150 435.390 2304.290 435.690 ;
        RECT 2207.390 434.710 2208.610 435.010 ;
        RECT 2303.990 435.010 2304.290 435.390 ;
        RECT 2304.910 435.010 2305.210 436.070 ;
        RECT 2352.750 435.690 2353.050 436.070 ;
        RECT 2401.510 436.070 2449.650 436.370 ;
        RECT 2352.750 435.390 2400.890 435.690 ;
        RECT 2303.990 434.710 2305.210 435.010 ;
        RECT 2400.590 435.010 2400.890 435.390 ;
        RECT 2401.510 435.010 2401.810 436.070 ;
        RECT 2449.350 435.690 2449.650 436.070 ;
        RECT 2498.110 436.070 2546.250 436.370 ;
        RECT 2449.350 435.390 2497.490 435.690 ;
        RECT 2400.590 434.710 2401.810 435.010 ;
        RECT 2497.190 435.010 2497.490 435.390 ;
        RECT 2498.110 435.010 2498.410 436.070 ;
        RECT 2545.950 435.690 2546.250 436.070 ;
        RECT 2594.710 436.070 2642.850 436.370 ;
        RECT 2545.950 435.390 2594.090 435.690 ;
        RECT 2497.190 434.710 2498.410 435.010 ;
        RECT 2593.790 435.010 2594.090 435.390 ;
        RECT 2594.710 435.010 2595.010 436.070 ;
        RECT 2642.550 435.690 2642.850 436.070 ;
        RECT 2691.310 436.070 2739.450 436.370 ;
        RECT 2642.550 435.390 2690.690 435.690 ;
        RECT 2593.790 434.710 2595.010 435.010 ;
        RECT 2690.390 435.010 2690.690 435.390 ;
        RECT 2691.310 435.010 2691.610 436.070 ;
        RECT 2739.150 435.690 2739.450 436.070 ;
        RECT 2787.910 436.070 2836.050 436.370 ;
        RECT 2739.150 435.390 2787.290 435.690 ;
        RECT 2690.390 434.710 2691.610 435.010 ;
        RECT 2786.990 435.010 2787.290 435.390 ;
        RECT 2787.910 435.010 2788.210 436.070 ;
        RECT 2835.750 435.690 2836.050 436.070 ;
        RECT 2916.710 435.690 2917.010 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
        RECT 2835.750 435.390 2883.890 435.690 ;
        RECT 2786.990 434.710 2788.210 435.010 ;
        RECT 2883.590 435.010 2883.890 435.390 ;
        RECT 2884.510 435.390 2917.010 435.690 ;
        RECT 2884.510 435.010 2884.810 435.390 ;
        RECT 2883.590 434.710 2884.810 435.010 ;
        RECT 2069.605 434.695 2069.935 434.710 ;
      LAYER via3 ;
        RECT 1177.900 2497.820 1178.220 2498.140 ;
        RECT 1177.900 436.740 1178.220 437.060 ;
        RECT 1738.180 436.060 1738.500 436.380 ;
        RECT 1834.780 436.060 1835.100 436.380 ;
        RECT 1738.180 434.700 1738.500 435.020 ;
        RECT 1834.780 434.700 1835.100 435.020 ;
      LAYER met4 ;
        RECT 1177.895 2497.815 1178.225 2498.145 ;
        RECT 1177.910 437.065 1178.210 2497.815 ;
        RECT 1177.895 436.735 1178.225 437.065 ;
        RECT 1738.175 436.055 1738.505 436.385 ;
        RECT 1834.775 436.055 1835.105 436.385 ;
        RECT 1738.190 435.025 1738.490 436.055 ;
        RECT 1834.790 435.025 1835.090 436.055 ;
        RECT 1738.175 434.695 1738.505 435.025 ;
        RECT 1834.775 434.695 1835.105 435.025 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3501.220 1014.230 3501.280 ;
        RECT 1535.090 3501.220 1535.410 3501.280 ;
        RECT 1013.910 3501.080 1535.410 3501.220 ;
        RECT 1013.910 3501.020 1014.230 3501.080 ;
        RECT 1535.090 3501.020 1535.410 3501.080 ;
        RECT 1535.090 2518.280 1535.410 2518.340 ;
        RECT 1554.870 2518.280 1555.190 2518.340 ;
        RECT 1535.090 2518.140 1555.190 2518.280 ;
        RECT 1535.090 2518.080 1535.410 2518.140 ;
        RECT 1554.870 2518.080 1555.190 2518.140 ;
      LAYER via ;
        RECT 1013.940 3501.020 1014.200 3501.280 ;
        RECT 1535.120 3501.020 1535.380 3501.280 ;
        RECT 1535.120 2518.080 1535.380 2518.340 ;
        RECT 1554.900 2518.080 1555.160 2518.340 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1013.790 3519.700 1014.350 3524.800 ;
=======
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3501.310 1014.140 3517.600 ;
        RECT 1013.940 3500.990 1014.200 3501.310 ;
        RECT 1535.120 3500.990 1535.380 3501.310 ;
        RECT 1535.180 2518.370 1535.320 3500.990 ;
        RECT 1535.120 2518.050 1535.380 2518.370 ;
        RECT 1554.900 2518.050 1555.160 2518.370 ;
        RECT 1554.960 2499.410 1555.100 2518.050 ;
        RECT 1556.270 2499.410 1556.550 2500.000 ;
        RECT 1554.960 2499.270 1556.550 2499.410 ;
        RECT 1556.270 2496.000 1556.550 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 689.150 3503.940 689.470 3504.000 ;
        RECT 1555.790 3503.940 1556.110 3504.000 ;
        RECT 689.150 3503.800 1556.110 3503.940 ;
        RECT 689.150 3503.740 689.470 3503.800 ;
        RECT 1555.790 3503.740 1556.110 3503.800 ;
        RECT 1562.320 2518.480 1563.840 2518.620 ;
        RECT 1555.790 2518.280 1556.110 2518.340 ;
        RECT 1562.320 2518.280 1562.460 2518.480 ;
        RECT 1555.790 2518.140 1562.460 2518.280 ;
        RECT 1555.790 2518.080 1556.110 2518.140 ;
        RECT 1563.700 2517.940 1563.840 2518.480 ;
        RECT 1576.030 2517.940 1576.350 2518.000 ;
        RECT 1563.700 2517.800 1576.350 2517.940 ;
        RECT 1576.030 2517.740 1576.350 2517.800 ;
      LAYER via ;
        RECT 689.180 3503.740 689.440 3504.000 ;
        RECT 1555.820 3503.740 1556.080 3504.000 ;
        RECT 1555.820 2518.080 1556.080 2518.340 ;
        RECT 1576.060 2517.740 1576.320 2518.000 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 689.030 3519.700 689.590 3524.800 ;
=======
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3504.030 689.380 3517.600 ;
        RECT 689.180 3503.710 689.440 3504.030 ;
        RECT 1555.820 3503.710 1556.080 3504.030 ;
        RECT 1555.880 2518.370 1556.020 3503.710 ;
        RECT 1555.820 2518.050 1556.080 2518.370 ;
        RECT 1576.060 2517.710 1576.320 2518.030 ;
        RECT 1576.120 2500.000 1576.260 2517.710 ;
        RECT 1576.050 2496.000 1576.330 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.240 365.170 3502.300 ;
        RECT 1576.490 3502.240 1576.810 3502.300 ;
        RECT 364.850 3502.100 1576.810 3502.240 ;
        RECT 364.850 3502.040 365.170 3502.100 ;
        RECT 1576.490 3502.040 1576.810 3502.100 ;
        RECT 1576.490 2517.940 1576.810 2518.000 ;
        RECT 1595.810 2517.940 1596.130 2518.000 ;
        RECT 1576.490 2517.800 1596.130 2517.940 ;
        RECT 1576.490 2517.740 1576.810 2517.800 ;
        RECT 1595.810 2517.740 1596.130 2517.800 ;
      LAYER via ;
        RECT 364.880 3502.040 365.140 3502.300 ;
        RECT 1576.520 3502.040 1576.780 3502.300 ;
        RECT 1576.520 2517.740 1576.780 2518.000 ;
        RECT 1595.840 2517.740 1596.100 2518.000 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 364.730 3519.700 365.290 3524.800 ;
=======
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3502.330 365.080 3517.600 ;
        RECT 364.880 3502.010 365.140 3502.330 ;
        RECT 1576.520 3502.010 1576.780 3502.330 ;
        RECT 1576.580 2518.030 1576.720 3502.010 ;
        RECT 1576.520 2517.710 1576.780 2518.030 ;
        RECT 1595.840 2517.710 1596.100 2518.030 ;
        RECT 1595.900 2500.000 1596.040 2517.710 ;
        RECT 1595.830 2496.000 1596.110 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1597.190 2517.940 1597.510 2518.000 ;
        RECT 1616.050 2517.940 1616.370 2518.000 ;
        RECT 1597.190 2517.800 1616.370 2517.940 ;
        RECT 1597.190 2517.740 1597.510 2517.800 ;
        RECT 1616.050 2517.740 1616.370 2517.800 ;
      LAYER via ;
        RECT 1597.220 2517.740 1597.480 2518.000 ;
        RECT 1616.080 2517.740 1616.340 2518.000 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 40.430 3519.700 40.990 3524.800 ;
=======
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
        RECT 1597.210 3501.475 1597.490 3501.845 ;
        RECT 1597.280 2518.030 1597.420 3501.475 ;
        RECT 1597.220 2517.710 1597.480 2518.030 ;
        RECT 1616.080 2517.710 1616.340 2518.030 ;
        RECT 1616.140 2500.000 1616.280 2517.710 ;
        RECT 1616.070 2496.000 1616.350 2500.000 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
        RECT 1597.210 3501.520 1597.490 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 1597.185 3501.810 1597.515 3501.825 ;
        RECT 40.545 3501.510 1597.515 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
        RECT 1597.185 3501.495 1597.515 3501.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 1635.370 3263.900 1635.690 3263.960 ;
        RECT 15.250 3263.760 1635.690 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 1635.370 3263.700 1635.690 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 1635.400 3263.700 1635.660 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 1635.400 3263.670 1635.660 3263.990 ;
        RECT 1635.460 2499.410 1635.600 3263.670 ;
        RECT 1635.850 2499.410 1636.130 2500.000 ;
        RECT 1635.460 2499.270 1636.130 2499.410 ;
        RECT 1635.850 2496.000 1636.130 2499.270 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3267.140 0.300 3268.340 ;
=======
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 2974.220 16.490 2974.280 ;
        RECT 1649.170 2974.220 1649.490 2974.280 ;
        RECT 16.170 2974.080 1649.490 2974.220 ;
        RECT 16.170 2974.020 16.490 2974.080 ;
        RECT 1649.170 2974.020 1649.490 2974.080 ;
      LAYER via ;
        RECT 16.200 2974.020 16.460 2974.280 ;
        RECT 1649.200 2974.020 1649.460 2974.280 ;
      LAYER met2 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 16.260 2974.310 16.400 2979.915 ;
        RECT 16.200 2973.990 16.460 2974.310 ;
        RECT 1649.200 2973.990 1649.460 2974.310 ;
        RECT 1649.260 2500.090 1649.400 2973.990 ;
        RECT 1649.260 2499.950 1653.080 2500.090 ;
        RECT 1652.940 2499.410 1653.080 2499.950 ;
        RECT 1655.630 2499.410 1655.910 2500.000 ;
        RECT 1652.940 2499.270 1655.910 2499.410 ;
        RECT 1655.630 2496.000 1655.910 2499.270 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2979.500 0.300 2980.700 ;
=======
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.800 2979.950 16.495 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2691.340 17.410 2691.400 ;
        RECT 1669.870 2691.340 1670.190 2691.400 ;
        RECT 17.090 2691.200 1670.190 2691.340 ;
        RECT 17.090 2691.140 17.410 2691.200 ;
        RECT 1669.870 2691.140 1670.190 2691.200 ;
      LAYER via ;
        RECT 17.120 2691.140 17.380 2691.400 ;
        RECT 1669.900 2691.140 1670.160 2691.400 ;
      LAYER met2 ;
        RECT 17.110 2692.955 17.390 2693.325 ;
        RECT 17.180 2691.430 17.320 2692.955 ;
        RECT 17.120 2691.110 17.380 2691.430 ;
        RECT 1669.900 2691.110 1670.160 2691.430 ;
        RECT 1669.960 2500.090 1670.100 2691.110 ;
        RECT 1669.960 2499.950 1672.400 2500.090 ;
        RECT 1672.260 2499.410 1672.400 2499.950 ;
        RECT 1675.410 2499.410 1675.690 2500.000 ;
        RECT 1672.260 2499.270 1675.690 2499.410 ;
        RECT 1675.410 2496.000 1675.690 2499.270 ;
      LAYER via2 ;
        RECT 17.110 2693.000 17.390 2693.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2692.540 0.300 2693.740 ;
=======
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 17.085 2693.290 17.415 2693.305 ;
        RECT -4.800 2692.990 17.415 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 17.085 2692.975 17.415 2692.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 22.150 2513.520 22.470 2513.580 ;
        RECT 1695.170 2513.520 1695.490 2513.580 ;
        RECT 22.150 2513.380 1695.490 2513.520 ;
        RECT 22.150 2513.320 22.470 2513.380 ;
        RECT 1695.170 2513.320 1695.490 2513.380 ;
        RECT 13.870 2405.740 14.190 2405.800 ;
        RECT 22.150 2405.740 22.470 2405.800 ;
        RECT 13.870 2405.600 22.470 2405.740 ;
        RECT 13.870 2405.540 14.190 2405.600 ;
        RECT 22.150 2405.540 22.470 2405.600 ;
      LAYER via ;
        RECT 22.180 2513.320 22.440 2513.580 ;
        RECT 1695.200 2513.320 1695.460 2513.580 ;
        RECT 13.900 2405.540 14.160 2405.800 ;
        RECT 22.180 2405.540 22.440 2405.800 ;
      LAYER met2 ;
        RECT 22.180 2513.290 22.440 2513.610 ;
        RECT 1695.200 2513.290 1695.460 2513.610 ;
        RECT 22.240 2405.830 22.380 2513.290 ;
        RECT 1695.260 2500.000 1695.400 2513.290 ;
        RECT 1695.190 2496.000 1695.470 2500.000 ;
        RECT 13.900 2405.685 14.160 2405.830 ;
        RECT 13.890 2405.315 14.170 2405.685 ;
        RECT 22.180 2405.510 22.440 2405.830 ;
      LAYER via2 ;
        RECT 13.890 2405.360 14.170 2405.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2404.900 0.300 2406.100 ;
=======
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 13.865 2405.650 14.195 2405.665 ;
        RECT -4.800 2405.350 14.195 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 13.865 2405.335 14.195 2405.350 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23.070 2512.840 23.390 2512.900 ;
        RECT 1714.950 2512.840 1715.270 2512.900 ;
        RECT 23.070 2512.700 1715.270 2512.840 ;
        RECT 23.070 2512.640 23.390 2512.700 ;
        RECT 1714.950 2512.640 1715.270 2512.700 ;
        RECT 13.870 2118.780 14.190 2118.840 ;
        RECT 23.070 2118.780 23.390 2118.840 ;
        RECT 13.870 2118.640 23.390 2118.780 ;
        RECT 13.870 2118.580 14.190 2118.640 ;
        RECT 23.070 2118.580 23.390 2118.640 ;
      LAYER via ;
        RECT 23.100 2512.640 23.360 2512.900 ;
        RECT 1714.980 2512.640 1715.240 2512.900 ;
        RECT 13.900 2118.580 14.160 2118.840 ;
        RECT 23.100 2118.580 23.360 2118.840 ;
      LAYER met2 ;
        RECT 23.100 2512.610 23.360 2512.930 ;
        RECT 1714.980 2512.610 1715.240 2512.930 ;
        RECT 23.160 2118.870 23.300 2512.610 ;
        RECT 1715.040 2500.000 1715.180 2512.610 ;
        RECT 1714.970 2496.000 1715.250 2500.000 ;
        RECT 13.900 2118.725 14.160 2118.870 ;
        RECT 13.890 2118.355 14.170 2118.725 ;
        RECT 23.100 2118.550 23.360 2118.870 ;
      LAYER via2 ;
        RECT 13.890 2118.400 14.170 2118.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2117.940 0.300 2119.140 ;
=======
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 13.865 2118.690 14.195 2118.705 ;
        RECT -4.800 2118.390 14.195 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 13.865 2118.375 14.195 2118.390 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2512.160 16.030 2512.220 ;
        RECT 1734.730 2512.160 1735.050 2512.220 ;
        RECT 15.710 2512.020 1735.050 2512.160 ;
        RECT 15.710 2511.960 16.030 2512.020 ;
        RECT 1734.730 2511.960 1735.050 2512.020 ;
      LAYER via ;
        RECT 15.740 2511.960 16.000 2512.220 ;
        RECT 1734.760 2511.960 1735.020 2512.220 ;
      LAYER met2 ;
        RECT 15.740 2511.930 16.000 2512.250 ;
        RECT 1734.760 2511.930 1735.020 2512.250 ;
        RECT 15.800 1831.085 15.940 2511.930 ;
        RECT 1734.820 2500.000 1734.960 2511.930 ;
        RECT 1734.750 2496.000 1735.030 2500.000 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1830.300 0.300 1831.500 ;
=======
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1200.670 670.720 1200.990 670.780 ;
        RECT 1231.490 670.720 1231.810 670.780 ;
        RECT 1200.670 670.580 1231.810 670.720 ;
        RECT 1200.670 670.520 1200.990 670.580 ;
        RECT 1231.490 670.520 1231.810 670.580 ;
        RECT 1490.470 670.720 1490.790 670.780 ;
        RECT 1514.850 670.720 1515.170 670.780 ;
        RECT 1490.470 670.580 1515.170 670.720 ;
        RECT 1490.470 670.520 1490.790 670.580 ;
        RECT 1514.850 670.520 1515.170 670.580 ;
        RECT 1352.010 670.380 1352.330 670.440 ;
        RECT 1355.230 670.380 1355.550 670.440 ;
        RECT 1352.010 670.240 1355.550 670.380 ;
        RECT 1352.010 670.180 1352.330 670.240 ;
        RECT 1355.230 670.180 1355.550 670.240 ;
        RECT 1400.770 670.380 1401.090 670.440 ;
        RECT 1403.070 670.380 1403.390 670.440 ;
        RECT 1400.770 670.240 1403.390 670.380 ;
        RECT 1400.770 670.180 1401.090 670.240 ;
        RECT 1403.070 670.180 1403.390 670.240 ;
        RECT 1798.670 670.380 1798.990 670.440 ;
        RECT 1811.550 670.380 1811.870 670.440 ;
        RECT 1798.670 670.240 1811.870 670.380 ;
        RECT 1798.670 670.180 1798.990 670.240 ;
        RECT 1811.550 670.180 1811.870 670.240 ;
        RECT 2090.310 670.380 2090.630 670.440 ;
        RECT 2124.810 670.380 2125.130 670.440 ;
        RECT 2090.310 670.240 2125.130 670.380 ;
        RECT 2090.310 670.180 2090.630 670.240 ;
        RECT 2124.810 670.180 2125.130 670.240 ;
        RECT 1606.390 670.040 1606.710 670.100 ;
        RECT 1607.770 670.040 1608.090 670.100 ;
        RECT 1606.390 669.900 1608.090 670.040 ;
        RECT 1606.390 669.840 1606.710 669.900 ;
        RECT 1607.770 669.840 1608.090 669.900 ;
        RECT 1702.070 670.040 1702.390 670.100 ;
        RECT 1714.490 670.040 1714.810 670.100 ;
        RECT 1702.070 669.900 1714.810 670.040 ;
        RECT 1702.070 669.840 1702.390 669.900 ;
        RECT 1714.490 669.840 1714.810 669.900 ;
        RECT 1544.750 669.700 1545.070 669.760 ;
        RECT 1561.310 669.700 1561.630 669.760 ;
        RECT 1544.750 669.560 1561.630 669.700 ;
        RECT 1544.750 669.500 1545.070 669.560 ;
        RECT 1561.310 669.500 1561.630 669.560 ;
        RECT 1932.070 669.700 1932.390 669.760 ;
        RECT 1946.330 669.700 1946.650 669.760 ;
        RECT 1932.070 669.560 1946.650 669.700 ;
        RECT 1932.070 669.500 1932.390 669.560 ;
        RECT 1946.330 669.500 1946.650 669.560 ;
      LAYER via ;
        RECT 1200.700 670.520 1200.960 670.780 ;
        RECT 1231.520 670.520 1231.780 670.780 ;
        RECT 1490.500 670.520 1490.760 670.780 ;
        RECT 1514.880 670.520 1515.140 670.780 ;
        RECT 1352.040 670.180 1352.300 670.440 ;
        RECT 1355.260 670.180 1355.520 670.440 ;
        RECT 1400.800 670.180 1401.060 670.440 ;
        RECT 1403.100 670.180 1403.360 670.440 ;
        RECT 1798.700 670.180 1798.960 670.440 ;
        RECT 1811.580 670.180 1811.840 670.440 ;
        RECT 2090.340 670.180 2090.600 670.440 ;
        RECT 2124.840 670.180 2125.100 670.440 ;
        RECT 1606.420 669.840 1606.680 670.100 ;
        RECT 1607.800 669.840 1608.060 670.100 ;
        RECT 1702.100 669.840 1702.360 670.100 ;
        RECT 1714.520 669.840 1714.780 670.100 ;
        RECT 1544.780 669.500 1545.040 669.760 ;
        RECT 1561.340 669.500 1561.600 669.760 ;
        RECT 1932.100 669.500 1932.360 669.760 ;
        RECT 1946.360 669.500 1946.620 669.760 ;
      LAYER met2 ;
        RECT 1199.310 2498.050 1199.590 2500.000 ;
        RECT 1199.770 2498.050 1200.050 2498.165 ;
        RECT 1199.310 2497.910 1200.050 2498.050 ;
        RECT 1199.310 2496.000 1199.590 2497.910 ;
        RECT 1199.770 2497.795 1200.050 2497.910 ;
        RECT 2028.230 671.995 2028.510 672.365 ;
        RECT 1200.690 670.635 1200.970 671.005 ;
        RECT 1200.700 670.490 1200.960 670.635 ;
        RECT 1231.520 670.490 1231.780 670.810 ;
        RECT 1266.010 670.635 1266.290 671.005 ;
        RECT 1403.090 670.635 1403.370 671.005 ;
        RECT 1490.490 670.635 1490.770 671.005 ;
        RECT 1231.580 670.325 1231.720 670.490 ;
        RECT 1231.510 669.955 1231.790 670.325 ;
        RECT 1266.080 669.645 1266.220 670.635 ;
        RECT 1403.160 670.470 1403.300 670.635 ;
        RECT 1490.500 670.490 1490.760 670.635 ;
        RECT 1514.880 670.490 1515.140 670.810 ;
        RECT 1561.330 670.635 1561.610 671.005 ;
        RECT 1946.350 670.635 1946.630 671.005 ;
        RECT 1352.040 670.325 1352.300 670.470 ;
        RECT 1355.260 670.325 1355.520 670.470 ;
        RECT 1400.800 670.325 1401.060 670.470 ;
        RECT 1352.030 669.955 1352.310 670.325 ;
        RECT 1355.250 669.955 1355.530 670.325 ;
        RECT 1400.790 669.955 1401.070 670.325 ;
        RECT 1403.100 670.150 1403.360 670.470 ;
        RECT 1514.940 669.645 1515.080 670.490 ;
        RECT 1561.400 669.790 1561.540 670.635 ;
        RECT 1798.700 670.325 1798.960 670.470 ;
        RECT 1811.580 670.325 1811.840 670.470 ;
        RECT 1606.410 669.955 1606.690 670.325 ;
        RECT 1607.790 669.955 1608.070 670.325 ;
        RECT 1702.090 669.955 1702.370 670.325 ;
        RECT 1714.510 669.955 1714.790 670.325 ;
        RECT 1798.690 669.955 1798.970 670.325 ;
        RECT 1811.570 669.955 1811.850 670.325 ;
        RECT 1895.290 669.955 1895.570 670.325 ;
        RECT 1606.420 669.810 1606.680 669.955 ;
        RECT 1607.800 669.810 1608.060 669.955 ;
        RECT 1702.100 669.810 1702.360 669.955 ;
        RECT 1714.520 669.810 1714.780 669.955 ;
        RECT 1544.780 669.645 1545.040 669.790 ;
        RECT 1266.010 669.275 1266.290 669.645 ;
        RECT 1514.870 669.275 1515.150 669.645 ;
        RECT 1544.770 669.275 1545.050 669.645 ;
        RECT 1561.340 669.470 1561.600 669.790 ;
        RECT 1895.360 668.285 1895.500 669.955 ;
        RECT 1946.420 669.790 1946.560 670.635 ;
        RECT 2028.300 670.325 2028.440 671.995 ;
        RECT 2052.610 671.315 2052.890 671.685 ;
        RECT 2028.230 669.955 2028.510 670.325 ;
        RECT 1932.100 669.645 1932.360 669.790 ;
        RECT 1932.090 669.275 1932.370 669.645 ;
        RECT 1946.360 669.470 1946.620 669.790 ;
        RECT 2052.680 669.645 2052.820 671.315 ;
        RECT 2124.830 670.635 2125.110 671.005 ;
        RECT 2124.900 670.470 2125.040 670.635 ;
        RECT 2090.340 670.325 2090.600 670.470 ;
        RECT 2090.330 669.955 2090.610 670.325 ;
        RECT 2124.840 670.150 2125.100 670.470 ;
        RECT 2052.610 669.275 2052.890 669.645 ;
        RECT 1895.290 667.915 1895.570 668.285 ;
      LAYER via2 ;
        RECT 1199.770 2497.840 1200.050 2498.120 ;
        RECT 2028.230 672.040 2028.510 672.320 ;
        RECT 1200.690 670.680 1200.970 670.960 ;
        RECT 1266.010 670.680 1266.290 670.960 ;
        RECT 1403.090 670.680 1403.370 670.960 ;
        RECT 1490.490 670.680 1490.770 670.960 ;
        RECT 1231.510 670.000 1231.790 670.280 ;
        RECT 1561.330 670.680 1561.610 670.960 ;
        RECT 1946.350 670.680 1946.630 670.960 ;
        RECT 1352.030 670.000 1352.310 670.280 ;
        RECT 1355.250 670.000 1355.530 670.280 ;
        RECT 1400.790 670.000 1401.070 670.280 ;
        RECT 1606.410 670.000 1606.690 670.280 ;
        RECT 1607.790 670.000 1608.070 670.280 ;
        RECT 1702.090 670.000 1702.370 670.280 ;
        RECT 1714.510 670.000 1714.790 670.280 ;
        RECT 1798.690 670.000 1798.970 670.280 ;
        RECT 1811.570 670.000 1811.850 670.280 ;
        RECT 1895.290 670.000 1895.570 670.280 ;
        RECT 1266.010 669.320 1266.290 669.600 ;
        RECT 1514.870 669.320 1515.150 669.600 ;
        RECT 1544.770 669.320 1545.050 669.600 ;
        RECT 2052.610 671.360 2052.890 671.640 ;
        RECT 2028.230 670.000 2028.510 670.280 ;
        RECT 1932.090 669.320 1932.370 669.600 ;
        RECT 2124.830 670.680 2125.110 670.960 ;
        RECT 2090.330 670.000 2090.610 670.280 ;
        RECT 2052.610 669.320 2052.890 669.600 ;
        RECT 1895.290 667.960 1895.570 668.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 673.620 2924.800 674.820 ;
=======
        RECT 1199.745 2498.140 1200.075 2498.145 ;
        RECT 1199.745 2498.130 1200.330 2498.140 ;
        RECT 1199.745 2497.830 1200.530 2498.130 ;
        RECT 1199.745 2497.820 1200.330 2497.830 ;
        RECT 1199.745 2497.815 1200.075 2497.820 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2916.710 674.070 2924.800 674.370 ;
        RECT 1980.110 672.330 1980.490 672.340 ;
        RECT 2028.205 672.330 2028.535 672.345 ;
        RECT 1980.110 672.030 2028.535 672.330 ;
        RECT 1980.110 672.020 1980.490 672.030 ;
        RECT 2028.205 672.015 2028.535 672.030 ;
        RECT 2052.585 671.650 2052.915 671.665 ;
        RECT 2028.910 671.350 2052.915 671.650 ;
        RECT 1199.950 670.970 1200.330 670.980 ;
        RECT 1200.665 670.970 1200.995 670.985 ;
        RECT 1199.950 670.670 1200.995 670.970 ;
        RECT 1199.950 670.660 1200.330 670.670 ;
        RECT 1200.665 670.655 1200.995 670.670 ;
        RECT 1265.985 670.970 1266.315 670.985 ;
        RECT 1403.065 670.970 1403.395 670.985 ;
        RECT 1490.465 670.970 1490.795 670.985 ;
        RECT 1265.985 670.800 1290.450 670.970 ;
        RECT 1265.985 670.670 1291.370 670.800 ;
        RECT 1265.985 670.655 1266.315 670.670 ;
        RECT 1290.150 670.500 1291.370 670.670 ;
        RECT 1403.065 670.670 1490.795 670.970 ;
        RECT 1403.065 670.655 1403.395 670.670 ;
        RECT 1490.465 670.655 1490.795 670.670 ;
        RECT 1561.305 670.970 1561.635 670.985 ;
        RECT 1946.325 670.970 1946.655 670.985 ;
        RECT 1980.110 670.970 1980.490 670.980 ;
        RECT 1561.305 670.670 1586.690 670.970 ;
        RECT 1561.305 670.655 1561.635 670.670 ;
        RECT 1231.485 670.290 1231.815 670.305 ;
        RECT 1291.070 670.290 1291.370 670.500 ;
        RECT 1352.005 670.290 1352.335 670.305 ;
        RECT 1231.485 669.990 1248.130 670.290 ;
        RECT 1291.070 669.990 1352.335 670.290 ;
        RECT 1231.485 669.975 1231.815 669.990 ;
        RECT 1247.830 669.610 1248.130 669.990 ;
        RECT 1352.005 669.975 1352.335 669.990 ;
        RECT 1355.225 670.290 1355.555 670.305 ;
        RECT 1400.765 670.290 1401.095 670.305 ;
        RECT 1355.225 669.990 1401.095 670.290 ;
        RECT 1586.390 670.290 1586.690 670.670 ;
        RECT 1946.325 670.670 1980.490 670.970 ;
        RECT 1946.325 670.655 1946.655 670.670 ;
        RECT 1980.110 670.660 1980.490 670.670 ;
        RECT 1606.385 670.290 1606.715 670.305 ;
        RECT 1586.390 669.990 1606.715 670.290 ;
        RECT 1355.225 669.975 1355.555 669.990 ;
        RECT 1400.765 669.975 1401.095 669.990 ;
        RECT 1606.385 669.975 1606.715 669.990 ;
        RECT 1607.765 670.290 1608.095 670.305 ;
        RECT 1702.065 670.290 1702.395 670.305 ;
        RECT 1607.765 669.990 1641.890 670.290 ;
        RECT 1607.765 669.975 1608.095 669.990 ;
        RECT 1265.985 669.610 1266.315 669.625 ;
        RECT 1247.830 669.310 1266.315 669.610 ;
        RECT 1265.985 669.295 1266.315 669.310 ;
        RECT 1514.845 669.610 1515.175 669.625 ;
        RECT 1544.745 669.610 1545.075 669.625 ;
        RECT 1514.845 669.310 1545.075 669.610 ;
        RECT 1641.590 669.610 1641.890 669.990 ;
        RECT 1656.310 669.990 1702.395 670.290 ;
        RECT 1656.310 669.610 1656.610 669.990 ;
        RECT 1702.065 669.975 1702.395 669.990 ;
        RECT 1714.485 670.290 1714.815 670.305 ;
        RECT 1798.665 670.290 1798.995 670.305 ;
        RECT 1714.485 669.990 1738.490 670.290 ;
        RECT 1714.485 669.975 1714.815 669.990 ;
        RECT 1641.590 669.310 1656.610 669.610 ;
        RECT 1738.190 669.610 1738.490 669.990 ;
        RECT 1752.910 669.990 1798.995 670.290 ;
        RECT 1752.910 669.610 1753.210 669.990 ;
        RECT 1798.665 669.975 1798.995 669.990 ;
        RECT 1811.545 670.290 1811.875 670.305 ;
        RECT 1895.265 670.290 1895.595 670.305 ;
        RECT 1811.545 669.990 1835.090 670.290 ;
        RECT 1811.545 669.975 1811.875 669.990 ;
        RECT 1738.190 669.310 1753.210 669.610 ;
        RECT 1834.790 669.610 1835.090 669.990 ;
        RECT 1849.510 669.990 1895.595 670.290 ;
        RECT 1849.510 669.610 1849.810 669.990 ;
        RECT 1895.265 669.975 1895.595 669.990 ;
        RECT 2028.205 670.290 2028.535 670.305 ;
        RECT 2028.910 670.290 2029.210 671.350 ;
        RECT 2052.585 671.335 2052.915 671.350 ;
        RECT 2124.805 670.970 2125.135 670.985 ;
        RECT 2124.805 670.670 2159.850 670.970 ;
        RECT 2124.805 670.655 2125.135 670.670 ;
        RECT 2090.305 670.290 2090.635 670.305 ;
        RECT 2028.205 669.990 2029.210 670.290 ;
        RECT 2076.750 669.990 2090.635 670.290 ;
        RECT 2159.550 670.290 2159.850 670.670 ;
        RECT 2208.310 670.670 2256.450 670.970 ;
        RECT 2159.550 669.990 2207.690 670.290 ;
        RECT 2028.205 669.975 2028.535 669.990 ;
        RECT 1932.065 669.610 1932.395 669.625 ;
        RECT 1834.790 669.310 1849.810 669.610 ;
        RECT 1931.390 669.310 1932.395 669.610 ;
        RECT 1514.845 669.295 1515.175 669.310 ;
        RECT 1544.745 669.295 1545.075 669.310 ;
        RECT 1895.265 668.250 1895.595 668.265 ;
        RECT 1931.390 668.250 1931.690 669.310 ;
        RECT 1932.065 669.295 1932.395 669.310 ;
        RECT 2052.585 669.610 2052.915 669.625 ;
        RECT 2076.750 669.610 2077.050 669.990 ;
        RECT 2090.305 669.975 2090.635 669.990 ;
        RECT 2052.585 669.310 2077.050 669.610 ;
        RECT 2207.390 669.610 2207.690 669.990 ;
        RECT 2208.310 669.610 2208.610 670.670 ;
        RECT 2256.150 670.290 2256.450 670.670 ;
        RECT 2304.910 670.670 2353.050 670.970 ;
        RECT 2256.150 669.990 2304.290 670.290 ;
        RECT 2207.390 669.310 2208.610 669.610 ;
        RECT 2303.990 669.610 2304.290 669.990 ;
        RECT 2304.910 669.610 2305.210 670.670 ;
        RECT 2352.750 670.290 2353.050 670.670 ;
        RECT 2401.510 670.670 2449.650 670.970 ;
        RECT 2352.750 669.990 2400.890 670.290 ;
        RECT 2303.990 669.310 2305.210 669.610 ;
        RECT 2400.590 669.610 2400.890 669.990 ;
        RECT 2401.510 669.610 2401.810 670.670 ;
        RECT 2449.350 670.290 2449.650 670.670 ;
        RECT 2498.110 670.670 2546.250 670.970 ;
        RECT 2449.350 669.990 2497.490 670.290 ;
        RECT 2400.590 669.310 2401.810 669.610 ;
        RECT 2497.190 669.610 2497.490 669.990 ;
        RECT 2498.110 669.610 2498.410 670.670 ;
        RECT 2545.950 670.290 2546.250 670.670 ;
        RECT 2594.710 670.670 2642.850 670.970 ;
        RECT 2545.950 669.990 2594.090 670.290 ;
        RECT 2497.190 669.310 2498.410 669.610 ;
        RECT 2593.790 669.610 2594.090 669.990 ;
        RECT 2594.710 669.610 2595.010 670.670 ;
        RECT 2642.550 670.290 2642.850 670.670 ;
        RECT 2691.310 670.670 2739.450 670.970 ;
        RECT 2642.550 669.990 2690.690 670.290 ;
        RECT 2593.790 669.310 2595.010 669.610 ;
        RECT 2690.390 669.610 2690.690 669.990 ;
        RECT 2691.310 669.610 2691.610 670.670 ;
        RECT 2739.150 670.290 2739.450 670.670 ;
        RECT 2787.910 670.670 2836.050 670.970 ;
        RECT 2739.150 669.990 2787.290 670.290 ;
        RECT 2690.390 669.310 2691.610 669.610 ;
        RECT 2786.990 669.610 2787.290 669.990 ;
        RECT 2787.910 669.610 2788.210 670.670 ;
        RECT 2835.750 670.290 2836.050 670.670 ;
        RECT 2916.710 670.290 2917.010 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
        RECT 2835.750 669.990 2883.890 670.290 ;
        RECT 2786.990 669.310 2788.210 669.610 ;
        RECT 2883.590 669.610 2883.890 669.990 ;
        RECT 2884.510 669.990 2917.010 670.290 ;
        RECT 2884.510 669.610 2884.810 669.990 ;
        RECT 2883.590 669.310 2884.810 669.610 ;
        RECT 2052.585 669.295 2052.915 669.310 ;
        RECT 1895.265 667.950 1931.690 668.250 ;
        RECT 1895.265 667.935 1895.595 667.950 ;
      LAYER via3 ;
        RECT 1199.980 2497.820 1200.300 2498.140 ;
        RECT 1980.140 672.020 1980.460 672.340 ;
        RECT 1199.980 670.660 1200.300 670.980 ;
        RECT 1980.140 670.660 1980.460 670.980 ;
      LAYER met4 ;
        RECT 1199.975 2497.815 1200.305 2498.145 ;
        RECT 1199.990 670.985 1200.290 2497.815 ;
        RECT 1980.135 672.015 1980.465 672.345 ;
        RECT 1980.150 670.985 1980.450 672.015 ;
        RECT 1199.975 670.655 1200.305 670.985 ;
        RECT 1980.135 670.655 1980.465 670.985 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1752.745 2494.325 1752.915 2496.875 ;
      LAYER mcon ;
        RECT 1752.745 2496.705 1752.915 2496.875 ;
      LAYER met1 ;
        RECT 1752.670 2496.860 1752.990 2496.920 ;
        RECT 1752.475 2496.720 1752.990 2496.860 ;
        RECT 1752.670 2496.660 1752.990 2496.720 ;
        RECT 16.630 2494.480 16.950 2494.540 ;
        RECT 1752.685 2494.480 1752.975 2494.525 ;
        RECT 16.630 2494.340 1752.975 2494.480 ;
        RECT 16.630 2494.280 16.950 2494.340 ;
        RECT 1752.685 2494.295 1752.975 2494.340 ;
      LAYER via ;
        RECT 1752.700 2496.660 1752.960 2496.920 ;
        RECT 16.660 2494.280 16.920 2494.540 ;
      LAYER met2 ;
        RECT 1752.700 2496.690 1752.960 2496.950 ;
        RECT 1754.530 2496.690 1754.810 2500.000 ;
        RECT 1752.700 2496.630 1754.810 2496.690 ;
        RECT 1752.760 2496.550 1754.810 2496.630 ;
        RECT 1754.530 2496.000 1754.810 2496.550 ;
        RECT 16.660 2494.250 16.920 2494.570 ;
        RECT 16.720 1544.125 16.860 2494.250 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1543.340 0.300 1544.540 ;
=======
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1773.905 2493.645 1774.075 2496.875 ;
      LAYER mcon ;
        RECT 1773.905 2496.705 1774.075 2496.875 ;
      LAYER met1 ;
        RECT 1773.830 2496.860 1774.150 2496.920 ;
        RECT 1773.635 2496.720 1774.150 2496.860 ;
        RECT 1773.830 2496.660 1774.150 2496.720 ;
        RECT 26.750 2493.800 27.070 2493.860 ;
        RECT 1773.845 2493.800 1774.135 2493.845 ;
        RECT 26.750 2493.660 1774.135 2493.800 ;
        RECT 26.750 2493.600 27.070 2493.660 ;
        RECT 1773.845 2493.615 1774.135 2493.660 ;
        RECT 13.870 1330.660 14.190 1330.720 ;
        RECT 26.750 1330.660 27.070 1330.720 ;
        RECT 13.870 1330.520 27.070 1330.660 ;
        RECT 13.870 1330.460 14.190 1330.520 ;
        RECT 26.750 1330.460 27.070 1330.520 ;
      LAYER via ;
        RECT 1773.860 2496.660 1774.120 2496.920 ;
        RECT 26.780 2493.600 27.040 2493.860 ;
        RECT 13.900 1330.460 14.160 1330.720 ;
        RECT 26.780 1330.460 27.040 1330.720 ;
      LAYER met2 ;
        RECT 1773.860 2496.690 1774.120 2496.950 ;
        RECT 1774.310 2496.690 1774.590 2500.000 ;
        RECT 1773.860 2496.630 1774.590 2496.690 ;
        RECT 1773.920 2496.550 1774.590 2496.630 ;
        RECT 1774.310 2496.000 1774.590 2496.550 ;
        RECT 26.780 2493.570 27.040 2493.890 ;
        RECT 26.840 1330.750 26.980 2493.570 ;
        RECT 13.900 1330.430 14.160 1330.750 ;
        RECT 26.780 1330.430 27.040 1330.750 ;
        RECT 13.960 1328.565 14.100 1330.430 ;
        RECT 13.890 1328.195 14.170 1328.565 ;
      LAYER via2 ;
        RECT 13.890 1328.240 14.170 1328.520 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1327.780 0.300 1328.980 ;
=======
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 13.865 1328.530 14.195 1328.545 ;
        RECT -4.800 1328.230 14.195 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 13.865 1328.215 14.195 1328.230 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1794.145 2492.965 1794.315 2496.875 ;
      LAYER mcon ;
        RECT 1794.145 2496.705 1794.315 2496.875 ;
      LAYER met1 ;
        RECT 1794.070 2496.860 1794.390 2496.920 ;
        RECT 1793.875 2496.720 1794.390 2496.860 ;
        RECT 1794.070 2496.660 1794.390 2496.720 ;
        RECT 25.830 2493.120 26.150 2493.180 ;
        RECT 1794.085 2493.120 1794.375 2493.165 ;
        RECT 25.830 2492.980 1794.375 2493.120 ;
        RECT 25.830 2492.920 26.150 2492.980 ;
        RECT 1794.085 2492.935 1794.375 2492.980 ;
        RECT 13.870 1115.440 14.190 1115.500 ;
        RECT 25.830 1115.440 26.150 1115.500 ;
        RECT 13.870 1115.300 26.150 1115.440 ;
        RECT 13.870 1115.240 14.190 1115.300 ;
        RECT 25.830 1115.240 26.150 1115.300 ;
      LAYER via ;
        RECT 1794.100 2496.660 1794.360 2496.920 ;
        RECT 25.860 2492.920 26.120 2493.180 ;
        RECT 13.900 1115.240 14.160 1115.500 ;
        RECT 25.860 1115.240 26.120 1115.500 ;
      LAYER met2 ;
        RECT 1794.100 2496.690 1794.360 2496.950 ;
        RECT 1794.550 2496.690 1794.830 2500.000 ;
        RECT 1794.100 2496.630 1794.830 2496.690 ;
        RECT 1794.160 2496.550 1794.830 2496.630 ;
        RECT 1794.550 2496.000 1794.830 2496.550 ;
        RECT 25.860 2492.890 26.120 2493.210 ;
        RECT 25.920 1115.530 26.060 2492.890 ;
        RECT 13.900 1115.210 14.160 1115.530 ;
        RECT 25.860 1115.210 26.120 1115.530 ;
        RECT 13.960 1113.005 14.100 1115.210 ;
        RECT 13.890 1112.635 14.170 1113.005 ;
      LAYER via2 ;
        RECT 13.890 1112.680 14.170 1112.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1112.220 0.300 1113.420 ;
=======
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 13.865 1112.970 14.195 1112.985 ;
        RECT -4.800 1112.670 14.195 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 13.865 1112.655 14.195 1112.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1812.545 2492.285 1812.715 2496.875 ;
      LAYER mcon ;
        RECT 1812.545 2496.705 1812.715 2496.875 ;
      LAYER met1 ;
        RECT 1812.470 2496.860 1812.790 2496.920 ;
        RECT 1812.275 2496.720 1812.790 2496.860 ;
        RECT 1812.470 2496.660 1812.790 2496.720 ;
        RECT 25.370 2492.440 25.690 2492.500 ;
        RECT 1812.485 2492.440 1812.775 2492.485 ;
        RECT 25.370 2492.300 1812.775 2492.440 ;
        RECT 25.370 2492.240 25.690 2492.300 ;
        RECT 1812.485 2492.255 1812.775 2492.300 ;
        RECT 13.870 899.200 14.190 899.260 ;
        RECT 25.370 899.200 25.690 899.260 ;
        RECT 13.870 899.060 25.690 899.200 ;
        RECT 13.870 899.000 14.190 899.060 ;
        RECT 25.370 899.000 25.690 899.060 ;
      LAYER via ;
        RECT 1812.500 2496.660 1812.760 2496.920 ;
        RECT 25.400 2492.240 25.660 2492.500 ;
        RECT 13.900 899.000 14.160 899.260 ;
        RECT 25.400 899.000 25.660 899.260 ;
      LAYER met2 ;
        RECT 1812.500 2496.690 1812.760 2496.950 ;
        RECT 1814.330 2496.690 1814.610 2500.000 ;
        RECT 1812.500 2496.630 1814.610 2496.690 ;
        RECT 1812.560 2496.550 1814.610 2496.630 ;
        RECT 1814.330 2496.000 1814.610 2496.550 ;
        RECT 25.400 2492.210 25.660 2492.530 ;
        RECT 25.460 899.290 25.600 2492.210 ;
        RECT 13.900 898.970 14.160 899.290 ;
        RECT 25.400 898.970 25.660 899.290 ;
        RECT 13.960 897.445 14.100 898.970 ;
        RECT 13.890 897.075 14.170 897.445 ;
      LAYER via2 ;
        RECT 13.890 897.120 14.170 897.400 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 896.660 0.300 897.860 ;
=======
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 13.865 897.410 14.195 897.425 ;
        RECT -4.800 897.110 14.195 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 13.865 897.095 14.195 897.110 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1832.785 2491.605 1832.955 2496.875 ;
      LAYER mcon ;
        RECT 1832.785 2496.705 1832.955 2496.875 ;
      LAYER met1 ;
        RECT 1832.710 2496.860 1833.030 2496.920 ;
        RECT 1832.515 2496.720 1833.030 2496.860 ;
        RECT 1832.710 2496.660 1833.030 2496.720 ;
        RECT 18.470 2491.760 18.790 2491.820 ;
        RECT 1832.725 2491.760 1833.015 2491.805 ;
        RECT 18.470 2491.620 1833.015 2491.760 ;
        RECT 18.470 2491.560 18.790 2491.620 ;
        RECT 1832.725 2491.575 1833.015 2491.620 ;
      LAYER via ;
        RECT 1832.740 2496.660 1833.000 2496.920 ;
        RECT 18.500 2491.560 18.760 2491.820 ;
      LAYER met2 ;
        RECT 1832.740 2496.690 1833.000 2496.950 ;
        RECT 1834.110 2496.690 1834.390 2500.000 ;
        RECT 1832.740 2496.630 1834.390 2496.690 ;
        RECT 1832.800 2496.550 1834.390 2496.630 ;
        RECT 1834.110 2496.000 1834.390 2496.550 ;
        RECT 18.500 2491.530 18.760 2491.850 ;
        RECT 18.560 681.885 18.700 2491.530 ;
        RECT 18.490 681.515 18.770 681.885 ;
      LAYER via2 ;
        RECT 18.490 681.560 18.770 681.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 681.100 0.300 682.300 ;
=======
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 18.465 681.850 18.795 681.865 ;
        RECT -4.800 681.550 18.795 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 18.465 681.535 18.795 681.550 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1852.105 2490.925 1852.275 2496.875 ;
      LAYER mcon ;
        RECT 1852.105 2496.705 1852.275 2496.875 ;
      LAYER met1 ;
        RECT 1852.030 2496.860 1852.350 2496.920 ;
        RECT 1851.835 2496.720 1852.350 2496.860 ;
        RECT 1852.030 2496.660 1852.350 2496.720 ;
        RECT 24.450 2491.080 24.770 2491.140 ;
        RECT 1852.045 2491.080 1852.335 2491.125 ;
        RECT 24.450 2490.940 1852.335 2491.080 ;
        RECT 24.450 2490.880 24.770 2490.940 ;
        RECT 1852.045 2490.895 1852.335 2490.940 ;
        RECT 13.870 466.380 14.190 466.440 ;
        RECT 24.450 466.380 24.770 466.440 ;
        RECT 13.870 466.240 24.770 466.380 ;
        RECT 13.870 466.180 14.190 466.240 ;
        RECT 24.450 466.180 24.770 466.240 ;
      LAYER via ;
        RECT 1852.060 2496.660 1852.320 2496.920 ;
        RECT 24.480 2490.880 24.740 2491.140 ;
        RECT 13.900 466.180 14.160 466.440 ;
        RECT 24.480 466.180 24.740 466.440 ;
      LAYER met2 ;
        RECT 1852.060 2496.690 1852.320 2496.950 ;
        RECT 1853.890 2496.690 1854.170 2500.000 ;
        RECT 1852.060 2496.630 1854.170 2496.690 ;
        RECT 1852.120 2496.550 1854.170 2496.630 ;
        RECT 1853.890 2496.000 1854.170 2496.550 ;
        RECT 24.480 2490.850 24.740 2491.170 ;
        RECT 24.540 466.470 24.680 2490.850 ;
        RECT 13.900 466.325 14.160 466.470 ;
        RECT 13.890 465.955 14.170 466.325 ;
        RECT 24.480 466.150 24.740 466.470 ;
      LAYER via2 ;
        RECT 13.890 466.000 14.170 466.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 465.540 0.300 466.740 ;
=======
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 13.865 466.290 14.195 466.305 ;
        RECT -4.800 465.990 14.195 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 13.865 465.975 14.195 465.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23.990 2498.220 24.310 2498.280 ;
        RECT 1872.270 2498.220 1872.590 2498.280 ;
        RECT 23.990 2498.080 1872.590 2498.220 ;
        RECT 23.990 2498.020 24.310 2498.080 ;
        RECT 1872.270 2498.020 1872.590 2498.080 ;
        RECT 13.870 252.520 14.190 252.580 ;
        RECT 23.990 252.520 24.310 252.580 ;
        RECT 13.870 252.380 24.310 252.520 ;
        RECT 13.870 252.320 14.190 252.380 ;
        RECT 23.990 252.320 24.310 252.380 ;
      LAYER via ;
        RECT 24.020 2498.020 24.280 2498.280 ;
        RECT 1872.300 2498.020 1872.560 2498.280 ;
        RECT 13.900 252.320 14.160 252.580 ;
        RECT 24.020 252.320 24.280 252.580 ;
      LAYER met2 ;
        RECT 24.020 2497.990 24.280 2498.310 ;
        RECT 1872.300 2498.050 1872.560 2498.310 ;
        RECT 1873.670 2498.050 1873.950 2500.000 ;
        RECT 1872.300 2497.990 1873.950 2498.050 ;
        RECT 24.080 252.610 24.220 2497.990 ;
        RECT 1872.360 2497.910 1873.950 2497.990 ;
        RECT 1873.670 2496.000 1873.950 2497.910 ;
        RECT 13.900 252.290 14.160 252.610 ;
        RECT 24.020 252.290 24.280 252.610 ;
        RECT 13.960 250.765 14.100 252.290 ;
        RECT 13.890 250.395 14.170 250.765 ;
      LAYER via2 ;
        RECT 13.890 250.440 14.170 250.720 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 249.980 0.300 251.180 ;
=======
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 13.865 250.730 14.195 250.745 ;
        RECT -4.800 250.430 14.195 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 13.865 250.415 14.195 250.430 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 2514.795 17.390 2515.165 ;
        RECT 1893.450 2514.795 1893.730 2515.165 ;
        RECT 17.180 35.885 17.320 2514.795 ;
        RECT 1893.520 2500.000 1893.660 2514.795 ;
        RECT 1893.450 2496.000 1893.730 2500.000 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 17.110 2514.840 17.390 2515.120 ;
        RECT 1893.450 2514.840 1893.730 2515.120 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 35.100 0.300 36.300 ;
=======
        RECT 17.085 2515.130 17.415 2515.145 ;
        RECT 1893.425 2515.130 1893.755 2515.145 ;
        RECT 17.085 2514.830 1893.755 2515.130 ;
        RECT 17.085 2514.815 17.415 2514.830 ;
        RECT 1893.425 2514.815 1893.755 2514.830 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2608.270 906.000 2608.590 906.060 ;
        RECT 2632.650 906.000 2632.970 906.060 ;
        RECT 2608.270 905.860 2632.970 906.000 ;
        RECT 2608.270 905.800 2608.590 905.860 ;
        RECT 2632.650 905.800 2632.970 905.860 ;
        RECT 2511.670 905.320 2511.990 905.380 ;
        RECT 2549.850 905.320 2550.170 905.380 ;
        RECT 2511.670 905.180 2550.170 905.320 ;
        RECT 2511.670 905.120 2511.990 905.180 ;
        RECT 2549.850 905.120 2550.170 905.180 ;
        RECT 1593.970 904.980 1594.290 905.040 ;
        RECT 1607.770 904.980 1608.090 905.040 ;
        RECT 1593.970 904.840 1608.090 904.980 ;
        RECT 1593.970 904.780 1594.290 904.840 ;
        RECT 1607.770 904.780 1608.090 904.840 ;
        RECT 1798.670 904.980 1798.990 905.040 ;
        RECT 1811.550 904.980 1811.870 905.040 ;
        RECT 1798.670 904.840 1811.870 904.980 ;
        RECT 1798.670 904.780 1798.990 904.840 ;
        RECT 1811.550 904.780 1811.870 904.840 ;
        RECT 1702.070 904.640 1702.390 904.700 ;
        RECT 1714.490 904.640 1714.810 904.700 ;
        RECT 1702.070 904.500 1714.810 904.640 ;
        RECT 1702.070 904.440 1702.390 904.500 ;
        RECT 1714.490 904.440 1714.810 904.500 ;
        RECT 1895.270 904.640 1895.590 904.700 ;
        RECT 1897.570 904.640 1897.890 904.700 ;
        RECT 1895.270 904.500 1897.890 904.640 ;
        RECT 1895.270 904.440 1895.590 904.500 ;
        RECT 1897.570 904.440 1897.890 904.500 ;
      LAYER via ;
        RECT 2608.300 905.800 2608.560 906.060 ;
        RECT 2632.680 905.800 2632.940 906.060 ;
        RECT 2511.700 905.120 2511.960 905.380 ;
        RECT 2549.880 905.120 2550.140 905.380 ;
        RECT 1594.000 904.780 1594.260 905.040 ;
        RECT 1607.800 904.780 1608.060 905.040 ;
        RECT 1798.700 904.780 1798.960 905.040 ;
        RECT 1811.580 904.780 1811.840 905.040 ;
        RECT 1702.100 904.440 1702.360 904.700 ;
        RECT 1714.520 904.440 1714.780 904.700 ;
        RECT 1895.300 904.440 1895.560 904.700 ;
        RECT 1897.600 904.440 1897.860 904.700 ;
      LAYER met2 ;
        RECT 1219.090 2498.050 1219.370 2500.000 ;
        RECT 1220.010 2498.050 1220.290 2498.165 ;
        RECT 1219.090 2497.910 1220.290 2498.050 ;
        RECT 1219.090 2496.000 1219.370 2497.910 ;
        RECT 1220.010 2497.795 1220.290 2497.910 ;
        RECT 2680.510 906.595 2680.790 906.965 ;
        RECT 1296.830 905.915 1297.110 906.285 ;
        RECT 2574.250 906.170 2574.530 906.285 ;
        RECT 2573.400 906.030 2574.530 906.170 ;
        RECT 1296.900 905.605 1297.040 905.915 ;
        RECT 1296.830 905.235 1297.110 905.605 ;
        RECT 2511.690 905.235 2511.970 905.605 ;
        RECT 2511.700 905.090 2511.960 905.235 ;
        RECT 2549.880 905.090 2550.140 905.410 ;
        RECT 1594.000 904.925 1594.260 905.070 ;
        RECT 1607.800 904.925 1608.060 905.070 ;
        RECT 1798.700 904.925 1798.960 905.070 ;
        RECT 1811.580 904.925 1811.840 905.070 ;
        RECT 1593.990 904.555 1594.270 904.925 ;
        RECT 1607.790 904.555 1608.070 904.925 ;
        RECT 1702.090 904.555 1702.370 904.925 ;
        RECT 1714.510 904.555 1714.790 904.925 ;
        RECT 1798.690 904.555 1798.970 904.925 ;
        RECT 1811.570 904.555 1811.850 904.925 ;
        RECT 1895.290 904.555 1895.570 904.925 ;
        RECT 1897.590 904.555 1897.870 904.925 ;
        RECT 1993.730 904.810 1994.010 904.925 ;
        RECT 1994.650 904.810 1994.930 904.925 ;
        RECT 1993.730 904.670 1994.930 904.810 ;
        RECT 1993.730 904.555 1994.010 904.670 ;
        RECT 1994.650 904.555 1994.930 904.670 ;
        RECT 1702.100 904.410 1702.360 904.555 ;
        RECT 1714.520 904.410 1714.780 904.555 ;
        RECT 1895.300 904.410 1895.560 904.555 ;
        RECT 1897.600 904.410 1897.860 904.555 ;
        RECT 2549.940 904.245 2550.080 905.090 ;
        RECT 2573.400 904.925 2573.540 906.030 ;
        RECT 2574.250 905.915 2574.530 906.030 ;
        RECT 2608.290 905.915 2608.570 906.285 ;
        RECT 2608.300 905.770 2608.560 905.915 ;
        RECT 2632.680 905.770 2632.940 906.090 ;
        RECT 2632.740 905.605 2632.880 905.770 ;
        RECT 2680.580 905.605 2680.720 906.595 ;
        RECT 2632.670 905.235 2632.950 905.605 ;
        RECT 2680.510 905.235 2680.790 905.605 ;
        RECT 2573.330 904.555 2573.610 904.925 ;
        RECT 2549.870 903.875 2550.150 904.245 ;
      LAYER via2 ;
        RECT 1220.010 2497.840 1220.290 2498.120 ;
        RECT 2680.510 906.640 2680.790 906.920 ;
        RECT 1296.830 905.960 1297.110 906.240 ;
        RECT 1296.830 905.280 1297.110 905.560 ;
        RECT 2511.690 905.280 2511.970 905.560 ;
        RECT 1593.990 904.600 1594.270 904.880 ;
        RECT 1607.790 904.600 1608.070 904.880 ;
        RECT 1702.090 904.600 1702.370 904.880 ;
        RECT 1714.510 904.600 1714.790 904.880 ;
        RECT 1798.690 904.600 1798.970 904.880 ;
        RECT 1811.570 904.600 1811.850 904.880 ;
        RECT 1895.290 904.600 1895.570 904.880 ;
        RECT 1897.590 904.600 1897.870 904.880 ;
        RECT 1993.730 904.600 1994.010 904.880 ;
        RECT 1994.650 904.600 1994.930 904.880 ;
        RECT 2574.250 905.960 2574.530 906.240 ;
        RECT 2608.290 905.960 2608.570 906.240 ;
        RECT 2632.670 905.280 2632.950 905.560 ;
        RECT 2680.510 905.280 2680.790 905.560 ;
        RECT 2573.330 904.600 2573.610 904.880 ;
        RECT 2549.870 903.920 2550.150 904.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 908.900 2924.800 910.100 ;
=======
        RECT 1219.985 2498.140 1220.315 2498.145 ;
        RECT 1219.985 2498.130 1220.570 2498.140 ;
        RECT 1219.985 2497.830 1220.770 2498.130 ;
        RECT 1219.985 2497.820 1220.570 2497.830 ;
        RECT 1219.985 2497.815 1220.315 2497.820 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2916.710 909.350 2924.800 909.650 ;
        RECT 2656.310 906.930 2656.690 906.940 ;
        RECT 2680.485 906.930 2680.815 906.945 ;
        RECT 2656.310 906.630 2680.815 906.930 ;
        RECT 2656.310 906.620 2656.690 906.630 ;
        RECT 2680.485 906.615 2680.815 906.630 ;
        RECT 1296.805 906.250 1297.135 906.265 ;
        RECT 2574.225 906.250 2574.555 906.265 ;
        RECT 2608.265 906.250 2608.595 906.265 ;
        RECT 1296.805 905.950 1321.730 906.250 ;
        RECT 1296.805 905.935 1297.135 905.950 ;
        RECT 1220.190 905.570 1220.570 905.580 ;
        RECT 1296.805 905.570 1297.135 905.585 ;
        RECT 1220.190 905.270 1297.135 905.570 ;
        RECT 1321.430 905.570 1321.730 905.950 ;
        RECT 2574.225 905.950 2608.595 906.250 ;
        RECT 2574.225 905.935 2574.555 905.950 ;
        RECT 2608.265 905.935 2608.595 905.950 ;
        RECT 2511.665 905.570 2511.995 905.585 ;
        RECT 1321.430 905.270 1345.650 905.570 ;
        RECT 1220.190 905.260 1220.570 905.270 ;
        RECT 1296.805 905.255 1297.135 905.270 ;
        RECT 1345.350 904.900 1345.650 905.270 ;
        RECT 1473.230 905.270 1511.250 905.570 ;
        RECT 1345.310 904.580 1345.690 904.900 ;
        RECT 1346.230 904.890 1346.610 904.900 ;
        RECT 1473.230 904.890 1473.530 905.270 ;
        RECT 1346.230 904.590 1473.530 904.890 ;
        RECT 1346.230 904.580 1346.610 904.590 ;
        RECT 1510.950 904.210 1511.250 905.270 ;
        RECT 2090.550 905.270 2138.690 905.570 ;
        RECT 1593.965 904.890 1594.295 904.905 ;
        RECT 1559.710 904.590 1594.295 904.890 ;
        RECT 1559.710 904.210 1560.010 904.590 ;
        RECT 1593.965 904.575 1594.295 904.590 ;
        RECT 1607.765 904.890 1608.095 904.905 ;
        RECT 1702.065 904.890 1702.395 904.905 ;
        RECT 1607.765 904.590 1641.890 904.890 ;
        RECT 1607.765 904.575 1608.095 904.590 ;
        RECT 1510.950 903.910 1560.010 904.210 ;
        RECT 1641.590 904.210 1641.890 904.590 ;
        RECT 1656.310 904.590 1702.395 904.890 ;
        RECT 1656.310 904.210 1656.610 904.590 ;
        RECT 1702.065 904.575 1702.395 904.590 ;
        RECT 1714.485 904.890 1714.815 904.905 ;
        RECT 1798.665 904.890 1798.995 904.905 ;
        RECT 1714.485 904.590 1738.490 904.890 ;
        RECT 1714.485 904.575 1714.815 904.590 ;
        RECT 1641.590 903.910 1656.610 904.210 ;
        RECT 1738.190 904.210 1738.490 904.590 ;
        RECT 1752.910 904.590 1798.995 904.890 ;
        RECT 1752.910 904.210 1753.210 904.590 ;
        RECT 1798.665 904.575 1798.995 904.590 ;
        RECT 1811.545 904.890 1811.875 904.905 ;
        RECT 1895.265 904.890 1895.595 904.905 ;
        RECT 1811.545 904.590 1835.090 904.890 ;
        RECT 1811.545 904.575 1811.875 904.590 ;
        RECT 1738.190 903.910 1753.210 904.210 ;
        RECT 1834.790 904.210 1835.090 904.590 ;
        RECT 1849.510 904.590 1895.595 904.890 ;
        RECT 1849.510 904.210 1849.810 904.590 ;
        RECT 1895.265 904.575 1895.595 904.590 ;
        RECT 1897.565 904.890 1897.895 904.905 ;
        RECT 1993.705 904.890 1994.035 904.905 ;
        RECT 1897.565 904.590 1931.690 904.890 ;
        RECT 1897.565 904.575 1897.895 904.590 ;
        RECT 1834.790 903.910 1849.810 904.210 ;
        RECT 1931.390 904.210 1931.690 904.590 ;
        RECT 1946.110 904.590 1994.035 904.890 ;
        RECT 1946.110 904.210 1946.410 904.590 ;
        RECT 1993.705 904.575 1994.035 904.590 ;
        RECT 1994.625 904.890 1994.955 904.905 ;
        RECT 1994.625 904.590 2042.090 904.890 ;
        RECT 1994.625 904.575 1994.955 904.590 ;
        RECT 1931.390 903.910 1946.410 904.210 ;
        RECT 2041.790 904.210 2042.090 904.590 ;
        RECT 2090.550 904.210 2090.850 905.270 ;
        RECT 2041.790 903.910 2090.850 904.210 ;
        RECT 2138.390 904.210 2138.690 905.270 ;
        RECT 2187.150 905.270 2235.290 905.570 ;
        RECT 2187.150 904.210 2187.450 905.270 ;
        RECT 2138.390 903.910 2187.450 904.210 ;
        RECT 2234.990 904.210 2235.290 905.270 ;
        RECT 2283.750 905.270 2331.890 905.570 ;
        RECT 2283.750 904.210 2284.050 905.270 ;
        RECT 2234.990 903.910 2284.050 904.210 ;
        RECT 2331.590 904.210 2331.890 905.270 ;
        RECT 2352.750 905.270 2400.890 905.570 ;
        RECT 2352.750 904.210 2353.050 905.270 ;
        RECT 2331.590 903.910 2353.050 904.210 ;
        RECT 2400.590 904.210 2400.890 905.270 ;
        RECT 2401.510 905.270 2449.650 905.570 ;
        RECT 2401.510 904.210 2401.810 905.270 ;
        RECT 2449.350 904.890 2449.650 905.270 ;
        RECT 2498.110 905.270 2511.995 905.570 ;
        RECT 2449.350 904.590 2497.490 904.890 ;
        RECT 2400.590 903.910 2401.810 904.210 ;
        RECT 2497.190 904.210 2497.490 904.590 ;
        RECT 2498.110 904.210 2498.410 905.270 ;
        RECT 2511.665 905.255 2511.995 905.270 ;
        RECT 2632.645 905.570 2632.975 905.585 ;
        RECT 2656.310 905.570 2656.690 905.580 ;
        RECT 2632.645 905.270 2656.690 905.570 ;
        RECT 2632.645 905.255 2632.975 905.270 ;
        RECT 2656.310 905.260 2656.690 905.270 ;
        RECT 2680.485 905.570 2680.815 905.585 ;
        RECT 2680.485 905.270 2739.450 905.570 ;
        RECT 2680.485 905.255 2680.815 905.270 ;
        RECT 2573.305 904.890 2573.635 904.905 ;
        RECT 2559.750 904.590 2573.635 904.890 ;
        RECT 2739.150 904.890 2739.450 905.270 ;
        RECT 2787.910 905.270 2836.050 905.570 ;
        RECT 2739.150 904.590 2787.290 904.890 ;
        RECT 2497.190 903.910 2498.410 904.210 ;
        RECT 2549.845 904.210 2550.175 904.225 ;
        RECT 2559.750 904.210 2560.050 904.590 ;
        RECT 2573.305 904.575 2573.635 904.590 ;
        RECT 2549.845 903.910 2560.050 904.210 ;
        RECT 2786.990 904.210 2787.290 904.590 ;
        RECT 2787.910 904.210 2788.210 905.270 ;
        RECT 2835.750 904.890 2836.050 905.270 ;
        RECT 2916.710 904.890 2917.010 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
        RECT 2835.750 904.590 2883.890 904.890 ;
        RECT 2786.990 903.910 2788.210 904.210 ;
        RECT 2883.590 904.210 2883.890 904.590 ;
        RECT 2884.510 904.590 2917.010 904.890 ;
        RECT 2884.510 904.210 2884.810 904.590 ;
        RECT 2883.590 903.910 2884.810 904.210 ;
        RECT 2549.845 903.895 2550.175 903.910 ;
      LAYER via3 ;
        RECT 1220.220 2497.820 1220.540 2498.140 ;
        RECT 2656.340 906.620 2656.660 906.940 ;
        RECT 1220.220 905.260 1220.540 905.580 ;
        RECT 1345.340 904.580 1345.660 904.900 ;
        RECT 1346.260 904.580 1346.580 904.900 ;
        RECT 2656.340 905.260 2656.660 905.580 ;
      LAYER met4 ;
        RECT 1220.215 2497.815 1220.545 2498.145 ;
        RECT 1220.230 905.585 1220.530 2497.815 ;
        RECT 2656.335 906.615 2656.665 906.945 ;
        RECT 2656.350 905.585 2656.650 906.615 ;
        RECT 1220.215 905.255 1220.545 905.585 ;
        RECT 2656.335 905.255 2656.665 905.585 ;
        RECT 1345.335 904.575 1345.665 904.905 ;
        RECT 1346.255 904.575 1346.585 904.905 ;
        RECT 1345.350 902.850 1345.650 904.575 ;
        RECT 1346.270 902.850 1346.570 904.575 ;
        RECT 1345.350 902.550 1346.570 902.850 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1351.550 1139.920 1351.870 1139.980 ;
        RECT 1393.410 1139.920 1393.730 1139.980 ;
        RECT 1351.550 1139.780 1393.730 1139.920 ;
        RECT 1351.550 1139.720 1351.870 1139.780 ;
        RECT 1393.410 1139.720 1393.730 1139.780 ;
        RECT 1798.670 1139.580 1798.990 1139.640 ;
        RECT 1811.550 1139.580 1811.870 1139.640 ;
        RECT 1798.670 1139.440 1811.870 1139.580 ;
        RECT 1798.670 1139.380 1798.990 1139.440 ;
        RECT 1811.550 1139.380 1811.870 1139.440 ;
        RECT 2090.310 1139.580 2090.630 1139.640 ;
        RECT 2124.810 1139.580 2125.130 1139.640 ;
        RECT 2090.310 1139.440 2125.130 1139.580 ;
        RECT 2090.310 1139.380 2090.630 1139.440 ;
        RECT 2124.810 1139.380 2125.130 1139.440 ;
        RECT 1606.390 1139.240 1606.710 1139.300 ;
        RECT 1607.770 1139.240 1608.090 1139.300 ;
        RECT 1606.390 1139.100 1608.090 1139.240 ;
        RECT 1606.390 1139.040 1606.710 1139.100 ;
        RECT 1607.770 1139.040 1608.090 1139.100 ;
        RECT 1702.070 1139.240 1702.390 1139.300 ;
        RECT 1714.490 1139.240 1714.810 1139.300 ;
        RECT 1702.070 1139.100 1714.810 1139.240 ;
        RECT 1702.070 1139.040 1702.390 1139.100 ;
        RECT 1714.490 1139.040 1714.810 1139.100 ;
        RECT 1932.070 1138.900 1932.390 1138.960 ;
        RECT 1946.330 1138.900 1946.650 1138.960 ;
        RECT 1932.070 1138.760 1946.650 1138.900 ;
        RECT 1932.070 1138.700 1932.390 1138.760 ;
        RECT 1946.330 1138.700 1946.650 1138.760 ;
      LAYER via ;
        RECT 1351.580 1139.720 1351.840 1139.980 ;
        RECT 1393.440 1139.720 1393.700 1139.980 ;
        RECT 1798.700 1139.380 1798.960 1139.640 ;
        RECT 1811.580 1139.380 1811.840 1139.640 ;
        RECT 2090.340 1139.380 2090.600 1139.640 ;
        RECT 2124.840 1139.380 2125.100 1139.640 ;
        RECT 1606.420 1139.040 1606.680 1139.300 ;
        RECT 1607.800 1139.040 1608.060 1139.300 ;
        RECT 1702.100 1139.040 1702.360 1139.300 ;
        RECT 1714.520 1139.040 1714.780 1139.300 ;
        RECT 1932.100 1138.700 1932.360 1138.960 ;
        RECT 1946.360 1138.700 1946.620 1138.960 ;
      LAYER met2 ;
        RECT 1238.870 2498.050 1239.150 2500.000 ;
        RECT 1240.710 2498.050 1240.990 2498.165 ;
        RECT 1238.870 2497.910 1240.990 2498.050 ;
        RECT 1238.870 2496.000 1239.150 2497.910 ;
        RECT 1240.710 2497.795 1240.990 2497.910 ;
        RECT 2028.230 1141.195 2028.510 1141.565 ;
        RECT 1351.570 1140.515 1351.850 1140.885 ;
        RECT 1351.640 1140.010 1351.780 1140.515 ;
        RECT 1351.580 1139.690 1351.840 1140.010 ;
        RECT 1393.440 1139.690 1393.700 1140.010 ;
        RECT 1946.350 1139.835 1946.630 1140.205 ;
        RECT 1393.500 1139.525 1393.640 1139.690 ;
        RECT 1798.700 1139.525 1798.960 1139.670 ;
        RECT 1811.580 1139.525 1811.840 1139.670 ;
        RECT 1393.430 1139.155 1393.710 1139.525 ;
        RECT 1606.410 1139.155 1606.690 1139.525 ;
        RECT 1607.790 1139.155 1608.070 1139.525 ;
        RECT 1702.090 1139.155 1702.370 1139.525 ;
        RECT 1714.510 1139.155 1714.790 1139.525 ;
        RECT 1798.690 1139.155 1798.970 1139.525 ;
        RECT 1811.570 1139.155 1811.850 1139.525 ;
        RECT 1895.290 1139.155 1895.570 1139.525 ;
        RECT 1606.420 1139.010 1606.680 1139.155 ;
        RECT 1607.800 1139.010 1608.060 1139.155 ;
        RECT 1702.100 1139.010 1702.360 1139.155 ;
        RECT 1714.520 1139.010 1714.780 1139.155 ;
        RECT 1895.360 1137.485 1895.500 1139.155 ;
        RECT 1946.420 1138.990 1946.560 1139.835 ;
        RECT 2028.300 1139.525 2028.440 1141.195 ;
        RECT 2052.610 1140.515 2052.890 1140.885 ;
        RECT 2028.230 1139.155 2028.510 1139.525 ;
        RECT 1932.100 1138.845 1932.360 1138.990 ;
        RECT 1932.090 1138.475 1932.370 1138.845 ;
        RECT 1946.360 1138.670 1946.620 1138.990 ;
        RECT 2052.680 1138.845 2052.820 1140.515 ;
        RECT 2124.830 1139.835 2125.110 1140.205 ;
        RECT 2124.900 1139.670 2125.040 1139.835 ;
        RECT 2090.340 1139.525 2090.600 1139.670 ;
        RECT 2090.330 1139.155 2090.610 1139.525 ;
        RECT 2124.840 1139.350 2125.100 1139.670 ;
        RECT 2052.610 1138.475 2052.890 1138.845 ;
        RECT 1895.290 1137.115 1895.570 1137.485 ;
      LAYER via2 ;
        RECT 1240.710 2497.840 1240.990 2498.120 ;
        RECT 2028.230 1141.240 2028.510 1141.520 ;
        RECT 1351.570 1140.560 1351.850 1140.840 ;
        RECT 1946.350 1139.880 1946.630 1140.160 ;
        RECT 1393.430 1139.200 1393.710 1139.480 ;
        RECT 1606.410 1139.200 1606.690 1139.480 ;
        RECT 1607.790 1139.200 1608.070 1139.480 ;
        RECT 1702.090 1139.200 1702.370 1139.480 ;
        RECT 1714.510 1139.200 1714.790 1139.480 ;
        RECT 1798.690 1139.200 1798.970 1139.480 ;
        RECT 1811.570 1139.200 1811.850 1139.480 ;
        RECT 1895.290 1139.200 1895.570 1139.480 ;
        RECT 2052.610 1140.560 2052.890 1140.840 ;
        RECT 2028.230 1139.200 2028.510 1139.480 ;
        RECT 1932.090 1138.520 1932.370 1138.800 ;
        RECT 2124.830 1139.880 2125.110 1140.160 ;
        RECT 2090.330 1139.200 2090.610 1139.480 ;
        RECT 2052.610 1138.520 2052.890 1138.800 ;
        RECT 1895.290 1137.160 1895.570 1137.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1143.500 2924.800 1144.700 ;
=======
        RECT 1240.685 2498.130 1241.015 2498.145 ;
        RECT 1241.350 2498.130 1241.730 2498.140 ;
        RECT 1240.685 2497.830 1241.730 2498.130 ;
        RECT 1240.685 2497.815 1241.015 2497.830 ;
        RECT 1241.350 2497.820 1241.730 2497.830 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2916.710 1143.950 2924.800 1144.250 ;
        RECT 1980.110 1141.530 1980.490 1141.540 ;
        RECT 2028.205 1141.530 2028.535 1141.545 ;
        RECT 1269.910 1141.230 1321.730 1141.530 ;
        RECT 1269.910 1140.850 1270.210 1141.230 ;
        RECT 1268.990 1140.550 1270.210 1140.850 ;
        RECT 1321.430 1140.850 1321.730 1141.230 ;
        RECT 1980.110 1141.230 2028.535 1141.530 ;
        RECT 1980.110 1141.220 1980.490 1141.230 ;
        RECT 2028.205 1141.215 2028.535 1141.230 ;
        RECT 1351.545 1140.850 1351.875 1140.865 ;
        RECT 2052.585 1140.850 2052.915 1140.865 ;
        RECT 1321.430 1140.550 1351.875 1140.850 ;
        RECT 1241.350 1140.170 1241.730 1140.180 ;
        RECT 1268.990 1140.170 1269.290 1140.550 ;
        RECT 1351.545 1140.535 1351.875 1140.550 ;
        RECT 2028.910 1140.550 2052.915 1140.850 ;
        RECT 1946.325 1140.170 1946.655 1140.185 ;
        RECT 1980.110 1140.170 1980.490 1140.180 ;
        RECT 1241.350 1139.870 1269.290 1140.170 ;
        RECT 1451.840 1139.870 1511.250 1140.170 ;
        RECT 1241.350 1139.860 1241.730 1139.870 ;
        RECT 1393.405 1139.490 1393.735 1139.505 ;
        RECT 1451.840 1139.490 1452.140 1139.870 ;
        RECT 1393.405 1139.190 1452.140 1139.490 ;
        RECT 1393.405 1139.175 1393.735 1139.190 ;
        RECT 1510.950 1138.810 1511.250 1139.870 ;
        RECT 1946.325 1139.870 1980.490 1140.170 ;
        RECT 1946.325 1139.855 1946.655 1139.870 ;
        RECT 1980.110 1139.860 1980.490 1139.870 ;
        RECT 1606.385 1139.490 1606.715 1139.505 ;
        RECT 1559.710 1139.190 1606.715 1139.490 ;
        RECT 1559.710 1138.810 1560.010 1139.190 ;
        RECT 1606.385 1139.175 1606.715 1139.190 ;
        RECT 1607.765 1139.490 1608.095 1139.505 ;
        RECT 1702.065 1139.490 1702.395 1139.505 ;
        RECT 1607.765 1139.190 1641.890 1139.490 ;
        RECT 1607.765 1139.175 1608.095 1139.190 ;
        RECT 1510.950 1138.510 1560.010 1138.810 ;
        RECT 1641.590 1138.810 1641.890 1139.190 ;
        RECT 1656.310 1139.190 1702.395 1139.490 ;
        RECT 1656.310 1138.810 1656.610 1139.190 ;
        RECT 1702.065 1139.175 1702.395 1139.190 ;
        RECT 1714.485 1139.490 1714.815 1139.505 ;
        RECT 1798.665 1139.490 1798.995 1139.505 ;
        RECT 1714.485 1139.190 1738.490 1139.490 ;
        RECT 1714.485 1139.175 1714.815 1139.190 ;
        RECT 1641.590 1138.510 1656.610 1138.810 ;
        RECT 1738.190 1138.810 1738.490 1139.190 ;
        RECT 1752.910 1139.190 1798.995 1139.490 ;
        RECT 1752.910 1138.810 1753.210 1139.190 ;
        RECT 1798.665 1139.175 1798.995 1139.190 ;
        RECT 1811.545 1139.490 1811.875 1139.505 ;
        RECT 1895.265 1139.490 1895.595 1139.505 ;
        RECT 1811.545 1139.190 1835.090 1139.490 ;
        RECT 1811.545 1139.175 1811.875 1139.190 ;
        RECT 1738.190 1138.510 1753.210 1138.810 ;
        RECT 1834.790 1138.810 1835.090 1139.190 ;
        RECT 1849.510 1139.190 1895.595 1139.490 ;
        RECT 1849.510 1138.810 1849.810 1139.190 ;
        RECT 1895.265 1139.175 1895.595 1139.190 ;
        RECT 2028.205 1139.490 2028.535 1139.505 ;
        RECT 2028.910 1139.490 2029.210 1140.550 ;
        RECT 2052.585 1140.535 2052.915 1140.550 ;
        RECT 2124.805 1140.170 2125.135 1140.185 ;
        RECT 2124.805 1139.870 2159.850 1140.170 ;
        RECT 2124.805 1139.855 2125.135 1139.870 ;
        RECT 2090.305 1139.490 2090.635 1139.505 ;
        RECT 2028.205 1139.190 2029.210 1139.490 ;
        RECT 2076.750 1139.190 2090.635 1139.490 ;
        RECT 2159.550 1139.490 2159.850 1139.870 ;
        RECT 2208.310 1139.870 2256.450 1140.170 ;
        RECT 2159.550 1139.190 2207.690 1139.490 ;
        RECT 2028.205 1139.175 2028.535 1139.190 ;
        RECT 1932.065 1138.810 1932.395 1138.825 ;
        RECT 1834.790 1138.510 1849.810 1138.810 ;
        RECT 1931.390 1138.510 1932.395 1138.810 ;
        RECT 1895.265 1137.450 1895.595 1137.465 ;
        RECT 1931.390 1137.450 1931.690 1138.510 ;
        RECT 1932.065 1138.495 1932.395 1138.510 ;
        RECT 2052.585 1138.810 2052.915 1138.825 ;
        RECT 2076.750 1138.810 2077.050 1139.190 ;
        RECT 2090.305 1139.175 2090.635 1139.190 ;
        RECT 2052.585 1138.510 2077.050 1138.810 ;
        RECT 2207.390 1138.810 2207.690 1139.190 ;
        RECT 2208.310 1138.810 2208.610 1139.870 ;
        RECT 2256.150 1139.490 2256.450 1139.870 ;
        RECT 2304.910 1139.870 2353.050 1140.170 ;
        RECT 2256.150 1139.190 2304.290 1139.490 ;
        RECT 2207.390 1138.510 2208.610 1138.810 ;
        RECT 2303.990 1138.810 2304.290 1139.190 ;
        RECT 2304.910 1138.810 2305.210 1139.870 ;
        RECT 2352.750 1139.490 2353.050 1139.870 ;
        RECT 2401.510 1139.870 2449.650 1140.170 ;
        RECT 2352.750 1139.190 2400.890 1139.490 ;
        RECT 2303.990 1138.510 2305.210 1138.810 ;
        RECT 2400.590 1138.810 2400.890 1139.190 ;
        RECT 2401.510 1138.810 2401.810 1139.870 ;
        RECT 2449.350 1139.490 2449.650 1139.870 ;
        RECT 2498.110 1139.870 2546.250 1140.170 ;
        RECT 2449.350 1139.190 2497.490 1139.490 ;
        RECT 2400.590 1138.510 2401.810 1138.810 ;
        RECT 2497.190 1138.810 2497.490 1139.190 ;
        RECT 2498.110 1138.810 2498.410 1139.870 ;
        RECT 2545.950 1139.490 2546.250 1139.870 ;
        RECT 2594.710 1139.870 2642.850 1140.170 ;
        RECT 2545.950 1139.190 2594.090 1139.490 ;
        RECT 2497.190 1138.510 2498.410 1138.810 ;
        RECT 2593.790 1138.810 2594.090 1139.190 ;
        RECT 2594.710 1138.810 2595.010 1139.870 ;
        RECT 2642.550 1139.490 2642.850 1139.870 ;
        RECT 2691.310 1139.870 2739.450 1140.170 ;
        RECT 2642.550 1139.190 2690.690 1139.490 ;
        RECT 2593.790 1138.510 2595.010 1138.810 ;
        RECT 2690.390 1138.810 2690.690 1139.190 ;
        RECT 2691.310 1138.810 2691.610 1139.870 ;
        RECT 2739.150 1139.490 2739.450 1139.870 ;
        RECT 2787.910 1139.870 2836.050 1140.170 ;
        RECT 2739.150 1139.190 2787.290 1139.490 ;
        RECT 2690.390 1138.510 2691.610 1138.810 ;
        RECT 2786.990 1138.810 2787.290 1139.190 ;
        RECT 2787.910 1138.810 2788.210 1139.870 ;
        RECT 2835.750 1139.490 2836.050 1139.870 ;
        RECT 2916.710 1139.490 2917.010 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT 2835.750 1139.190 2883.890 1139.490 ;
        RECT 2786.990 1138.510 2788.210 1138.810 ;
        RECT 2883.590 1138.810 2883.890 1139.190 ;
        RECT 2884.510 1139.190 2917.010 1139.490 ;
        RECT 2884.510 1138.810 2884.810 1139.190 ;
        RECT 2883.590 1138.510 2884.810 1138.810 ;
        RECT 2052.585 1138.495 2052.915 1138.510 ;
        RECT 1895.265 1137.150 1931.690 1137.450 ;
        RECT 1895.265 1137.135 1895.595 1137.150 ;
      LAYER via3 ;
        RECT 1241.380 2497.820 1241.700 2498.140 ;
        RECT 1980.140 1141.220 1980.460 1141.540 ;
        RECT 1241.380 1139.860 1241.700 1140.180 ;
        RECT 1980.140 1139.860 1980.460 1140.180 ;
      LAYER met4 ;
        RECT 1241.375 2497.815 1241.705 2498.145 ;
        RECT 1241.390 1140.185 1241.690 2497.815 ;
        RECT 1980.135 1141.215 1980.465 1141.545 ;
        RECT 1980.150 1140.185 1980.450 1141.215 ;
        RECT 1241.375 1139.855 1241.705 1140.185 ;
        RECT 1980.135 1139.855 1980.465 1140.185 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1798.670 1374.180 1798.990 1374.240 ;
        RECT 1811.550 1374.180 1811.870 1374.240 ;
        RECT 1798.670 1374.040 1811.870 1374.180 ;
        RECT 1798.670 1373.980 1798.990 1374.040 ;
        RECT 1811.550 1373.980 1811.870 1374.040 ;
        RECT 2090.310 1374.180 2090.630 1374.240 ;
        RECT 2124.810 1374.180 2125.130 1374.240 ;
        RECT 2090.310 1374.040 2125.130 1374.180 ;
        RECT 2090.310 1373.980 2090.630 1374.040 ;
        RECT 2124.810 1373.980 2125.130 1374.040 ;
        RECT 1606.390 1373.840 1606.710 1373.900 ;
        RECT 1607.770 1373.840 1608.090 1373.900 ;
        RECT 1606.390 1373.700 1608.090 1373.840 ;
        RECT 1606.390 1373.640 1606.710 1373.700 ;
        RECT 1607.770 1373.640 1608.090 1373.700 ;
        RECT 1702.070 1373.840 1702.390 1373.900 ;
        RECT 1714.490 1373.840 1714.810 1373.900 ;
        RECT 1702.070 1373.700 1714.810 1373.840 ;
        RECT 1702.070 1373.640 1702.390 1373.700 ;
        RECT 1714.490 1373.640 1714.810 1373.700 ;
        RECT 1932.070 1373.500 1932.390 1373.560 ;
        RECT 1946.330 1373.500 1946.650 1373.560 ;
        RECT 1932.070 1373.360 1946.650 1373.500 ;
        RECT 1932.070 1373.300 1932.390 1373.360 ;
        RECT 1946.330 1373.300 1946.650 1373.360 ;
      LAYER via ;
        RECT 1798.700 1373.980 1798.960 1374.240 ;
        RECT 1811.580 1373.980 1811.840 1374.240 ;
        RECT 2090.340 1373.980 2090.600 1374.240 ;
        RECT 2124.840 1373.980 2125.100 1374.240 ;
        RECT 1606.420 1373.640 1606.680 1373.900 ;
        RECT 1607.800 1373.640 1608.060 1373.900 ;
        RECT 1702.100 1373.640 1702.360 1373.900 ;
        RECT 1714.520 1373.640 1714.780 1373.900 ;
        RECT 1932.100 1373.300 1932.360 1373.560 ;
        RECT 1946.360 1373.300 1946.620 1373.560 ;
      LAYER met2 ;
        RECT 1258.650 2498.050 1258.930 2500.000 ;
        RECT 1260.030 2498.050 1260.310 2498.165 ;
        RECT 1258.650 2497.910 1260.310 2498.050 ;
        RECT 1258.650 2496.000 1258.930 2497.910 ;
        RECT 1260.030 2497.795 1260.310 2497.910 ;
        RECT 2028.230 1375.795 2028.510 1376.165 ;
        RECT 1434.830 1375.115 1435.110 1375.485 ;
        RECT 1379.630 1374.435 1379.910 1374.805 ;
        RECT 1296.830 1374.010 1297.110 1374.125 ;
        RECT 1296.830 1373.870 1297.500 1374.010 ;
        RECT 1296.830 1373.755 1297.110 1373.870 ;
        RECT 1297.360 1373.445 1297.500 1373.870 ;
        RECT 1379.700 1373.445 1379.840 1374.435 ;
        RECT 1386.530 1373.755 1386.810 1374.125 ;
        RECT 1386.600 1373.445 1386.740 1373.755 ;
        RECT 1434.900 1373.445 1435.040 1375.115 ;
        RECT 1946.350 1374.435 1946.630 1374.805 ;
        RECT 1798.700 1374.125 1798.960 1374.270 ;
        RECT 1811.580 1374.125 1811.840 1374.270 ;
        RECT 1606.410 1373.755 1606.690 1374.125 ;
        RECT 1607.790 1373.755 1608.070 1374.125 ;
        RECT 1702.090 1373.755 1702.370 1374.125 ;
        RECT 1714.510 1373.755 1714.790 1374.125 ;
        RECT 1798.690 1373.755 1798.970 1374.125 ;
        RECT 1811.570 1373.755 1811.850 1374.125 ;
        RECT 1895.290 1373.755 1895.570 1374.125 ;
        RECT 1606.420 1373.610 1606.680 1373.755 ;
        RECT 1607.800 1373.610 1608.060 1373.755 ;
        RECT 1702.100 1373.610 1702.360 1373.755 ;
        RECT 1714.520 1373.610 1714.780 1373.755 ;
        RECT 1297.290 1373.075 1297.570 1373.445 ;
        RECT 1379.630 1373.075 1379.910 1373.445 ;
        RECT 1386.530 1373.075 1386.810 1373.445 ;
        RECT 1434.830 1373.075 1435.110 1373.445 ;
        RECT 1895.360 1372.085 1895.500 1373.755 ;
        RECT 1946.420 1373.590 1946.560 1374.435 ;
        RECT 2028.300 1374.125 2028.440 1375.795 ;
        RECT 2052.610 1375.115 2052.890 1375.485 ;
        RECT 2028.230 1373.755 2028.510 1374.125 ;
        RECT 1932.100 1373.445 1932.360 1373.590 ;
        RECT 1932.090 1373.075 1932.370 1373.445 ;
        RECT 1946.360 1373.270 1946.620 1373.590 ;
        RECT 2052.680 1373.445 2052.820 1375.115 ;
        RECT 2124.830 1374.435 2125.110 1374.805 ;
        RECT 2124.900 1374.270 2125.040 1374.435 ;
        RECT 2090.340 1374.125 2090.600 1374.270 ;
        RECT 2090.330 1373.755 2090.610 1374.125 ;
        RECT 2124.840 1373.950 2125.100 1374.270 ;
        RECT 2052.610 1373.075 2052.890 1373.445 ;
        RECT 1895.290 1371.715 1895.570 1372.085 ;
      LAYER via2 ;
        RECT 1260.030 2497.840 1260.310 2498.120 ;
        RECT 2028.230 1375.840 2028.510 1376.120 ;
        RECT 1434.830 1375.160 1435.110 1375.440 ;
        RECT 1379.630 1374.480 1379.910 1374.760 ;
        RECT 1296.830 1373.800 1297.110 1374.080 ;
        RECT 1386.530 1373.800 1386.810 1374.080 ;
        RECT 1946.350 1374.480 1946.630 1374.760 ;
        RECT 1606.410 1373.800 1606.690 1374.080 ;
        RECT 1607.790 1373.800 1608.070 1374.080 ;
        RECT 1702.090 1373.800 1702.370 1374.080 ;
        RECT 1714.510 1373.800 1714.790 1374.080 ;
        RECT 1798.690 1373.800 1798.970 1374.080 ;
        RECT 1811.570 1373.800 1811.850 1374.080 ;
        RECT 1895.290 1373.800 1895.570 1374.080 ;
        RECT 1297.290 1373.120 1297.570 1373.400 ;
        RECT 1379.630 1373.120 1379.910 1373.400 ;
        RECT 1386.530 1373.120 1386.810 1373.400 ;
        RECT 1434.830 1373.120 1435.110 1373.400 ;
        RECT 2052.610 1375.160 2052.890 1375.440 ;
        RECT 2028.230 1373.800 2028.510 1374.080 ;
        RECT 1932.090 1373.120 1932.370 1373.400 ;
        RECT 2124.830 1374.480 2125.110 1374.760 ;
        RECT 2090.330 1373.800 2090.610 1374.080 ;
        RECT 2052.610 1373.120 2052.890 1373.400 ;
        RECT 1895.290 1371.760 1895.570 1372.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1378.100 2924.800 1379.300 ;
=======
        RECT 1260.005 2498.130 1260.335 2498.145 ;
        RECT 1261.590 2498.130 1261.970 2498.140 ;
        RECT 1260.005 2497.830 1261.970 2498.130 ;
        RECT 1260.005 2497.815 1260.335 2497.830 ;
        RECT 1261.590 2497.820 1261.970 2497.830 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2916.710 1378.550 2924.800 1378.850 ;
        RECT 1980.110 1376.130 1980.490 1376.140 ;
        RECT 2028.205 1376.130 2028.535 1376.145 ;
        RECT 1980.110 1375.830 2028.535 1376.130 ;
        RECT 1980.110 1375.820 1980.490 1375.830 ;
        RECT 2028.205 1375.815 2028.535 1375.830 ;
        RECT 1386.710 1375.450 1387.090 1375.460 ;
        RECT 1434.805 1375.450 1435.135 1375.465 ;
        RECT 2052.585 1375.450 2052.915 1375.465 ;
        RECT 1386.710 1375.150 1435.135 1375.450 ;
        RECT 1386.710 1375.140 1387.090 1375.150 ;
        RECT 1434.805 1375.135 1435.135 1375.150 ;
        RECT 2028.910 1375.150 2052.915 1375.450 ;
        RECT 1331.510 1374.770 1331.890 1374.780 ;
        RECT 1379.605 1374.770 1379.935 1374.785 ;
        RECT 1331.510 1374.470 1379.935 1374.770 ;
        RECT 1331.510 1374.460 1331.890 1374.470 ;
        RECT 1379.605 1374.455 1379.935 1374.470 ;
        RECT 1441.910 1374.770 1442.290 1374.780 ;
        RECT 1946.325 1374.770 1946.655 1374.785 ;
        RECT 1980.110 1374.770 1980.490 1374.780 ;
        RECT 1441.910 1374.470 1562.770 1374.770 ;
        RECT 1441.910 1374.460 1442.290 1374.470 ;
        RECT 1261.590 1374.090 1261.970 1374.100 ;
        RECT 1296.805 1374.090 1297.135 1374.105 ;
        RECT 1261.590 1373.790 1297.135 1374.090 ;
        RECT 1261.590 1373.780 1261.970 1373.790 ;
        RECT 1296.805 1373.775 1297.135 1373.790 ;
        RECT 1386.505 1374.100 1386.835 1374.105 ;
        RECT 1386.505 1374.090 1387.090 1374.100 ;
        RECT 1562.470 1374.090 1562.770 1374.470 ;
        RECT 1946.325 1374.470 1980.490 1374.770 ;
        RECT 1946.325 1374.455 1946.655 1374.470 ;
        RECT 1980.110 1374.460 1980.490 1374.470 ;
        RECT 1606.385 1374.090 1606.715 1374.105 ;
        RECT 1386.505 1373.790 1387.470 1374.090 ;
        RECT 1562.470 1373.790 1606.715 1374.090 ;
        RECT 1386.505 1373.780 1387.090 1373.790 ;
        RECT 1386.505 1373.775 1386.835 1373.780 ;
        RECT 1606.385 1373.775 1606.715 1373.790 ;
        RECT 1607.765 1374.090 1608.095 1374.105 ;
        RECT 1702.065 1374.090 1702.395 1374.105 ;
        RECT 1607.765 1373.790 1641.890 1374.090 ;
        RECT 1607.765 1373.775 1608.095 1373.790 ;
        RECT 1297.265 1373.410 1297.595 1373.425 ;
        RECT 1331.510 1373.410 1331.890 1373.420 ;
        RECT 1297.265 1373.110 1331.890 1373.410 ;
        RECT 1297.265 1373.095 1297.595 1373.110 ;
        RECT 1331.510 1373.100 1331.890 1373.110 ;
        RECT 1379.605 1373.410 1379.935 1373.425 ;
        RECT 1386.505 1373.410 1386.835 1373.425 ;
        RECT 1379.605 1373.110 1386.835 1373.410 ;
        RECT 1379.605 1373.095 1379.935 1373.110 ;
        RECT 1386.505 1373.095 1386.835 1373.110 ;
        RECT 1434.805 1373.410 1435.135 1373.425 ;
        RECT 1441.910 1373.410 1442.290 1373.420 ;
        RECT 1434.805 1373.110 1442.290 1373.410 ;
        RECT 1641.590 1373.410 1641.890 1373.790 ;
        RECT 1656.310 1373.790 1702.395 1374.090 ;
        RECT 1656.310 1373.410 1656.610 1373.790 ;
        RECT 1702.065 1373.775 1702.395 1373.790 ;
        RECT 1714.485 1374.090 1714.815 1374.105 ;
        RECT 1798.665 1374.090 1798.995 1374.105 ;
        RECT 1714.485 1373.790 1738.490 1374.090 ;
        RECT 1714.485 1373.775 1714.815 1373.790 ;
        RECT 1641.590 1373.110 1656.610 1373.410 ;
        RECT 1738.190 1373.410 1738.490 1373.790 ;
        RECT 1752.910 1373.790 1798.995 1374.090 ;
        RECT 1752.910 1373.410 1753.210 1373.790 ;
        RECT 1798.665 1373.775 1798.995 1373.790 ;
        RECT 1811.545 1374.090 1811.875 1374.105 ;
        RECT 1895.265 1374.090 1895.595 1374.105 ;
        RECT 1811.545 1373.790 1835.090 1374.090 ;
        RECT 1811.545 1373.775 1811.875 1373.790 ;
        RECT 1738.190 1373.110 1753.210 1373.410 ;
        RECT 1834.790 1373.410 1835.090 1373.790 ;
        RECT 1849.510 1373.790 1895.595 1374.090 ;
        RECT 1849.510 1373.410 1849.810 1373.790 ;
        RECT 1895.265 1373.775 1895.595 1373.790 ;
        RECT 2028.205 1374.090 2028.535 1374.105 ;
        RECT 2028.910 1374.090 2029.210 1375.150 ;
        RECT 2052.585 1375.135 2052.915 1375.150 ;
        RECT 2124.805 1374.770 2125.135 1374.785 ;
        RECT 2124.805 1374.470 2159.850 1374.770 ;
        RECT 2124.805 1374.455 2125.135 1374.470 ;
        RECT 2090.305 1374.090 2090.635 1374.105 ;
        RECT 2028.205 1373.790 2029.210 1374.090 ;
        RECT 2076.750 1373.790 2090.635 1374.090 ;
        RECT 2159.550 1374.090 2159.850 1374.470 ;
        RECT 2208.310 1374.470 2256.450 1374.770 ;
        RECT 2159.550 1373.790 2207.690 1374.090 ;
        RECT 2028.205 1373.775 2028.535 1373.790 ;
        RECT 1932.065 1373.410 1932.395 1373.425 ;
        RECT 1834.790 1373.110 1849.810 1373.410 ;
        RECT 1931.390 1373.110 1932.395 1373.410 ;
        RECT 1434.805 1373.095 1435.135 1373.110 ;
        RECT 1441.910 1373.100 1442.290 1373.110 ;
        RECT 1895.265 1372.050 1895.595 1372.065 ;
        RECT 1931.390 1372.050 1931.690 1373.110 ;
        RECT 1932.065 1373.095 1932.395 1373.110 ;
        RECT 2052.585 1373.410 2052.915 1373.425 ;
        RECT 2076.750 1373.410 2077.050 1373.790 ;
        RECT 2090.305 1373.775 2090.635 1373.790 ;
        RECT 2052.585 1373.110 2077.050 1373.410 ;
        RECT 2207.390 1373.410 2207.690 1373.790 ;
        RECT 2208.310 1373.410 2208.610 1374.470 ;
        RECT 2256.150 1374.090 2256.450 1374.470 ;
        RECT 2304.910 1374.470 2353.050 1374.770 ;
        RECT 2256.150 1373.790 2304.290 1374.090 ;
        RECT 2207.390 1373.110 2208.610 1373.410 ;
        RECT 2303.990 1373.410 2304.290 1373.790 ;
        RECT 2304.910 1373.410 2305.210 1374.470 ;
        RECT 2352.750 1374.090 2353.050 1374.470 ;
        RECT 2401.510 1374.470 2449.650 1374.770 ;
        RECT 2352.750 1373.790 2400.890 1374.090 ;
        RECT 2303.990 1373.110 2305.210 1373.410 ;
        RECT 2400.590 1373.410 2400.890 1373.790 ;
        RECT 2401.510 1373.410 2401.810 1374.470 ;
        RECT 2449.350 1374.090 2449.650 1374.470 ;
        RECT 2498.110 1374.470 2546.250 1374.770 ;
        RECT 2449.350 1373.790 2497.490 1374.090 ;
        RECT 2400.590 1373.110 2401.810 1373.410 ;
        RECT 2497.190 1373.410 2497.490 1373.790 ;
        RECT 2498.110 1373.410 2498.410 1374.470 ;
        RECT 2545.950 1374.090 2546.250 1374.470 ;
        RECT 2594.710 1374.470 2642.850 1374.770 ;
        RECT 2545.950 1373.790 2594.090 1374.090 ;
        RECT 2497.190 1373.110 2498.410 1373.410 ;
        RECT 2593.790 1373.410 2594.090 1373.790 ;
        RECT 2594.710 1373.410 2595.010 1374.470 ;
        RECT 2642.550 1374.090 2642.850 1374.470 ;
        RECT 2691.310 1374.470 2739.450 1374.770 ;
        RECT 2642.550 1373.790 2690.690 1374.090 ;
        RECT 2593.790 1373.110 2595.010 1373.410 ;
        RECT 2690.390 1373.410 2690.690 1373.790 ;
        RECT 2691.310 1373.410 2691.610 1374.470 ;
        RECT 2739.150 1374.090 2739.450 1374.470 ;
        RECT 2787.910 1374.470 2836.050 1374.770 ;
        RECT 2739.150 1373.790 2787.290 1374.090 ;
        RECT 2690.390 1373.110 2691.610 1373.410 ;
        RECT 2786.990 1373.410 2787.290 1373.790 ;
        RECT 2787.910 1373.410 2788.210 1374.470 ;
        RECT 2835.750 1374.090 2836.050 1374.470 ;
        RECT 2916.710 1374.090 2917.010 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 2835.750 1373.790 2883.890 1374.090 ;
        RECT 2786.990 1373.110 2788.210 1373.410 ;
        RECT 2883.590 1373.410 2883.890 1373.790 ;
        RECT 2884.510 1373.790 2917.010 1374.090 ;
        RECT 2884.510 1373.410 2884.810 1373.790 ;
        RECT 2883.590 1373.110 2884.810 1373.410 ;
        RECT 2052.585 1373.095 2052.915 1373.110 ;
        RECT 1895.265 1371.750 1931.690 1372.050 ;
        RECT 1895.265 1371.735 1895.595 1371.750 ;
      LAYER via3 ;
        RECT 1261.620 2497.820 1261.940 2498.140 ;
        RECT 1980.140 1375.820 1980.460 1376.140 ;
        RECT 1386.740 1375.140 1387.060 1375.460 ;
        RECT 1331.540 1374.460 1331.860 1374.780 ;
        RECT 1441.940 1374.460 1442.260 1374.780 ;
        RECT 1261.620 1373.780 1261.940 1374.100 ;
        RECT 1386.740 1373.780 1387.060 1374.100 ;
        RECT 1980.140 1374.460 1980.460 1374.780 ;
        RECT 1331.540 1373.100 1331.860 1373.420 ;
        RECT 1441.940 1373.100 1442.260 1373.420 ;
      LAYER met4 ;
        RECT 1261.615 2497.815 1261.945 2498.145 ;
        RECT 1261.630 1374.105 1261.930 2497.815 ;
        RECT 1980.135 1375.815 1980.465 1376.145 ;
        RECT 1386.735 1375.135 1387.065 1375.465 ;
        RECT 1331.535 1374.455 1331.865 1374.785 ;
        RECT 1261.615 1373.775 1261.945 1374.105 ;
        RECT 1331.550 1373.425 1331.850 1374.455 ;
        RECT 1386.750 1374.105 1387.050 1375.135 ;
        RECT 1980.150 1374.785 1980.450 1375.815 ;
        RECT 1441.935 1374.455 1442.265 1374.785 ;
        RECT 1980.135 1374.455 1980.465 1374.785 ;
        RECT 1386.735 1373.775 1387.065 1374.105 ;
        RECT 1441.950 1373.425 1442.250 1374.455 ;
        RECT 1331.535 1373.095 1331.865 1373.425 ;
        RECT 1441.935 1373.095 1442.265 1373.425 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2090.310 1608.780 2090.630 1608.840 ;
        RECT 2124.810 1608.780 2125.130 1608.840 ;
        RECT 2090.310 1608.640 2125.130 1608.780 ;
        RECT 2090.310 1608.580 2090.630 1608.640 ;
        RECT 2124.810 1608.580 2125.130 1608.640 ;
        RECT 1825.810 1608.440 1826.130 1608.500 ;
        RECT 1881.930 1608.440 1882.250 1608.500 ;
        RECT 1825.810 1608.300 1882.250 1608.440 ;
        RECT 1825.810 1608.240 1826.130 1608.300 ;
        RECT 1881.930 1608.240 1882.250 1608.300 ;
        RECT 1895.270 1608.440 1895.590 1608.500 ;
        RECT 1973.010 1608.440 1973.330 1608.500 ;
        RECT 1895.270 1608.300 1973.330 1608.440 ;
        RECT 1895.270 1608.240 1895.590 1608.300 ;
        RECT 1973.010 1608.240 1973.330 1608.300 ;
      LAYER via ;
        RECT 2090.340 1608.580 2090.600 1608.840 ;
        RECT 2124.840 1608.580 2125.100 1608.840 ;
        RECT 1825.840 1608.240 1826.100 1608.500 ;
        RECT 1881.960 1608.240 1882.220 1608.500 ;
        RECT 1895.300 1608.240 1895.560 1608.500 ;
        RECT 1973.040 1608.240 1973.300 1608.500 ;
      LAYER met2 ;
        RECT 1278.890 2498.050 1279.170 2500.000 ;
        RECT 1280.270 2498.050 1280.550 2498.165 ;
        RECT 1278.890 2497.910 1280.550 2498.050 ;
        RECT 1278.890 2496.000 1279.170 2497.910 ;
        RECT 1280.270 2497.795 1280.550 2497.910 ;
        RECT 2052.610 1609.715 2052.890 1610.085 ;
        RECT 1606.410 1609.035 1606.690 1609.405 ;
        RECT 1606.480 1608.045 1606.620 1609.035 ;
        RECT 1883.330 1608.610 1883.610 1608.725 ;
        RECT 1882.020 1608.530 1883.610 1608.610 ;
        RECT 1825.840 1608.210 1826.100 1608.530 ;
        RECT 1881.960 1608.470 1883.610 1608.530 ;
        RECT 1881.960 1608.210 1882.220 1608.470 ;
        RECT 1883.330 1608.355 1883.610 1608.470 ;
        RECT 1895.290 1608.355 1895.570 1608.725 ;
        RECT 1994.650 1608.610 1994.930 1608.725 ;
        RECT 1895.300 1608.210 1895.560 1608.355 ;
        RECT 1973.040 1608.210 1973.300 1608.530 ;
        RECT 1993.800 1608.470 1994.930 1608.610 ;
        RECT 1606.410 1607.675 1606.690 1608.045 ;
        RECT 1642.290 1607.675 1642.570 1608.045 ;
        RECT 1738.890 1607.675 1739.170 1608.045 ;
        RECT 1642.360 1606.685 1642.500 1607.675 ;
        RECT 1738.960 1606.685 1739.100 1607.675 ;
        RECT 1825.900 1607.365 1826.040 1608.210 ;
        RECT 1973.100 1608.045 1973.240 1608.210 ;
        RECT 1993.800 1608.045 1993.940 1608.470 ;
        RECT 1994.650 1608.355 1994.930 1608.470 ;
        RECT 2052.680 1608.045 2052.820 1609.715 ;
        RECT 2124.830 1609.035 2125.110 1609.405 ;
        RECT 2124.900 1608.870 2125.040 1609.035 ;
        RECT 2090.340 1608.725 2090.600 1608.870 ;
        RECT 2090.330 1608.355 2090.610 1608.725 ;
        RECT 2124.840 1608.550 2125.100 1608.870 ;
        RECT 1973.030 1607.675 1973.310 1608.045 ;
        RECT 1993.730 1607.675 1994.010 1608.045 ;
        RECT 2052.610 1607.675 2052.890 1608.045 ;
        RECT 1825.830 1606.995 1826.110 1607.365 ;
        RECT 1642.290 1606.315 1642.570 1606.685 ;
        RECT 1687.830 1606.315 1688.110 1606.685 ;
        RECT 1738.890 1606.315 1739.170 1606.685 ;
        RECT 1687.900 1605.325 1688.040 1606.315 ;
        RECT 1687.830 1604.955 1688.110 1605.325 ;
      LAYER via2 ;
        RECT 1280.270 2497.840 1280.550 2498.120 ;
        RECT 2052.610 1609.760 2052.890 1610.040 ;
        RECT 1606.410 1609.080 1606.690 1609.360 ;
        RECT 1883.330 1608.400 1883.610 1608.680 ;
        RECT 1895.290 1608.400 1895.570 1608.680 ;
        RECT 1606.410 1607.720 1606.690 1608.000 ;
        RECT 1642.290 1607.720 1642.570 1608.000 ;
        RECT 1738.890 1607.720 1739.170 1608.000 ;
        RECT 1994.650 1608.400 1994.930 1608.680 ;
        RECT 2124.830 1609.080 2125.110 1609.360 ;
        RECT 2090.330 1608.400 2090.610 1608.680 ;
        RECT 1973.030 1607.720 1973.310 1608.000 ;
        RECT 1993.730 1607.720 1994.010 1608.000 ;
        RECT 2052.610 1607.720 2052.890 1608.000 ;
        RECT 1825.830 1607.040 1826.110 1607.320 ;
        RECT 1642.290 1606.360 1642.570 1606.640 ;
        RECT 1687.830 1606.360 1688.110 1606.640 ;
        RECT 1738.890 1606.360 1739.170 1606.640 ;
        RECT 1687.830 1605.000 1688.110 1605.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1612.700 2924.800 1613.900 ;
=======
        RECT 1280.245 2498.130 1280.575 2498.145 ;
        RECT 1280.910 2498.130 1281.290 2498.140 ;
        RECT 1280.245 2497.830 1281.290 2498.130 ;
        RECT 1280.245 2497.815 1280.575 2497.830 ;
        RECT 1280.910 2497.820 1281.290 2497.830 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2916.710 1613.150 2924.800 1613.450 ;
        RECT 2052.585 1610.050 2052.915 1610.065 ;
        RECT 1352.710 1609.750 1376.930 1610.050 ;
        RECT 1280.910 1609.370 1281.290 1609.380 ;
        RECT 1352.710 1609.370 1353.010 1609.750 ;
        RECT 1280.910 1609.070 1353.010 1609.370 ;
        RECT 1376.630 1609.370 1376.930 1609.750 ;
        RECT 2028.910 1609.750 2052.915 1610.050 ;
        RECT 1400.510 1609.370 1400.890 1609.380 ;
        RECT 1376.630 1609.070 1400.890 1609.370 ;
        RECT 1280.910 1609.060 1281.290 1609.070 ;
        RECT 1400.510 1609.060 1400.890 1609.070 ;
        RECT 1441.910 1609.370 1442.290 1609.380 ;
        RECT 1606.385 1609.370 1606.715 1609.385 ;
        RECT 1441.910 1609.070 1521.370 1609.370 ;
        RECT 1441.910 1609.060 1442.290 1609.070 ;
        RECT 1521.070 1608.690 1521.370 1609.070 ;
        RECT 1545.910 1609.070 1606.715 1609.370 ;
        RECT 1545.910 1608.690 1546.210 1609.070 ;
        RECT 1606.385 1609.055 1606.715 1609.070 ;
        RECT 1521.070 1608.390 1546.210 1608.690 ;
        RECT 1883.305 1608.690 1883.635 1608.705 ;
        RECT 1895.265 1608.690 1895.595 1608.705 ;
        RECT 1883.305 1608.390 1895.595 1608.690 ;
        RECT 1883.305 1608.375 1883.635 1608.390 ;
        RECT 1895.265 1608.375 1895.595 1608.390 ;
        RECT 1994.625 1608.690 1994.955 1608.705 ;
        RECT 2028.910 1608.690 2029.210 1609.750 ;
        RECT 2052.585 1609.735 2052.915 1609.750 ;
        RECT 2124.805 1609.370 2125.135 1609.385 ;
        RECT 2124.805 1609.070 2159.850 1609.370 ;
        RECT 2124.805 1609.055 2125.135 1609.070 ;
        RECT 2090.305 1608.690 2090.635 1608.705 ;
        RECT 1994.625 1608.390 2029.210 1608.690 ;
        RECT 2076.750 1608.390 2090.635 1608.690 ;
        RECT 2159.550 1608.690 2159.850 1609.070 ;
        RECT 2208.310 1609.070 2256.450 1609.370 ;
        RECT 2159.550 1608.390 2207.690 1608.690 ;
        RECT 1994.625 1608.375 1994.955 1608.390 ;
        RECT 1400.510 1608.010 1400.890 1608.020 ;
        RECT 1441.910 1608.010 1442.290 1608.020 ;
        RECT 1400.510 1607.710 1442.290 1608.010 ;
        RECT 1400.510 1607.700 1400.890 1607.710 ;
        RECT 1441.910 1607.700 1442.290 1607.710 ;
        RECT 1606.385 1608.010 1606.715 1608.025 ;
        RECT 1642.265 1608.010 1642.595 1608.025 ;
        RECT 1606.385 1607.710 1642.595 1608.010 ;
        RECT 1606.385 1607.695 1606.715 1607.710 ;
        RECT 1642.265 1607.695 1642.595 1607.710 ;
        RECT 1730.790 1608.010 1731.170 1608.020 ;
        RECT 1738.865 1608.010 1739.195 1608.025 ;
        RECT 1730.790 1607.710 1739.195 1608.010 ;
        RECT 1730.790 1607.700 1731.170 1607.710 ;
        RECT 1738.865 1607.695 1739.195 1607.710 ;
        RECT 1973.005 1608.010 1973.335 1608.025 ;
        RECT 1993.705 1608.010 1994.035 1608.025 ;
        RECT 1973.005 1607.710 1994.035 1608.010 ;
        RECT 1973.005 1607.695 1973.335 1607.710 ;
        RECT 1993.705 1607.695 1994.035 1607.710 ;
        RECT 2052.585 1608.010 2052.915 1608.025 ;
        RECT 2076.750 1608.010 2077.050 1608.390 ;
        RECT 2090.305 1608.375 2090.635 1608.390 ;
        RECT 2052.585 1607.710 2077.050 1608.010 ;
        RECT 2207.390 1608.010 2207.690 1608.390 ;
        RECT 2208.310 1608.010 2208.610 1609.070 ;
        RECT 2256.150 1608.690 2256.450 1609.070 ;
        RECT 2304.910 1609.070 2353.050 1609.370 ;
        RECT 2256.150 1608.390 2304.290 1608.690 ;
        RECT 2207.390 1607.710 2208.610 1608.010 ;
        RECT 2303.990 1608.010 2304.290 1608.390 ;
        RECT 2304.910 1608.010 2305.210 1609.070 ;
        RECT 2352.750 1608.690 2353.050 1609.070 ;
        RECT 2401.510 1609.070 2449.650 1609.370 ;
        RECT 2352.750 1608.390 2400.890 1608.690 ;
        RECT 2303.990 1607.710 2305.210 1608.010 ;
        RECT 2400.590 1608.010 2400.890 1608.390 ;
        RECT 2401.510 1608.010 2401.810 1609.070 ;
        RECT 2449.350 1608.690 2449.650 1609.070 ;
        RECT 2498.110 1609.070 2546.250 1609.370 ;
        RECT 2449.350 1608.390 2497.490 1608.690 ;
        RECT 2400.590 1607.710 2401.810 1608.010 ;
        RECT 2497.190 1608.010 2497.490 1608.390 ;
        RECT 2498.110 1608.010 2498.410 1609.070 ;
        RECT 2545.950 1608.690 2546.250 1609.070 ;
        RECT 2594.710 1609.070 2642.850 1609.370 ;
        RECT 2545.950 1608.390 2594.090 1608.690 ;
        RECT 2497.190 1607.710 2498.410 1608.010 ;
        RECT 2593.790 1608.010 2594.090 1608.390 ;
        RECT 2594.710 1608.010 2595.010 1609.070 ;
        RECT 2642.550 1608.690 2642.850 1609.070 ;
        RECT 2691.310 1609.070 2739.450 1609.370 ;
        RECT 2642.550 1608.390 2690.690 1608.690 ;
        RECT 2593.790 1607.710 2595.010 1608.010 ;
        RECT 2690.390 1608.010 2690.690 1608.390 ;
        RECT 2691.310 1608.010 2691.610 1609.070 ;
        RECT 2739.150 1608.690 2739.450 1609.070 ;
        RECT 2787.910 1609.070 2836.050 1609.370 ;
        RECT 2739.150 1608.390 2787.290 1608.690 ;
        RECT 2690.390 1607.710 2691.610 1608.010 ;
        RECT 2786.990 1608.010 2787.290 1608.390 ;
        RECT 2787.910 1608.010 2788.210 1609.070 ;
        RECT 2835.750 1608.690 2836.050 1609.070 ;
        RECT 2916.710 1608.690 2917.010 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 2835.750 1608.390 2883.890 1608.690 ;
        RECT 2786.990 1607.710 2788.210 1608.010 ;
        RECT 2883.590 1608.010 2883.890 1608.390 ;
        RECT 2884.510 1608.390 2917.010 1608.690 ;
        RECT 2884.510 1608.010 2884.810 1608.390 ;
        RECT 2883.590 1607.710 2884.810 1608.010 ;
        RECT 2052.585 1607.695 2052.915 1607.710 ;
        RECT 1825.805 1607.330 1826.135 1607.345 ;
        RECT 1785.110 1607.030 1826.135 1607.330 ;
        RECT 1642.265 1606.650 1642.595 1606.665 ;
        RECT 1687.805 1606.650 1688.135 1606.665 ;
        RECT 1642.265 1606.350 1688.135 1606.650 ;
        RECT 1642.265 1606.335 1642.595 1606.350 ;
        RECT 1687.805 1606.335 1688.135 1606.350 ;
        RECT 1738.865 1606.650 1739.195 1606.665 ;
        RECT 1785.110 1606.650 1785.410 1607.030 ;
        RECT 1825.805 1607.015 1826.135 1607.030 ;
        RECT 1738.865 1606.350 1785.410 1606.650 ;
        RECT 1738.865 1606.335 1739.195 1606.350 ;
        RECT 1687.805 1605.290 1688.135 1605.305 ;
        RECT 1730.790 1605.290 1731.170 1605.300 ;
        RECT 1687.805 1604.990 1731.170 1605.290 ;
        RECT 1687.805 1604.975 1688.135 1604.990 ;
        RECT 1730.790 1604.980 1731.170 1604.990 ;
      LAYER via3 ;
        RECT 1280.940 2497.820 1281.260 2498.140 ;
        RECT 1280.940 1609.060 1281.260 1609.380 ;
        RECT 1400.540 1609.060 1400.860 1609.380 ;
        RECT 1441.940 1609.060 1442.260 1609.380 ;
        RECT 1400.540 1607.700 1400.860 1608.020 ;
        RECT 1441.940 1607.700 1442.260 1608.020 ;
        RECT 1730.820 1607.700 1731.140 1608.020 ;
        RECT 1730.820 1604.980 1731.140 1605.300 ;
      LAYER met4 ;
        RECT 1280.935 2497.815 1281.265 2498.145 ;
        RECT 1280.950 1609.385 1281.250 2497.815 ;
        RECT 1280.935 1609.055 1281.265 1609.385 ;
        RECT 1400.535 1609.055 1400.865 1609.385 ;
        RECT 1441.935 1609.055 1442.265 1609.385 ;
        RECT 1400.550 1608.025 1400.850 1609.055 ;
        RECT 1441.950 1608.025 1442.250 1609.055 ;
        RECT 1400.535 1607.695 1400.865 1608.025 ;
        RECT 1441.935 1607.695 1442.265 1608.025 ;
        RECT 1730.815 1607.695 1731.145 1608.025 ;
        RECT 1730.830 1605.305 1731.130 1607.695 ;
        RECT 1730.815 1604.975 1731.145 1605.305 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1298.650 2514.200 1298.970 2514.260 ;
        RECT 1949.550 2514.200 1949.870 2514.260 ;
        RECT 1298.650 2514.060 1949.870 2514.200 ;
        RECT 1298.650 2514.000 1298.970 2514.060 ;
        RECT 1949.550 2514.000 1949.870 2514.060 ;
        RECT 1949.550 1849.160 1949.870 1849.220 ;
        RECT 2900.830 1849.160 2901.150 1849.220 ;
        RECT 1949.550 1849.020 2901.150 1849.160 ;
        RECT 1949.550 1848.960 1949.870 1849.020 ;
        RECT 2900.830 1848.960 2901.150 1849.020 ;
      LAYER via ;
        RECT 1298.680 2514.000 1298.940 2514.260 ;
        RECT 1949.580 2514.000 1949.840 2514.260 ;
        RECT 1949.580 1848.960 1949.840 1849.220 ;
        RECT 2900.860 1848.960 2901.120 1849.220 ;
      LAYER met2 ;
        RECT 1298.680 2513.970 1298.940 2514.290 ;
        RECT 1949.580 2513.970 1949.840 2514.290 ;
        RECT 1298.740 2500.000 1298.880 2513.970 ;
        RECT 1298.670 2496.000 1298.950 2500.000 ;
        RECT 1949.640 1849.250 1949.780 2513.970 ;
        RECT 1949.580 1848.930 1949.840 1849.250 ;
        RECT 2900.860 1848.930 2901.120 1849.250 ;
        RECT 2900.920 1848.085 2901.060 1848.930 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1847.300 2924.800 1848.500 ;
=======
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1318.430 2515.900 1318.750 2515.960 ;
        RECT 1950.930 2515.900 1951.250 2515.960 ;
        RECT 1318.430 2515.760 1951.250 2515.900 ;
        RECT 1318.430 2515.700 1318.750 2515.760 ;
        RECT 1950.930 2515.700 1951.250 2515.760 ;
        RECT 1950.930 2083.760 1951.250 2083.820 ;
        RECT 2900.830 2083.760 2901.150 2083.820 ;
        RECT 1950.930 2083.620 2901.150 2083.760 ;
        RECT 1950.930 2083.560 1951.250 2083.620 ;
        RECT 2900.830 2083.560 2901.150 2083.620 ;
      LAYER via ;
        RECT 1318.460 2515.700 1318.720 2515.960 ;
        RECT 1950.960 2515.700 1951.220 2515.960 ;
        RECT 1950.960 2083.560 1951.220 2083.820 ;
        RECT 2900.860 2083.560 2901.120 2083.820 ;
      LAYER met2 ;
        RECT 1318.460 2515.670 1318.720 2515.990 ;
        RECT 1950.960 2515.670 1951.220 2515.990 ;
        RECT 1318.520 2500.000 1318.660 2515.670 ;
        RECT 1318.450 2496.000 1318.730 2500.000 ;
        RECT 1951.020 2083.850 1951.160 2515.670 ;
        RECT 1950.960 2083.530 1951.220 2083.850 ;
        RECT 2900.860 2083.530 2901.120 2083.850 ;
        RECT 2900.920 2082.685 2901.060 2083.530 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2081.900 2924.800 2083.100 ;
=======
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1338.210 2516.920 1338.530 2516.980 ;
        RECT 1948.630 2516.920 1948.950 2516.980 ;
        RECT 1338.210 2516.780 1948.950 2516.920 ;
        RECT 1338.210 2516.720 1338.530 2516.780 ;
        RECT 1948.630 2516.720 1948.950 2516.780 ;
        RECT 1948.630 2318.360 1948.950 2318.420 ;
        RECT 2900.830 2318.360 2901.150 2318.420 ;
        RECT 1948.630 2318.220 2901.150 2318.360 ;
        RECT 1948.630 2318.160 1948.950 2318.220 ;
        RECT 2900.830 2318.160 2901.150 2318.220 ;
      LAYER via ;
        RECT 1338.240 2516.720 1338.500 2516.980 ;
        RECT 1948.660 2516.720 1948.920 2516.980 ;
        RECT 1948.660 2318.160 1948.920 2318.420 ;
        RECT 2900.860 2318.160 2901.120 2318.420 ;
      LAYER met2 ;
        RECT 1338.240 2516.690 1338.500 2517.010 ;
        RECT 1948.660 2516.690 1948.920 2517.010 ;
        RECT 1338.300 2500.000 1338.440 2516.690 ;
        RECT 1338.230 2496.000 1338.510 2500.000 ;
        RECT 1948.720 2318.450 1948.860 2516.690 ;
        RECT 1948.660 2318.130 1948.920 2318.450 ;
        RECT 2900.860 2318.130 2901.120 2318.450 ;
        RECT 2900.920 2317.285 2901.060 2318.130 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2316.500 2924.800 2317.700 ;
=======
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1200.670 146.780 1200.990 146.840 ;
        RECT 1265.990 146.780 1266.310 146.840 ;
        RECT 1200.670 146.640 1266.310 146.780 ;
        RECT 1200.670 146.580 1200.990 146.640 ;
        RECT 1265.990 146.580 1266.310 146.640 ;
        RECT 2090.310 146.100 2090.630 146.160 ;
        RECT 2124.810 146.100 2125.130 146.160 ;
        RECT 2090.310 145.960 2125.130 146.100 ;
        RECT 2090.310 145.900 2090.630 145.960 ;
        RECT 2124.810 145.900 2125.130 145.960 ;
        RECT 1344.650 145.760 1344.970 145.820 ;
        RECT 1386.510 145.760 1386.830 145.820 ;
        RECT 1344.650 145.620 1386.830 145.760 ;
        RECT 1344.650 145.560 1344.970 145.620 ;
        RECT 1386.510 145.560 1386.830 145.620 ;
        RECT 1895.270 145.420 1895.590 145.480 ;
        RECT 1930.230 145.420 1930.550 145.480 ;
        RECT 1895.270 145.280 1930.550 145.420 ;
        RECT 1895.270 145.220 1895.590 145.280 ;
        RECT 1930.230 145.220 1930.550 145.280 ;
        RECT 1932.070 145.420 1932.390 145.480 ;
        RECT 1956.450 145.420 1956.770 145.480 ;
        RECT 1932.070 145.280 1956.770 145.420 ;
        RECT 1932.070 145.220 1932.390 145.280 ;
        RECT 1956.450 145.220 1956.770 145.280 ;
        RECT 2042.010 145.080 2042.330 145.140 ;
        RECT 2069.610 145.080 2069.930 145.140 ;
        RECT 2042.010 144.940 2069.930 145.080 ;
        RECT 2042.010 144.880 2042.330 144.940 ;
        RECT 2069.610 144.880 2069.930 144.940 ;
      LAYER via ;
        RECT 1200.700 146.580 1200.960 146.840 ;
        RECT 1266.020 146.580 1266.280 146.840 ;
        RECT 2090.340 145.900 2090.600 146.160 ;
        RECT 2124.840 145.900 2125.100 146.160 ;
        RECT 1344.680 145.560 1344.940 145.820 ;
        RECT 1386.540 145.560 1386.800 145.820 ;
        RECT 1895.300 145.220 1895.560 145.480 ;
        RECT 1930.260 145.220 1930.520 145.480 ;
        RECT 1932.100 145.220 1932.360 145.480 ;
        RECT 1956.480 145.220 1956.740 145.480 ;
        RECT 2042.040 144.880 2042.300 145.140 ;
        RECT 2069.640 144.880 2069.900 145.140 ;
      LAYER met2 ;
        RECT 1166.190 2498.050 1166.470 2500.000 ;
        RECT 1168.030 2498.050 1168.310 2498.165 ;
        RECT 1166.190 2497.910 1168.310 2498.050 ;
        RECT 1166.190 2496.000 1166.470 2497.910 ;
        RECT 1168.030 2497.795 1168.310 2497.910 ;
        RECT 1318.910 149.075 1319.190 149.445 ;
        RECT 1266.010 147.715 1266.290 148.085 ;
        RECT 1266.080 146.870 1266.220 147.715 ;
        RECT 1200.700 146.725 1200.960 146.870 ;
        RECT 1200.690 146.355 1200.970 146.725 ;
        RECT 1266.020 146.550 1266.280 146.870 ;
        RECT 1318.980 146.725 1319.120 149.075 ;
        RECT 1318.910 146.355 1319.190 146.725 ;
        RECT 1344.670 146.355 1344.950 146.725 ;
        RECT 1956.470 146.355 1956.750 146.725 ;
        RECT 1993.730 146.355 1994.010 146.725 ;
        RECT 2124.830 146.355 2125.110 146.725 ;
        RECT 1344.740 145.850 1344.880 146.355 ;
        RECT 1344.680 145.530 1344.940 145.850 ;
        RECT 1386.540 145.530 1386.800 145.850 ;
        RECT 1895.290 145.675 1895.570 146.045 ;
        RECT 1386.600 145.365 1386.740 145.530 ;
        RECT 1895.360 145.510 1895.500 145.675 ;
        RECT 1386.530 144.995 1386.810 145.365 ;
        RECT 1895.300 145.190 1895.560 145.510 ;
        RECT 1930.250 145.165 1930.530 145.535 ;
        RECT 1956.540 145.510 1956.680 146.355 ;
        RECT 1993.800 145.930 1993.940 146.355 ;
        RECT 2124.900 146.190 2125.040 146.355 ;
        RECT 2090.340 146.045 2090.600 146.190 ;
        RECT 1994.650 145.930 1994.930 146.045 ;
        RECT 1993.800 145.790 1994.930 145.930 ;
        RECT 1994.650 145.675 1994.930 145.790 ;
        RECT 2090.330 145.675 2090.610 146.045 ;
        RECT 2124.840 145.870 2125.100 146.190 ;
        RECT 1932.100 145.365 1932.360 145.510 ;
        RECT 1932.090 144.995 1932.370 145.365 ;
        RECT 1956.480 145.190 1956.740 145.510 ;
        RECT 2042.030 144.995 2042.310 145.365 ;
        RECT 2069.630 144.995 2069.910 145.365 ;
        RECT 2042.040 144.850 2042.300 144.995 ;
        RECT 2069.640 144.850 2069.900 144.995 ;
      LAYER via2 ;
        RECT 1168.030 2497.840 1168.310 2498.120 ;
        RECT 1318.910 149.120 1319.190 149.400 ;
        RECT 1266.010 147.760 1266.290 148.040 ;
        RECT 1200.690 146.400 1200.970 146.680 ;
        RECT 1318.910 146.400 1319.190 146.680 ;
        RECT 1344.670 146.400 1344.950 146.680 ;
        RECT 1956.470 146.400 1956.750 146.680 ;
        RECT 1993.730 146.400 1994.010 146.680 ;
        RECT 2124.830 146.400 2125.110 146.680 ;
        RECT 1895.290 145.720 1895.570 146.000 ;
        RECT 1386.530 145.040 1386.810 145.320 ;
        RECT 1994.650 145.720 1994.930 146.000 ;
        RECT 2090.330 145.720 2090.610 146.000 ;
        RECT 1930.250 145.210 1930.530 145.490 ;
        RECT 1932.090 145.040 1932.370 145.320 ;
        RECT 2042.030 145.040 2042.310 145.320 ;
        RECT 2069.630 145.040 2069.910 145.320 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 145.940 2924.800 147.140 ;
=======
        RECT 1168.005 2498.130 1168.335 2498.145 ;
        RECT 1169.590 2498.130 1169.970 2498.140 ;
        RECT 1168.005 2497.830 1169.970 2498.130 ;
        RECT 1168.005 2497.815 1168.335 2497.830 ;
        RECT 1169.590 2497.820 1169.970 2497.830 ;
        RECT 1290.110 149.410 1290.490 149.420 ;
        RECT 1318.885 149.410 1319.215 149.425 ;
        RECT 1290.110 149.110 1319.215 149.410 ;
        RECT 1290.110 149.100 1290.490 149.110 ;
        RECT 1318.885 149.095 1319.215 149.110 ;
        RECT 1447.470 148.430 1483.650 148.730 ;
        RECT 1169.590 148.050 1169.970 148.060 ;
        RECT 1265.985 148.050 1266.315 148.065 ;
        RECT 1290.110 148.050 1290.490 148.060 ;
        RECT 1169.590 147.750 1200.290 148.050 ;
        RECT 1169.590 147.740 1169.970 147.750 ;
        RECT 1199.990 146.690 1200.290 147.750 ;
        RECT 1265.985 147.750 1290.490 148.050 ;
        RECT 1265.985 147.735 1266.315 147.750 ;
        RECT 1290.110 147.740 1290.490 147.750 ;
        RECT 1200.665 146.690 1200.995 146.705 ;
        RECT 1199.990 146.390 1200.995 146.690 ;
        RECT 1200.665 146.375 1200.995 146.390 ;
        RECT 1318.885 146.690 1319.215 146.705 ;
        RECT 1344.645 146.690 1344.975 146.705 ;
        RECT 1447.470 146.690 1447.770 148.430 ;
        RECT 1483.350 148.050 1483.650 148.430 ;
        RECT 1483.350 147.750 1531.490 148.050 ;
        RECT 1531.190 147.370 1531.490 147.750 ;
        RECT 1702.310 147.750 1738.490 148.050 ;
        RECT 1531.190 147.070 1545.290 147.370 ;
        RECT 1318.885 146.390 1344.975 146.690 ;
        RECT 1318.885 146.375 1319.215 146.390 ;
        RECT 1344.645 146.375 1344.975 146.390 ;
        RECT 1394.110 146.390 1447.770 146.690 ;
        RECT 1394.110 146.010 1394.410 146.390 ;
        RECT 1393.190 145.710 1394.410 146.010 ;
        RECT 1544.990 146.010 1545.290 147.070 ;
        RECT 1617.670 146.390 1641.890 146.690 ;
        RECT 1617.670 146.010 1617.970 146.390 ;
        RECT 1544.990 145.710 1617.970 146.010 ;
        RECT 1386.505 145.330 1386.835 145.345 ;
        RECT 1393.190 145.330 1393.490 145.710 ;
        RECT 1386.505 145.030 1393.490 145.330 ;
        RECT 1641.590 145.330 1641.890 146.390 ;
        RECT 1702.310 146.010 1702.610 147.750 ;
        RECT 1738.190 147.380 1738.490 147.750 ;
        RECT 1798.910 147.750 1835.090 148.050 ;
        RECT 1738.150 147.060 1738.530 147.380 ;
        RECT 1798.910 146.010 1799.210 147.750 ;
        RECT 1834.790 147.380 1835.090 147.750 ;
        RECT 1834.750 147.060 1835.130 147.380 ;
        RECT 1956.445 146.690 1956.775 146.705 ;
        RECT 1993.705 146.690 1994.035 146.705 ;
        RECT 1956.445 146.390 1994.035 146.690 ;
        RECT 1956.445 146.375 1956.775 146.390 ;
        RECT 1993.705 146.375 1994.035 146.390 ;
        RECT 2124.805 146.690 2125.135 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2124.805 146.390 2159.850 146.690 ;
        RECT 2124.805 146.375 2125.135 146.390 ;
        RECT 1895.265 146.010 1895.595 146.025 ;
        RECT 1656.310 145.710 1702.610 146.010 ;
        RECT 1752.910 145.710 1799.210 146.010 ;
        RECT 1849.510 145.710 1895.595 146.010 ;
        RECT 1656.310 145.330 1656.610 145.710 ;
        RECT 1641.590 145.030 1656.610 145.330 ;
        RECT 1738.150 145.330 1738.530 145.340 ;
        RECT 1752.910 145.330 1753.210 145.710 ;
        RECT 1738.150 145.030 1753.210 145.330 ;
        RECT 1834.750 145.330 1835.130 145.340 ;
        RECT 1849.510 145.330 1849.810 145.710 ;
        RECT 1895.265 145.695 1895.595 145.710 ;
        RECT 1994.625 146.010 1994.955 146.025 ;
        RECT 2090.305 146.010 2090.635 146.025 ;
        RECT 1994.625 145.710 2021.850 146.010 ;
        RECT 1994.625 145.695 1994.955 145.710 ;
        RECT 1834.750 145.030 1849.810 145.330 ;
        RECT 1930.225 145.500 1930.555 145.515 ;
        RECT 1930.225 145.330 1931.690 145.500 ;
        RECT 1932.065 145.330 1932.395 145.345 ;
        RECT 1930.225 145.200 1932.395 145.330 ;
        RECT 1930.225 145.185 1930.555 145.200 ;
        RECT 1931.390 145.030 1932.395 145.200 ;
        RECT 2021.550 145.330 2021.850 145.710 ;
        RECT 2076.750 145.710 2090.635 146.010 ;
        RECT 2159.550 146.010 2159.850 146.390 ;
        RECT 2208.310 146.390 2256.450 146.690 ;
        RECT 2159.550 145.710 2207.690 146.010 ;
        RECT 2042.005 145.330 2042.335 145.345 ;
        RECT 2021.550 145.030 2042.335 145.330 ;
        RECT 1386.505 145.015 1386.835 145.030 ;
        RECT 1738.150 145.020 1738.530 145.030 ;
        RECT 1834.750 145.020 1835.130 145.030 ;
        RECT 1932.065 145.015 1932.395 145.030 ;
        RECT 2042.005 145.015 2042.335 145.030 ;
        RECT 2069.605 145.330 2069.935 145.345 ;
        RECT 2076.750 145.330 2077.050 145.710 ;
        RECT 2090.305 145.695 2090.635 145.710 ;
        RECT 2069.605 145.030 2077.050 145.330 ;
        RECT 2207.390 145.330 2207.690 145.710 ;
        RECT 2208.310 145.330 2208.610 146.390 ;
        RECT 2256.150 146.010 2256.450 146.390 ;
        RECT 2304.910 146.390 2353.050 146.690 ;
        RECT 2256.150 145.710 2304.290 146.010 ;
        RECT 2207.390 145.030 2208.610 145.330 ;
        RECT 2303.990 145.330 2304.290 145.710 ;
        RECT 2304.910 145.330 2305.210 146.390 ;
        RECT 2352.750 146.010 2353.050 146.390 ;
        RECT 2401.510 146.390 2449.650 146.690 ;
        RECT 2352.750 145.710 2400.890 146.010 ;
        RECT 2303.990 145.030 2305.210 145.330 ;
        RECT 2400.590 145.330 2400.890 145.710 ;
        RECT 2401.510 145.330 2401.810 146.390 ;
        RECT 2449.350 146.010 2449.650 146.390 ;
        RECT 2498.110 146.390 2546.250 146.690 ;
        RECT 2449.350 145.710 2497.490 146.010 ;
        RECT 2400.590 145.030 2401.810 145.330 ;
        RECT 2497.190 145.330 2497.490 145.710 ;
        RECT 2498.110 145.330 2498.410 146.390 ;
        RECT 2545.950 146.010 2546.250 146.390 ;
        RECT 2594.710 146.390 2642.850 146.690 ;
        RECT 2545.950 145.710 2594.090 146.010 ;
        RECT 2497.190 145.030 2498.410 145.330 ;
        RECT 2593.790 145.330 2594.090 145.710 ;
        RECT 2594.710 145.330 2595.010 146.390 ;
        RECT 2642.550 146.010 2642.850 146.390 ;
        RECT 2691.310 146.390 2739.450 146.690 ;
        RECT 2642.550 145.710 2690.690 146.010 ;
        RECT 2593.790 145.030 2595.010 145.330 ;
        RECT 2690.390 145.330 2690.690 145.710 ;
        RECT 2691.310 145.330 2691.610 146.390 ;
        RECT 2739.150 146.010 2739.450 146.390 ;
        RECT 2787.910 146.390 2836.050 146.690 ;
        RECT 2739.150 145.710 2787.290 146.010 ;
        RECT 2690.390 145.030 2691.610 145.330 ;
        RECT 2786.990 145.330 2787.290 145.710 ;
        RECT 2787.910 145.330 2788.210 146.390 ;
        RECT 2835.750 146.010 2836.050 146.390 ;
        RECT 2916.710 146.390 2924.800 146.690 ;
        RECT 2916.710 146.010 2917.010 146.390 ;
        RECT 2835.750 145.710 2883.890 146.010 ;
        RECT 2786.990 145.030 2788.210 145.330 ;
        RECT 2883.590 145.330 2883.890 145.710 ;
        RECT 2884.510 145.710 2917.010 146.010 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT 2884.510 145.330 2884.810 145.710 ;
        RECT 2883.590 145.030 2884.810 145.330 ;
        RECT 2069.605 145.015 2069.935 145.030 ;
      LAYER via3 ;
        RECT 1169.620 2497.820 1169.940 2498.140 ;
        RECT 1290.140 149.100 1290.460 149.420 ;
        RECT 1169.620 147.740 1169.940 148.060 ;
        RECT 1290.140 147.740 1290.460 148.060 ;
        RECT 1738.180 147.060 1738.500 147.380 ;
        RECT 1834.780 147.060 1835.100 147.380 ;
        RECT 1738.180 145.020 1738.500 145.340 ;
        RECT 1834.780 145.020 1835.100 145.340 ;
      LAYER met4 ;
        RECT 1169.615 2497.815 1169.945 2498.145 ;
        RECT 1169.630 148.065 1169.930 2497.815 ;
        RECT 1290.135 149.095 1290.465 149.425 ;
        RECT 1290.150 148.065 1290.450 149.095 ;
        RECT 1169.615 147.735 1169.945 148.065 ;
        RECT 1290.135 147.735 1290.465 148.065 ;
        RECT 1738.175 147.055 1738.505 147.385 ;
        RECT 1834.775 147.055 1835.105 147.385 ;
        RECT 1738.190 145.345 1738.490 147.055 ;
        RECT 1834.790 145.345 1835.090 147.055 ;
        RECT 1738.175 145.015 1738.505 145.345 ;
        RECT 1834.775 145.015 1835.105 145.345 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1365.885 2496.025 1366.055 2497.215 ;
      LAYER mcon ;
        RECT 1365.885 2497.045 1366.055 2497.215 ;
      LAYER met1 ;
        RECT 1365.810 2497.200 1366.130 2497.260 ;
        RECT 1365.615 2497.060 1366.130 2497.200 ;
        RECT 1365.810 2497.000 1366.130 2497.060 ;
        RECT 1365.825 2496.180 1366.115 2496.225 ;
        RECT 2900.830 2496.180 2901.150 2496.240 ;
        RECT 1365.825 2496.040 2901.150 2496.180 ;
        RECT 1365.825 2495.995 1366.115 2496.040 ;
        RECT 2900.830 2495.980 2901.150 2496.040 ;
      LAYER via ;
        RECT 1365.840 2497.000 1366.100 2497.260 ;
        RECT 2900.860 2495.980 2901.120 2496.240 ;
      LAYER met2 ;
        RECT 1364.450 2497.370 1364.730 2500.000 ;
        RECT 1364.450 2497.290 1366.040 2497.370 ;
        RECT 1364.450 2497.230 1366.100 2497.290 ;
        RECT 1364.450 2496.000 1364.730 2497.230 ;
        RECT 1365.840 2496.970 1366.100 2497.230 ;
        RECT 2900.860 2495.950 2901.120 2496.270 ;
        RECT 2900.920 2493.405 2901.060 2495.950 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2492.620 2924.800 2493.820 ;
=======
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1386.510 2725.680 1386.830 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 1386.510 2725.540 2901.150 2725.680 ;
        RECT 1386.510 2725.480 1386.830 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
      LAYER via ;
        RECT 1386.540 2725.480 1386.800 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 1386.540 2725.450 1386.800 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 1384.690 2499.410 1384.970 2500.000 ;
        RECT 1386.600 2499.410 1386.740 2725.450 ;
        RECT 1384.690 2499.270 1386.740 2499.410 ;
        RECT 1384.690 2496.000 1384.970 2499.270 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2727.220 2924.800 2728.420 ;
=======
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1407.210 2960.280 1407.530 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 1407.210 2960.140 2901.150 2960.280 ;
        RECT 1407.210 2960.080 1407.530 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 1407.240 2960.080 1407.500 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 1407.240 2960.050 1407.500 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 1404.470 2498.730 1404.750 2500.000 ;
        RECT 1407.300 2498.730 1407.440 2960.050 ;
        RECT 1404.470 2498.590 1407.440 2498.730 ;
        RECT 1404.470 2496.000 1404.750 2498.590 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2961.820 2924.800 2963.020 ;
=======
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1427.910 3195.220 1428.230 3195.280 ;
        RECT 2900.830 3195.220 2901.150 3195.280 ;
        RECT 1427.910 3195.080 2901.150 3195.220 ;
        RECT 1427.910 3195.020 1428.230 3195.080 ;
        RECT 2900.830 3195.020 2901.150 3195.080 ;
        RECT 1424.230 2514.880 1424.550 2514.940 ;
        RECT 1427.910 2514.880 1428.230 2514.940 ;
        RECT 1424.230 2514.740 1428.230 2514.880 ;
        RECT 1424.230 2514.680 1424.550 2514.740 ;
        RECT 1427.910 2514.680 1428.230 2514.740 ;
      LAYER via ;
        RECT 1427.940 3195.020 1428.200 3195.280 ;
        RECT 2900.860 3195.020 2901.120 3195.280 ;
        RECT 1424.260 2514.680 1424.520 2514.940 ;
        RECT 1427.940 2514.680 1428.200 2514.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3195.310 2901.060 3196.835 ;
        RECT 1427.940 3194.990 1428.200 3195.310 ;
        RECT 2900.860 3194.990 2901.120 3195.310 ;
        RECT 1428.000 2514.970 1428.140 3194.990 ;
        RECT 1424.260 2514.650 1424.520 2514.970 ;
        RECT 1427.940 2514.650 1428.200 2514.970 ;
        RECT 1424.320 2500.000 1424.460 2514.650 ;
        RECT 1424.250 2496.000 1424.530 2500.000 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3196.420 2924.800 3197.620 ;
=======
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2028.760 3429.680 2065.700 3429.820 ;
        RECT 1448.610 3429.480 1448.930 3429.540 ;
        RECT 2028.760 3429.480 2028.900 3429.680 ;
        RECT 1448.610 3429.340 2028.900 3429.480 ;
        RECT 2065.560 3429.480 2065.700 3429.680 ;
        RECT 2146.060 3429.680 2149.880 3429.820 ;
        RECT 2146.060 3429.480 2146.200 3429.680 ;
        RECT 2065.560 3429.340 2146.200 3429.480 ;
        RECT 2149.740 3429.480 2149.880 3429.680 ;
        RECT 2704.960 3429.680 2714.300 3429.820 ;
        RECT 2704.960 3429.480 2705.100 3429.680 ;
        RECT 2149.740 3429.340 2705.100 3429.480 ;
        RECT 2714.160 3429.480 2714.300 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2714.160 3429.340 2901.150 3429.480 ;
        RECT 1448.610 3429.280 1448.930 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
        RECT 1444.010 2514.880 1444.330 2514.940 ;
        RECT 1448.610 2514.880 1448.930 2514.940 ;
        RECT 1444.010 2514.740 1448.930 2514.880 ;
        RECT 1444.010 2514.680 1444.330 2514.740 ;
        RECT 1448.610 2514.680 1448.930 2514.740 ;
      LAYER via ;
        RECT 1448.640 3429.280 1448.900 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
        RECT 1444.040 2514.680 1444.300 2514.940 ;
        RECT 1448.640 2514.680 1448.900 2514.940 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1448.640 3429.250 1448.900 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1448.700 2514.970 1448.840 3429.250 ;
        RECT 1444.040 2514.650 1444.300 2514.970 ;
        RECT 1448.640 2514.650 1448.900 2514.970 ;
        RECT 1444.100 2500.000 1444.240 2514.650 ;
        RECT 1444.030 2496.000 1444.310 2500.000 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3431.020 2924.800 3432.220 ;
=======
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2713.685 3332.765 2713.855 3422.355 ;
        RECT 2713.225 3139.645 2713.395 3187.755 ;
        RECT 2712.765 3088.645 2712.935 3132.675 ;
        RECT 2713.685 2946.525 2713.855 3035.775 ;
        RECT 2712.305 2753.065 2712.475 2801.175 ;
      LAYER mcon ;
        RECT 2713.685 3422.185 2713.855 3422.355 ;
        RECT 2713.225 3187.585 2713.395 3187.755 ;
        RECT 2712.765 3132.505 2712.935 3132.675 ;
        RECT 2713.685 3035.605 2713.855 3035.775 ;
        RECT 2712.305 2801.005 2712.475 2801.175 ;
      LAYER met1 ;
        RECT 2713.610 3491.360 2713.930 3491.420 ;
        RECT 2717.750 3491.360 2718.070 3491.420 ;
        RECT 2713.610 3491.220 2718.070 3491.360 ;
        RECT 2713.610 3491.160 2713.930 3491.220 ;
        RECT 2717.750 3491.160 2718.070 3491.220 ;
        RECT 2713.610 3443.220 2713.930 3443.480 ;
        RECT 2712.690 3443.080 2713.010 3443.140 ;
        RECT 2713.700 3443.080 2713.840 3443.220 ;
        RECT 2712.690 3442.940 2713.840 3443.080 ;
        RECT 2712.690 3442.880 2713.010 3442.940 ;
        RECT 2712.230 3422.340 2712.550 3422.400 ;
        RECT 2713.625 3422.340 2713.915 3422.385 ;
        RECT 2712.230 3422.200 2713.915 3422.340 ;
        RECT 2712.230 3422.140 2712.550 3422.200 ;
        RECT 2713.625 3422.155 2713.915 3422.200 ;
        RECT 2713.625 3332.920 2713.915 3332.965 ;
        RECT 2714.070 3332.920 2714.390 3332.980 ;
        RECT 2713.625 3332.780 2714.390 3332.920 ;
        RECT 2713.625 3332.735 2713.915 3332.780 ;
        RECT 2714.070 3332.720 2714.390 3332.780 ;
        RECT 2712.690 3236.360 2713.010 3236.420 ;
        RECT 2713.150 3236.360 2713.470 3236.420 ;
        RECT 2712.690 3236.220 2713.470 3236.360 ;
        RECT 2712.690 3236.160 2713.010 3236.220 ;
        RECT 2713.150 3236.160 2713.470 3236.220 ;
        RECT 2713.150 3187.740 2713.470 3187.800 ;
        RECT 2712.955 3187.600 2713.470 3187.740 ;
        RECT 2713.150 3187.540 2713.470 3187.600 ;
        RECT 2713.165 3139.800 2713.455 3139.845 ;
        RECT 2713.610 3139.800 2713.930 3139.860 ;
        RECT 2713.165 3139.660 2713.930 3139.800 ;
        RECT 2713.165 3139.615 2713.455 3139.660 ;
        RECT 2713.610 3139.600 2713.930 3139.660 ;
        RECT 2712.705 3132.660 2712.995 3132.705 ;
        RECT 2713.610 3132.660 2713.930 3132.720 ;
        RECT 2712.705 3132.520 2713.930 3132.660 ;
        RECT 2712.705 3132.475 2712.995 3132.520 ;
        RECT 2713.610 3132.460 2713.930 3132.520 ;
        RECT 2712.690 3088.800 2713.010 3088.860 ;
        RECT 2712.495 3088.660 2713.010 3088.800 ;
        RECT 2712.690 3088.600 2713.010 3088.660 ;
        RECT 2713.150 3036.440 2713.470 3036.500 ;
        RECT 2713.610 3036.440 2713.930 3036.500 ;
        RECT 2713.150 3036.300 2713.930 3036.440 ;
        RECT 2713.150 3036.240 2713.470 3036.300 ;
        RECT 2713.610 3036.240 2713.930 3036.300 ;
        RECT 2713.610 3035.760 2713.930 3035.820 ;
        RECT 2713.415 3035.620 2713.930 3035.760 ;
        RECT 2713.610 3035.560 2713.930 3035.620 ;
        RECT 2713.625 2946.680 2713.915 2946.725 ;
        RECT 2714.070 2946.680 2714.390 2946.740 ;
        RECT 2713.625 2946.540 2714.390 2946.680 ;
        RECT 2713.625 2946.495 2713.915 2946.540 ;
        RECT 2714.070 2946.480 2714.390 2946.540 ;
        RECT 2714.070 2912.340 2714.390 2912.400 ;
        RECT 2713.700 2912.200 2714.390 2912.340 ;
        RECT 2713.700 2911.720 2713.840 2912.200 ;
        RECT 2714.070 2912.140 2714.390 2912.200 ;
        RECT 2713.610 2911.460 2713.930 2911.720 ;
        RECT 2712.230 2815.580 2712.550 2815.840 ;
        RECT 2712.320 2815.160 2712.460 2815.580 ;
        RECT 2712.230 2814.900 2712.550 2815.160 ;
        RECT 2712.230 2801.160 2712.550 2801.220 ;
        RECT 2712.035 2801.020 2712.550 2801.160 ;
        RECT 2712.230 2800.960 2712.550 2801.020 ;
        RECT 2712.245 2753.220 2712.535 2753.265 ;
        RECT 2713.150 2753.220 2713.470 2753.280 ;
        RECT 2712.245 2753.080 2713.470 2753.220 ;
        RECT 2712.245 2753.035 2712.535 2753.080 ;
        RECT 2713.150 2753.020 2713.470 2753.080 ;
        RECT 2712.230 2718.200 2712.550 2718.260 ;
        RECT 2713.150 2718.200 2713.470 2718.260 ;
        RECT 2712.230 2718.060 2713.470 2718.200 ;
        RECT 2712.230 2718.000 2712.550 2718.060 ;
        RECT 2713.150 2718.000 2713.470 2718.060 ;
        RECT 2712.230 2670.260 2712.550 2670.320 ;
        RECT 2713.150 2670.260 2713.470 2670.320 ;
        RECT 2712.230 2670.120 2713.470 2670.260 ;
        RECT 2712.230 2670.060 2712.550 2670.120 ;
        RECT 2713.150 2670.060 2713.470 2670.120 ;
        RECT 2713.150 2622.120 2713.470 2622.380 ;
        RECT 2713.240 2621.980 2713.380 2622.120 ;
        RECT 2713.610 2621.980 2713.930 2622.040 ;
        RECT 2713.240 2621.840 2713.930 2621.980 ;
        RECT 2713.610 2621.780 2713.930 2621.840 ;
        RECT 2712.690 2560.100 2713.010 2560.160 ;
        RECT 2714.070 2560.100 2714.390 2560.160 ;
        RECT 2712.690 2559.960 2714.390 2560.100 ;
        RECT 2712.690 2559.900 2713.010 2559.960 ;
        RECT 2714.070 2559.900 2714.390 2559.960 ;
        RECT 1463.790 2515.220 1464.110 2515.280 ;
        RECT 1463.790 2515.080 1483.800 2515.220 ;
        RECT 1463.790 2515.020 1464.110 2515.080 ;
        RECT 1483.660 2514.880 1483.800 2515.080 ;
        RECT 2714.070 2514.880 2714.390 2514.940 ;
        RECT 1483.660 2514.740 2714.390 2514.880 ;
        RECT 2714.070 2514.680 2714.390 2514.740 ;
      LAYER via ;
        RECT 2713.640 3491.160 2713.900 3491.420 ;
        RECT 2717.780 3491.160 2718.040 3491.420 ;
        RECT 2713.640 3443.220 2713.900 3443.480 ;
        RECT 2712.720 3442.880 2712.980 3443.140 ;
        RECT 2712.260 3422.140 2712.520 3422.400 ;
        RECT 2714.100 3332.720 2714.360 3332.980 ;
        RECT 2712.720 3236.160 2712.980 3236.420 ;
        RECT 2713.180 3236.160 2713.440 3236.420 ;
        RECT 2713.180 3187.540 2713.440 3187.800 ;
        RECT 2713.640 3139.600 2713.900 3139.860 ;
        RECT 2713.640 3132.460 2713.900 3132.720 ;
        RECT 2712.720 3088.600 2712.980 3088.860 ;
        RECT 2713.180 3036.240 2713.440 3036.500 ;
        RECT 2713.640 3036.240 2713.900 3036.500 ;
        RECT 2713.640 3035.560 2713.900 3035.820 ;
        RECT 2714.100 2946.480 2714.360 2946.740 ;
        RECT 2714.100 2912.140 2714.360 2912.400 ;
        RECT 2713.640 2911.460 2713.900 2911.720 ;
        RECT 2712.260 2815.580 2712.520 2815.840 ;
        RECT 2712.260 2814.900 2712.520 2815.160 ;
        RECT 2712.260 2800.960 2712.520 2801.220 ;
        RECT 2713.180 2753.020 2713.440 2753.280 ;
        RECT 2712.260 2718.000 2712.520 2718.260 ;
        RECT 2713.180 2718.000 2713.440 2718.260 ;
        RECT 2712.260 2670.060 2712.520 2670.320 ;
        RECT 2713.180 2670.060 2713.440 2670.320 ;
        RECT 2713.180 2622.120 2713.440 2622.380 ;
        RECT 2713.640 2621.780 2713.900 2622.040 ;
        RECT 2712.720 2559.900 2712.980 2560.160 ;
        RECT 2714.100 2559.900 2714.360 2560.160 ;
        RECT 1463.820 2515.020 1464.080 2515.280 ;
        RECT 2714.100 2514.680 2714.360 2514.940 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2717.170 3519.700 2717.730 3524.800 ;
=======
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3517.370 2717.520 3517.600 ;
        RECT 2717.380 3517.230 2717.980 3517.370 ;
        RECT 2717.840 3491.450 2717.980 3517.230 ;
        RECT 2713.640 3491.130 2713.900 3491.450 ;
        RECT 2717.780 3491.130 2718.040 3491.450 ;
        RECT 2713.700 3443.510 2713.840 3491.130 ;
        RECT 2713.640 3443.190 2713.900 3443.510 ;
        RECT 2712.720 3442.850 2712.980 3443.170 ;
        RECT 2712.780 3429.650 2712.920 3442.850 ;
        RECT 2712.320 3429.510 2712.920 3429.650 ;
        RECT 2712.320 3422.430 2712.460 3429.510 ;
        RECT 2712.260 3422.110 2712.520 3422.430 ;
        RECT 2714.100 3332.690 2714.360 3333.010 ;
        RECT 2714.160 3298.410 2714.300 3332.690 ;
        RECT 2713.240 3298.270 2714.300 3298.410 ;
        RECT 2713.240 3236.450 2713.380 3298.270 ;
        RECT 2712.720 3236.130 2712.980 3236.450 ;
        RECT 2713.180 3236.130 2713.440 3236.450 ;
        RECT 2712.780 3201.850 2712.920 3236.130 ;
        RECT 2712.780 3201.710 2713.380 3201.850 ;
        RECT 2713.240 3187.830 2713.380 3201.710 ;
        RECT 2713.180 3187.510 2713.440 3187.830 ;
        RECT 2713.640 3139.570 2713.900 3139.890 ;
        RECT 2713.700 3132.750 2713.840 3139.570 ;
        RECT 2713.640 3132.430 2713.900 3132.750 ;
        RECT 2712.720 3088.570 2712.980 3088.890 ;
        RECT 2712.780 3084.325 2712.920 3088.570 ;
        RECT 2712.710 3083.955 2712.990 3084.325 ;
        RECT 2713.630 3083.955 2713.910 3084.325 ;
        RECT 2713.700 3036.530 2713.840 3083.955 ;
        RECT 2713.180 3036.210 2713.440 3036.530 ;
        RECT 2713.640 3036.210 2713.900 3036.530 ;
        RECT 2713.240 3035.930 2713.380 3036.210 ;
        RECT 2713.240 3035.850 2713.840 3035.930 ;
        RECT 2713.240 3035.790 2713.900 3035.850 ;
        RECT 2713.640 3035.530 2713.900 3035.790 ;
        RECT 2714.100 2946.450 2714.360 2946.770 ;
        RECT 2714.160 2912.430 2714.300 2946.450 ;
        RECT 2714.100 2912.110 2714.360 2912.430 ;
        RECT 2713.640 2911.430 2713.900 2911.750 ;
        RECT 2713.700 2863.210 2713.840 2911.430 ;
        RECT 2712.780 2863.070 2713.840 2863.210 ;
        RECT 2712.780 2849.610 2712.920 2863.070 ;
        RECT 2712.320 2849.470 2712.920 2849.610 ;
        RECT 2712.320 2815.870 2712.460 2849.470 ;
        RECT 2712.260 2815.550 2712.520 2815.870 ;
        RECT 2712.260 2814.870 2712.520 2815.190 ;
        RECT 2712.320 2801.250 2712.460 2814.870 ;
        RECT 2712.260 2800.930 2712.520 2801.250 ;
        RECT 2713.180 2752.990 2713.440 2753.310 ;
        RECT 2713.240 2718.290 2713.380 2752.990 ;
        RECT 2712.260 2717.970 2712.520 2718.290 ;
        RECT 2713.180 2717.970 2713.440 2718.290 ;
        RECT 2712.320 2670.350 2712.460 2717.970 ;
        RECT 2712.260 2670.030 2712.520 2670.350 ;
        RECT 2713.180 2670.030 2713.440 2670.350 ;
        RECT 2713.240 2622.410 2713.380 2670.030 ;
        RECT 2713.180 2622.090 2713.440 2622.410 ;
        RECT 2713.640 2621.750 2713.900 2622.070 ;
        RECT 2713.700 2608.325 2713.840 2621.750 ;
        RECT 2712.710 2607.955 2712.990 2608.325 ;
        RECT 2713.630 2607.955 2713.910 2608.325 ;
        RECT 2712.780 2560.190 2712.920 2607.955 ;
        RECT 2712.720 2559.870 2712.980 2560.190 ;
        RECT 2714.100 2559.870 2714.360 2560.190 ;
        RECT 1463.820 2514.990 1464.080 2515.310 ;
        RECT 1463.880 2500.000 1464.020 2514.990 ;
        RECT 2714.160 2514.970 2714.300 2559.870 ;
        RECT 2714.100 2514.650 2714.360 2514.970 ;
        RECT 1463.810 2496.000 1464.090 2500.000 ;
      LAYER via2 ;
        RECT 2712.710 3084.000 2712.990 3084.280 ;
        RECT 2713.630 3084.000 2713.910 3084.280 ;
        RECT 2712.710 2608.000 2712.990 2608.280 ;
        RECT 2713.630 2608.000 2713.910 2608.280 ;
      LAYER met3 ;
        RECT 2712.685 3084.290 2713.015 3084.305 ;
        RECT 2713.605 3084.290 2713.935 3084.305 ;
        RECT 2712.685 3083.990 2713.935 3084.290 ;
        RECT 2712.685 3083.975 2713.015 3083.990 ;
        RECT 2713.605 3083.975 2713.935 3083.990 ;
        RECT 2712.685 2608.290 2713.015 2608.305 ;
        RECT 2713.605 2608.290 2713.935 2608.305 ;
        RECT 2712.685 2607.990 2713.935 2608.290 ;
        RECT 2712.685 2607.975 2713.015 2607.990 ;
        RECT 2713.605 2607.975 2713.935 2607.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2387.545 3332.765 2387.715 3380.875 ;
        RECT 2388.005 2815.285 2388.175 2849.455 ;
      LAYER mcon ;
        RECT 2387.545 3380.705 2387.715 3380.875 ;
        RECT 2388.005 2849.285 2388.175 2849.455 ;
      LAYER met1 ;
        RECT 2387.470 3380.860 2387.790 3380.920 ;
        RECT 2387.275 3380.720 2387.790 3380.860 ;
        RECT 2387.470 3380.660 2387.790 3380.720 ;
        RECT 2387.485 3332.920 2387.775 3332.965 ;
        RECT 2387.930 3332.920 2388.250 3332.980 ;
        RECT 2387.485 3332.780 2388.250 3332.920 ;
        RECT 2387.485 3332.735 2387.775 3332.780 ;
        RECT 2387.930 3332.720 2388.250 3332.780 ;
        RECT 2387.470 3270.700 2387.790 3270.760 ;
        RECT 2388.390 3270.700 2388.710 3270.760 ;
        RECT 2387.470 3270.560 2388.710 3270.700 ;
        RECT 2387.470 3270.500 2387.790 3270.560 ;
        RECT 2388.390 3270.500 2388.710 3270.560 ;
        RECT 2387.470 3174.140 2387.790 3174.200 ;
        RECT 2388.390 3174.140 2388.710 3174.200 ;
        RECT 2387.470 3174.000 2388.710 3174.140 ;
        RECT 2387.470 3173.940 2387.790 3174.000 ;
        RECT 2388.390 3173.940 2388.710 3174.000 ;
        RECT 2387.470 3077.580 2387.790 3077.640 ;
        RECT 2388.390 3077.580 2388.710 3077.640 ;
        RECT 2387.470 3077.440 2388.710 3077.580 ;
        RECT 2387.470 3077.380 2387.790 3077.440 ;
        RECT 2388.390 3077.380 2388.710 3077.440 ;
        RECT 2387.470 2981.020 2387.790 2981.080 ;
        RECT 2388.390 2981.020 2388.710 2981.080 ;
        RECT 2387.470 2980.880 2388.710 2981.020 ;
        RECT 2387.470 2980.820 2387.790 2980.880 ;
        RECT 2388.390 2980.820 2388.710 2980.880 ;
        RECT 2386.550 2946.340 2386.870 2946.400 ;
        RECT 2387.930 2946.340 2388.250 2946.400 ;
        RECT 2386.550 2946.200 2388.250 2946.340 ;
        RECT 2386.550 2946.140 2386.870 2946.200 ;
        RECT 2387.930 2946.140 2388.250 2946.200 ;
        RECT 2387.930 2849.440 2388.250 2849.500 ;
        RECT 2387.735 2849.300 2388.250 2849.440 ;
        RECT 2387.930 2849.240 2388.250 2849.300 ;
        RECT 2387.945 2815.440 2388.235 2815.485 ;
        RECT 2388.850 2815.440 2389.170 2815.500 ;
        RECT 2387.945 2815.300 2389.170 2815.440 ;
        RECT 2387.945 2815.255 2388.235 2815.300 ;
        RECT 2388.850 2815.240 2389.170 2815.300 ;
        RECT 2387.930 2753.220 2388.250 2753.280 ;
        RECT 2389.310 2753.220 2389.630 2753.280 ;
        RECT 2387.930 2753.080 2389.630 2753.220 ;
        RECT 2387.930 2753.020 2388.250 2753.080 ;
        RECT 2389.310 2753.020 2389.630 2753.080 ;
        RECT 2389.310 2719.220 2389.630 2719.280 ;
        RECT 2388.940 2719.080 2389.630 2719.220 ;
        RECT 2388.940 2718.600 2389.080 2719.080 ;
        RECT 2389.310 2719.020 2389.630 2719.080 ;
        RECT 2388.850 2718.340 2389.170 2718.600 ;
        RECT 2388.850 2670.400 2389.170 2670.660 ;
        RECT 2388.940 2669.920 2389.080 2670.400 ;
        RECT 2389.310 2669.920 2389.630 2669.980 ;
        RECT 2388.940 2669.780 2389.630 2669.920 ;
        RECT 2389.310 2669.720 2389.630 2669.780 ;
        RECT 2389.310 2649.520 2389.630 2649.580 ;
        RECT 2390.230 2649.520 2390.550 2649.580 ;
        RECT 2389.310 2649.380 2390.550 2649.520 ;
        RECT 2389.310 2649.320 2389.630 2649.380 ;
        RECT 2390.230 2649.320 2390.550 2649.380 ;
        RECT 2389.310 2573.360 2389.630 2573.420 ;
        RECT 2390.230 2573.360 2390.550 2573.420 ;
        RECT 2389.310 2573.220 2390.550 2573.360 ;
        RECT 2389.310 2573.160 2389.630 2573.220 ;
        RECT 2390.230 2573.160 2390.550 2573.220 ;
        RECT 1485.410 2515.220 1485.730 2515.280 ;
        RECT 2389.310 2515.220 2389.630 2515.280 ;
        RECT 1485.410 2515.080 2389.630 2515.220 ;
        RECT 1485.410 2515.020 1485.730 2515.080 ;
        RECT 2389.310 2515.020 2389.630 2515.080 ;
      LAYER via ;
        RECT 2387.500 3380.660 2387.760 3380.920 ;
        RECT 2387.960 3332.720 2388.220 3332.980 ;
        RECT 2387.500 3270.500 2387.760 3270.760 ;
        RECT 2388.420 3270.500 2388.680 3270.760 ;
        RECT 2387.500 3173.940 2387.760 3174.200 ;
        RECT 2388.420 3173.940 2388.680 3174.200 ;
        RECT 2387.500 3077.380 2387.760 3077.640 ;
        RECT 2388.420 3077.380 2388.680 3077.640 ;
        RECT 2387.500 2980.820 2387.760 2981.080 ;
        RECT 2388.420 2980.820 2388.680 2981.080 ;
        RECT 2386.580 2946.140 2386.840 2946.400 ;
        RECT 2387.960 2946.140 2388.220 2946.400 ;
        RECT 2387.960 2849.240 2388.220 2849.500 ;
        RECT 2388.880 2815.240 2389.140 2815.500 ;
        RECT 2387.960 2753.020 2388.220 2753.280 ;
        RECT 2389.340 2753.020 2389.600 2753.280 ;
        RECT 2389.340 2719.020 2389.600 2719.280 ;
        RECT 2388.880 2718.340 2389.140 2718.600 ;
        RECT 2388.880 2670.400 2389.140 2670.660 ;
        RECT 2389.340 2669.720 2389.600 2669.980 ;
        RECT 2389.340 2649.320 2389.600 2649.580 ;
        RECT 2390.260 2649.320 2390.520 2649.580 ;
        RECT 2389.340 2573.160 2389.600 2573.420 ;
        RECT 2390.260 2573.160 2390.520 2573.420 ;
        RECT 1485.440 2515.020 1485.700 2515.280 ;
        RECT 2389.340 2515.020 2389.600 2515.280 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2392.410 3519.700 2392.970 3524.800 ;
=======
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3517.370 2392.760 3517.600 ;
        RECT 2392.620 3517.230 2393.220 3517.370 ;
        RECT 2393.080 3430.445 2393.220 3517.230 ;
        RECT 2393.010 3430.075 2393.290 3430.445 ;
        RECT 2388.410 3429.395 2388.690 3429.765 ;
        RECT 2388.480 3394.970 2388.620 3429.395 ;
        RECT 2387.560 3394.830 2388.620 3394.970 ;
        RECT 2387.560 3380.950 2387.700 3394.830 ;
        RECT 2387.500 3380.630 2387.760 3380.950 ;
        RECT 2387.960 3332.690 2388.220 3333.010 ;
        RECT 2388.020 3298.410 2388.160 3332.690 ;
        RECT 2388.020 3298.270 2388.620 3298.410 ;
        RECT 2388.480 3270.790 2388.620 3298.270 ;
        RECT 2387.500 3270.470 2387.760 3270.790 ;
        RECT 2388.420 3270.470 2388.680 3270.790 ;
        RECT 2387.560 3222.250 2387.700 3270.470 ;
        RECT 2387.560 3222.110 2388.620 3222.250 ;
        RECT 2388.480 3174.230 2388.620 3222.110 ;
        RECT 2387.500 3173.910 2387.760 3174.230 ;
        RECT 2388.420 3173.910 2388.680 3174.230 ;
        RECT 2387.560 3125.690 2387.700 3173.910 ;
        RECT 2387.560 3125.550 2388.620 3125.690 ;
        RECT 2388.480 3077.670 2388.620 3125.550 ;
        RECT 2387.500 3077.350 2387.760 3077.670 ;
        RECT 2388.420 3077.350 2388.680 3077.670 ;
        RECT 2387.560 3029.130 2387.700 3077.350 ;
        RECT 2387.560 3028.990 2388.620 3029.130 ;
        RECT 2388.480 2981.110 2388.620 3028.990 ;
        RECT 2387.500 2980.850 2387.760 2981.110 ;
        RECT 2387.500 2980.790 2388.160 2980.850 ;
        RECT 2388.420 2980.790 2388.680 2981.110 ;
        RECT 2387.560 2980.710 2388.160 2980.790 ;
        RECT 2388.020 2980.170 2388.160 2980.710 ;
        RECT 2388.020 2980.030 2388.620 2980.170 ;
        RECT 2388.480 2959.770 2388.620 2980.030 ;
        RECT 2388.020 2959.630 2388.620 2959.770 ;
        RECT 2388.020 2946.430 2388.160 2959.630 ;
        RECT 2386.580 2946.110 2386.840 2946.430 ;
        RECT 2387.960 2946.110 2388.220 2946.430 ;
        RECT 2386.640 2898.685 2386.780 2946.110 ;
        RECT 2386.570 2898.315 2386.850 2898.685 ;
        RECT 2387.490 2898.315 2387.770 2898.685 ;
        RECT 2387.560 2863.210 2387.700 2898.315 ;
        RECT 2387.560 2863.070 2388.160 2863.210 ;
        RECT 2388.020 2849.530 2388.160 2863.070 ;
        RECT 2387.960 2849.210 2388.220 2849.530 ;
        RECT 2388.880 2815.210 2389.140 2815.530 ;
        RECT 2388.940 2801.445 2389.080 2815.210 ;
        RECT 2387.950 2801.075 2388.230 2801.445 ;
        RECT 2388.870 2801.075 2389.150 2801.445 ;
        RECT 2388.020 2753.310 2388.160 2801.075 ;
        RECT 2387.960 2752.990 2388.220 2753.310 ;
        RECT 2389.340 2752.990 2389.600 2753.310 ;
        RECT 2389.400 2719.310 2389.540 2752.990 ;
        RECT 2389.340 2718.990 2389.600 2719.310 ;
        RECT 2388.880 2718.310 2389.140 2718.630 ;
        RECT 2388.940 2670.690 2389.080 2718.310 ;
        RECT 2388.880 2670.370 2389.140 2670.690 ;
        RECT 2389.340 2669.690 2389.600 2670.010 ;
        RECT 2389.400 2649.610 2389.540 2669.690 ;
        RECT 2389.340 2649.290 2389.600 2649.610 ;
        RECT 2390.260 2649.290 2390.520 2649.610 ;
        RECT 2390.320 2573.450 2390.460 2649.290 ;
        RECT 2389.340 2573.130 2389.600 2573.450 ;
        RECT 2390.260 2573.130 2390.520 2573.450 ;
        RECT 2389.400 2515.310 2389.540 2573.130 ;
        RECT 1485.440 2514.990 1485.700 2515.310 ;
        RECT 2389.340 2514.990 2389.600 2515.310 ;
        RECT 1483.590 2499.410 1483.870 2500.000 ;
        RECT 1485.500 2499.410 1485.640 2514.990 ;
        RECT 1483.590 2499.270 1485.640 2499.410 ;
        RECT 1483.590 2496.000 1483.870 2499.270 ;
      LAYER via2 ;
        RECT 2393.010 3430.120 2393.290 3430.400 ;
        RECT 2388.410 3429.440 2388.690 3429.720 ;
        RECT 2386.570 2898.360 2386.850 2898.640 ;
        RECT 2387.490 2898.360 2387.770 2898.640 ;
        RECT 2387.950 2801.120 2388.230 2801.400 ;
        RECT 2388.870 2801.120 2389.150 2801.400 ;
      LAYER met3 ;
        RECT 2392.985 3430.410 2393.315 3430.425 ;
        RECT 2387.710 3430.110 2393.315 3430.410 ;
        RECT 2387.710 3429.730 2388.010 3430.110 ;
        RECT 2392.985 3430.095 2393.315 3430.110 ;
        RECT 2388.385 3429.730 2388.715 3429.745 ;
        RECT 2387.710 3429.430 2388.715 3429.730 ;
        RECT 2388.385 3429.415 2388.715 3429.430 ;
        RECT 2386.545 2898.650 2386.875 2898.665 ;
        RECT 2387.465 2898.650 2387.795 2898.665 ;
        RECT 2386.545 2898.350 2387.795 2898.650 ;
        RECT 2386.545 2898.335 2386.875 2898.350 ;
        RECT 2387.465 2898.335 2387.795 2898.350 ;
        RECT 2387.925 2801.410 2388.255 2801.425 ;
        RECT 2388.845 2801.410 2389.175 2801.425 ;
        RECT 2387.925 2801.110 2389.175 2801.410 ;
        RECT 2387.925 2801.095 2388.255 2801.110 ;
        RECT 2388.845 2801.095 2389.175 2801.110 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2065.085 3332.765 2065.255 3422.355 ;
        RECT 2064.165 3008.405 2064.335 3042.915 ;
        RECT 2065.085 2946.525 2065.255 2994.635 ;
        RECT 2063.705 2753.065 2063.875 2801.175 ;
      LAYER mcon ;
        RECT 2065.085 3422.185 2065.255 3422.355 ;
        RECT 2064.165 3042.745 2064.335 3042.915 ;
        RECT 2065.085 2994.465 2065.255 2994.635 ;
        RECT 2063.705 2801.005 2063.875 2801.175 ;
      LAYER met1 ;
        RECT 2065.010 3491.360 2065.330 3491.420 ;
        RECT 2068.690 3491.360 2069.010 3491.420 ;
        RECT 2065.010 3491.220 2069.010 3491.360 ;
        RECT 2065.010 3491.160 2065.330 3491.220 ;
        RECT 2068.690 3491.160 2069.010 3491.220 ;
        RECT 2065.010 3443.220 2065.330 3443.480 ;
        RECT 2064.090 3443.080 2064.410 3443.140 ;
        RECT 2065.100 3443.080 2065.240 3443.220 ;
        RECT 2064.090 3442.940 2065.240 3443.080 ;
        RECT 2064.090 3442.880 2064.410 3442.940 ;
        RECT 2063.630 3422.340 2063.950 3422.400 ;
        RECT 2065.025 3422.340 2065.315 3422.385 ;
        RECT 2063.630 3422.200 2065.315 3422.340 ;
        RECT 2063.630 3422.140 2063.950 3422.200 ;
        RECT 2065.025 3422.155 2065.315 3422.200 ;
        RECT 2065.025 3332.920 2065.315 3332.965 ;
        RECT 2065.470 3332.920 2065.790 3332.980 ;
        RECT 2065.025 3332.780 2065.790 3332.920 ;
        RECT 2065.025 3332.735 2065.315 3332.780 ;
        RECT 2065.470 3332.720 2065.790 3332.780 ;
        RECT 2064.090 3236.360 2064.410 3236.420 ;
        RECT 2064.550 3236.360 2064.870 3236.420 ;
        RECT 2064.090 3236.220 2064.870 3236.360 ;
        RECT 2064.090 3236.160 2064.410 3236.220 ;
        RECT 2064.550 3236.160 2064.870 3236.220 ;
        RECT 2064.090 3202.020 2064.410 3202.080 ;
        RECT 2064.550 3202.020 2064.870 3202.080 ;
        RECT 2064.090 3201.880 2064.870 3202.020 ;
        RECT 2064.090 3201.820 2064.410 3201.880 ;
        RECT 2064.550 3201.820 2064.870 3201.880 ;
        RECT 2063.630 3153.400 2063.950 3153.460 ;
        RECT 2064.550 3153.400 2064.870 3153.460 ;
        RECT 2063.630 3153.260 2064.870 3153.400 ;
        RECT 2063.630 3153.200 2063.950 3153.260 ;
        RECT 2064.550 3153.200 2064.870 3153.260 ;
        RECT 2063.630 3056.840 2063.950 3056.900 ;
        RECT 2064.550 3056.840 2064.870 3056.900 ;
        RECT 2063.630 3056.700 2064.870 3056.840 ;
        RECT 2063.630 3056.640 2063.950 3056.700 ;
        RECT 2064.550 3056.640 2064.870 3056.700 ;
        RECT 2064.090 3042.900 2064.410 3042.960 ;
        RECT 2063.895 3042.760 2064.410 3042.900 ;
        RECT 2064.090 3042.700 2064.410 3042.760 ;
        RECT 2064.105 3008.560 2064.395 3008.605 ;
        RECT 2065.010 3008.560 2065.330 3008.620 ;
        RECT 2064.105 3008.420 2065.330 3008.560 ;
        RECT 2064.105 3008.375 2064.395 3008.420 ;
        RECT 2065.010 3008.360 2065.330 3008.420 ;
        RECT 2065.010 2994.620 2065.330 2994.680 ;
        RECT 2064.815 2994.480 2065.330 2994.620 ;
        RECT 2065.010 2994.420 2065.330 2994.480 ;
        RECT 2065.025 2946.680 2065.315 2946.725 ;
        RECT 2065.470 2946.680 2065.790 2946.740 ;
        RECT 2065.025 2946.540 2065.790 2946.680 ;
        RECT 2065.025 2946.495 2065.315 2946.540 ;
        RECT 2065.470 2946.480 2065.790 2946.540 ;
        RECT 2065.470 2912.340 2065.790 2912.400 ;
        RECT 2065.100 2912.200 2065.790 2912.340 ;
        RECT 2065.100 2911.720 2065.240 2912.200 ;
        RECT 2065.470 2912.140 2065.790 2912.200 ;
        RECT 2065.010 2911.460 2065.330 2911.720 ;
        RECT 2063.630 2815.580 2063.950 2815.840 ;
        RECT 2063.720 2815.160 2063.860 2815.580 ;
        RECT 2063.630 2814.900 2063.950 2815.160 ;
        RECT 2063.630 2801.160 2063.950 2801.220 ;
        RECT 2063.435 2801.020 2063.950 2801.160 ;
        RECT 2063.630 2800.960 2063.950 2801.020 ;
        RECT 2063.645 2753.220 2063.935 2753.265 ;
        RECT 2064.550 2753.220 2064.870 2753.280 ;
        RECT 2063.645 2753.080 2064.870 2753.220 ;
        RECT 2063.645 2753.035 2063.935 2753.080 ;
        RECT 2064.550 2753.020 2064.870 2753.080 ;
        RECT 2063.630 2718.200 2063.950 2718.260 ;
        RECT 2064.550 2718.200 2064.870 2718.260 ;
        RECT 2063.630 2718.060 2064.870 2718.200 ;
        RECT 2063.630 2718.000 2063.950 2718.060 ;
        RECT 2064.550 2718.000 2064.870 2718.060 ;
        RECT 2063.630 2670.260 2063.950 2670.320 ;
        RECT 2064.550 2670.260 2064.870 2670.320 ;
        RECT 2063.630 2670.120 2064.870 2670.260 ;
        RECT 2063.630 2670.060 2063.950 2670.120 ;
        RECT 2064.550 2670.060 2064.870 2670.120 ;
        RECT 2064.550 2622.120 2064.870 2622.380 ;
        RECT 2064.640 2621.980 2064.780 2622.120 ;
        RECT 2065.010 2621.980 2065.330 2622.040 ;
        RECT 2064.640 2621.840 2065.330 2621.980 ;
        RECT 2065.010 2621.780 2065.330 2621.840 ;
        RECT 2064.090 2560.100 2064.410 2560.160 ;
        RECT 2065.470 2560.100 2065.790 2560.160 ;
        RECT 2064.090 2559.960 2065.790 2560.100 ;
        RECT 2064.090 2559.900 2064.410 2559.960 ;
        RECT 2065.470 2559.900 2065.790 2559.960 ;
        RECT 1503.350 2517.940 1503.670 2518.000 ;
        RECT 1503.350 2517.800 1556.020 2517.940 ;
        RECT 1503.350 2517.740 1503.670 2517.800 ;
        RECT 1555.880 2517.600 1556.020 2517.800 ;
        RECT 2065.470 2517.600 2065.790 2517.660 ;
        RECT 1555.880 2517.460 2065.790 2517.600 ;
        RECT 2065.470 2517.400 2065.790 2517.460 ;
      LAYER via ;
        RECT 2065.040 3491.160 2065.300 3491.420 ;
        RECT 2068.720 3491.160 2068.980 3491.420 ;
        RECT 2065.040 3443.220 2065.300 3443.480 ;
        RECT 2064.120 3442.880 2064.380 3443.140 ;
        RECT 2063.660 3422.140 2063.920 3422.400 ;
        RECT 2065.500 3332.720 2065.760 3332.980 ;
        RECT 2064.120 3236.160 2064.380 3236.420 ;
        RECT 2064.580 3236.160 2064.840 3236.420 ;
        RECT 2064.120 3201.820 2064.380 3202.080 ;
        RECT 2064.580 3201.820 2064.840 3202.080 ;
        RECT 2063.660 3153.200 2063.920 3153.460 ;
        RECT 2064.580 3153.200 2064.840 3153.460 ;
        RECT 2063.660 3056.640 2063.920 3056.900 ;
        RECT 2064.580 3056.640 2064.840 3056.900 ;
        RECT 2064.120 3042.700 2064.380 3042.960 ;
        RECT 2065.040 3008.360 2065.300 3008.620 ;
        RECT 2065.040 2994.420 2065.300 2994.680 ;
        RECT 2065.500 2946.480 2065.760 2946.740 ;
        RECT 2065.500 2912.140 2065.760 2912.400 ;
        RECT 2065.040 2911.460 2065.300 2911.720 ;
        RECT 2063.660 2815.580 2063.920 2815.840 ;
        RECT 2063.660 2814.900 2063.920 2815.160 ;
        RECT 2063.660 2800.960 2063.920 2801.220 ;
        RECT 2064.580 2753.020 2064.840 2753.280 ;
        RECT 2063.660 2718.000 2063.920 2718.260 ;
        RECT 2064.580 2718.000 2064.840 2718.260 ;
        RECT 2063.660 2670.060 2063.920 2670.320 ;
        RECT 2064.580 2670.060 2064.840 2670.320 ;
        RECT 2064.580 2622.120 2064.840 2622.380 ;
        RECT 2065.040 2621.780 2065.300 2622.040 ;
        RECT 2064.120 2559.900 2064.380 2560.160 ;
        RECT 2065.500 2559.900 2065.760 2560.160 ;
        RECT 1503.380 2517.740 1503.640 2518.000 ;
        RECT 2065.500 2517.400 2065.760 2517.660 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2068.110 3519.700 2068.670 3524.800 ;
=======
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3517.370 2068.460 3517.600 ;
        RECT 2068.320 3517.230 2068.920 3517.370 ;
        RECT 2068.780 3491.450 2068.920 3517.230 ;
        RECT 2065.040 3491.130 2065.300 3491.450 ;
        RECT 2068.720 3491.130 2068.980 3491.450 ;
        RECT 2065.100 3443.510 2065.240 3491.130 ;
        RECT 2065.040 3443.190 2065.300 3443.510 ;
        RECT 2064.120 3442.850 2064.380 3443.170 ;
        RECT 2064.180 3429.650 2064.320 3442.850 ;
        RECT 2063.720 3429.510 2064.320 3429.650 ;
        RECT 2063.720 3422.430 2063.860 3429.510 ;
        RECT 2063.660 3422.110 2063.920 3422.430 ;
        RECT 2065.500 3332.690 2065.760 3333.010 ;
        RECT 2065.560 3298.410 2065.700 3332.690 ;
        RECT 2064.640 3298.270 2065.700 3298.410 ;
        RECT 2064.640 3236.450 2064.780 3298.270 ;
        RECT 2064.120 3236.130 2064.380 3236.450 ;
        RECT 2064.580 3236.130 2064.840 3236.450 ;
        RECT 2064.180 3202.110 2064.320 3236.130 ;
        RECT 2064.120 3201.790 2064.380 3202.110 ;
        RECT 2064.580 3201.790 2064.840 3202.110 ;
        RECT 2064.640 3153.490 2064.780 3201.790 ;
        RECT 2063.660 3153.170 2063.920 3153.490 ;
        RECT 2064.580 3153.170 2064.840 3153.490 ;
        RECT 2063.720 3152.890 2063.860 3153.170 ;
        RECT 2063.720 3152.750 2064.320 3152.890 ;
        RECT 2064.180 3105.290 2064.320 3152.750 ;
        RECT 2064.180 3105.150 2064.780 3105.290 ;
        RECT 2064.640 3056.930 2064.780 3105.150 ;
        RECT 2063.660 3056.610 2063.920 3056.930 ;
        RECT 2064.580 3056.610 2064.840 3056.930 ;
        RECT 2063.720 3056.330 2063.860 3056.610 ;
        RECT 2063.720 3056.190 2064.320 3056.330 ;
        RECT 2064.180 3042.990 2064.320 3056.190 ;
        RECT 2064.120 3042.670 2064.380 3042.990 ;
        RECT 2065.040 3008.330 2065.300 3008.650 ;
        RECT 2065.100 2994.710 2065.240 3008.330 ;
        RECT 2065.040 2994.390 2065.300 2994.710 ;
        RECT 2065.500 2946.450 2065.760 2946.770 ;
        RECT 2065.560 2912.430 2065.700 2946.450 ;
        RECT 2065.500 2912.110 2065.760 2912.430 ;
        RECT 2065.040 2911.430 2065.300 2911.750 ;
        RECT 2065.100 2863.210 2065.240 2911.430 ;
        RECT 2064.180 2863.070 2065.240 2863.210 ;
        RECT 2064.180 2849.610 2064.320 2863.070 ;
        RECT 2063.720 2849.470 2064.320 2849.610 ;
        RECT 2063.720 2815.870 2063.860 2849.470 ;
        RECT 2063.660 2815.550 2063.920 2815.870 ;
        RECT 2063.660 2814.870 2063.920 2815.190 ;
        RECT 2063.720 2801.250 2063.860 2814.870 ;
        RECT 2063.660 2800.930 2063.920 2801.250 ;
        RECT 2064.580 2752.990 2064.840 2753.310 ;
        RECT 2064.640 2718.290 2064.780 2752.990 ;
        RECT 2063.660 2717.970 2063.920 2718.290 ;
        RECT 2064.580 2717.970 2064.840 2718.290 ;
        RECT 2063.720 2670.350 2063.860 2717.970 ;
        RECT 2063.660 2670.030 2063.920 2670.350 ;
        RECT 2064.580 2670.030 2064.840 2670.350 ;
        RECT 2064.640 2622.410 2064.780 2670.030 ;
        RECT 2064.580 2622.090 2064.840 2622.410 ;
        RECT 2065.040 2621.750 2065.300 2622.070 ;
        RECT 2065.100 2608.325 2065.240 2621.750 ;
        RECT 2064.110 2607.955 2064.390 2608.325 ;
        RECT 2065.030 2607.955 2065.310 2608.325 ;
        RECT 2064.180 2560.190 2064.320 2607.955 ;
        RECT 2064.120 2559.870 2064.380 2560.190 ;
        RECT 2065.500 2559.870 2065.760 2560.190 ;
        RECT 1503.380 2517.710 1503.640 2518.030 ;
        RECT 1503.440 2500.000 1503.580 2517.710 ;
        RECT 2065.560 2517.690 2065.700 2559.870 ;
        RECT 2065.500 2517.370 2065.760 2517.690 ;
        RECT 1503.370 2496.000 1503.650 2500.000 ;
      LAYER via2 ;
        RECT 2064.110 2608.000 2064.390 2608.280 ;
        RECT 2065.030 2608.000 2065.310 2608.280 ;
      LAYER met3 ;
        RECT 2064.085 2608.290 2064.415 2608.305 ;
        RECT 2065.005 2608.290 2065.335 2608.305 ;
        RECT 2064.085 2607.990 2065.335 2608.290 ;
        RECT 2064.085 2607.975 2064.415 2607.990 ;
        RECT 2065.005 2607.975 2065.335 2607.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1524.510 3499.520 1524.830 3499.580 ;
        RECT 1743.930 3499.520 1744.250 3499.580 ;
        RECT 1524.510 3499.380 1744.250 3499.520 ;
        RECT 1524.510 3499.320 1524.830 3499.380 ;
        RECT 1743.930 3499.320 1744.250 3499.380 ;
      LAYER via ;
        RECT 1524.540 3499.320 1524.800 3499.580 ;
        RECT 1743.960 3499.320 1744.220 3499.580 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1743.810 3519.700 1744.370 3524.800 ;
=======
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3499.610 1744.160 3517.600 ;
        RECT 1524.540 3499.290 1524.800 3499.610 ;
        RECT 1743.960 3499.290 1744.220 3499.610 ;
        RECT 1523.150 2499.410 1523.430 2500.000 ;
        RECT 1524.600 2499.410 1524.740 3499.290 ;
        RECT 1523.150 2499.270 1524.740 2499.410 ;
        RECT 1523.150 2496.000 1523.430 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1420.165 3381.045 1420.335 3429.155 ;
        RECT 1531.485 2517.445 1531.655 2518.635 ;
        RECT 1531.945 2517.445 1532.115 2518.635 ;
      LAYER mcon ;
        RECT 1420.165 3428.985 1420.335 3429.155 ;
        RECT 1531.485 2518.465 1531.655 2518.635 ;
        RECT 1531.945 2518.465 1532.115 2518.635 ;
      LAYER met1 ;
        RECT 1418.710 3478.100 1419.030 3478.160 ;
        RECT 1419.630 3478.100 1419.950 3478.160 ;
        RECT 1418.710 3477.960 1419.950 3478.100 ;
        RECT 1418.710 3477.900 1419.030 3477.960 ;
        RECT 1419.630 3477.900 1419.950 3477.960 ;
        RECT 1419.630 3443.080 1419.950 3443.140 ;
        RECT 1420.550 3443.080 1420.870 3443.140 ;
        RECT 1419.630 3442.940 1420.870 3443.080 ;
        RECT 1419.630 3442.880 1419.950 3442.940 ;
        RECT 1420.550 3442.880 1420.870 3442.940 ;
        RECT 1420.105 3429.140 1420.395 3429.185 ;
        RECT 1420.550 3429.140 1420.870 3429.200 ;
        RECT 1420.105 3429.000 1420.870 3429.140 ;
        RECT 1420.105 3428.955 1420.395 3429.000 ;
        RECT 1420.550 3428.940 1420.870 3429.000 ;
        RECT 1420.090 3381.200 1420.410 3381.260 ;
        RECT 1419.895 3381.060 1420.410 3381.200 ;
        RECT 1420.090 3381.000 1420.410 3381.060 ;
        RECT 1420.090 3367.600 1420.410 3367.660 ;
        RECT 1421.010 3367.600 1421.330 3367.660 ;
        RECT 1420.090 3367.460 1421.330 3367.600 ;
        RECT 1420.090 3367.400 1420.410 3367.460 ;
        RECT 1421.010 3367.400 1421.330 3367.460 ;
        RECT 1420.090 3270.700 1420.410 3270.760 ;
        RECT 1421.010 3270.700 1421.330 3270.760 ;
        RECT 1420.090 3270.560 1421.330 3270.700 ;
        RECT 1420.090 3270.500 1420.410 3270.560 ;
        RECT 1421.010 3270.500 1421.330 3270.560 ;
        RECT 1419.630 3222.080 1419.950 3222.140 ;
        RECT 1421.010 3222.080 1421.330 3222.140 ;
        RECT 1419.630 3221.940 1421.330 3222.080 ;
        RECT 1419.630 3221.880 1419.950 3221.940 ;
        RECT 1421.010 3221.880 1421.330 3221.940 ;
        RECT 1419.630 3174.140 1419.950 3174.200 ;
        RECT 1421.010 3174.140 1421.330 3174.200 ;
        RECT 1419.630 3174.000 1421.330 3174.140 ;
        RECT 1419.630 3173.940 1419.950 3174.000 ;
        RECT 1421.010 3173.940 1421.330 3174.000 ;
        RECT 1419.630 3125.520 1419.950 3125.580 ;
        RECT 1421.010 3125.520 1421.330 3125.580 ;
        RECT 1419.630 3125.380 1421.330 3125.520 ;
        RECT 1419.630 3125.320 1419.950 3125.380 ;
        RECT 1421.010 3125.320 1421.330 3125.380 ;
        RECT 1419.630 3077.580 1419.950 3077.640 ;
        RECT 1421.010 3077.580 1421.330 3077.640 ;
        RECT 1419.630 3077.440 1421.330 3077.580 ;
        RECT 1419.630 3077.380 1419.950 3077.440 ;
        RECT 1421.010 3077.380 1421.330 3077.440 ;
        RECT 1419.630 3028.960 1419.950 3029.020 ;
        RECT 1421.010 3028.960 1421.330 3029.020 ;
        RECT 1419.630 3028.820 1421.330 3028.960 ;
        RECT 1419.630 3028.760 1419.950 3028.820 ;
        RECT 1421.010 3028.760 1421.330 3028.820 ;
        RECT 1419.630 2981.020 1419.950 2981.080 ;
        RECT 1421.010 2981.020 1421.330 2981.080 ;
        RECT 1419.630 2980.880 1421.330 2981.020 ;
        RECT 1419.630 2980.820 1419.950 2980.880 ;
        RECT 1421.010 2980.820 1421.330 2980.880 ;
        RECT 1419.630 2932.400 1419.950 2932.460 ;
        RECT 1421.010 2932.400 1421.330 2932.460 ;
        RECT 1419.630 2932.260 1421.330 2932.400 ;
        RECT 1419.630 2932.200 1419.950 2932.260 ;
        RECT 1421.010 2932.200 1421.330 2932.260 ;
        RECT 1419.630 2884.460 1419.950 2884.520 ;
        RECT 1421.010 2884.460 1421.330 2884.520 ;
        RECT 1419.630 2884.320 1421.330 2884.460 ;
        RECT 1419.630 2884.260 1419.950 2884.320 ;
        RECT 1421.010 2884.260 1421.330 2884.320 ;
        RECT 1419.630 2835.840 1419.950 2835.900 ;
        RECT 1421.010 2835.840 1421.330 2835.900 ;
        RECT 1419.630 2835.700 1421.330 2835.840 ;
        RECT 1419.630 2835.640 1419.950 2835.700 ;
        RECT 1421.010 2835.640 1421.330 2835.700 ;
        RECT 1419.630 2787.900 1419.950 2787.960 ;
        RECT 1421.010 2787.900 1421.330 2787.960 ;
        RECT 1419.630 2787.760 1421.330 2787.900 ;
        RECT 1419.630 2787.700 1419.950 2787.760 ;
        RECT 1421.010 2787.700 1421.330 2787.760 ;
        RECT 1419.630 2739.280 1419.950 2739.340 ;
        RECT 1421.010 2739.280 1421.330 2739.340 ;
        RECT 1419.630 2739.140 1421.330 2739.280 ;
        RECT 1419.630 2739.080 1419.950 2739.140 ;
        RECT 1421.010 2739.080 1421.330 2739.140 ;
        RECT 1419.630 2642.720 1419.950 2642.780 ;
        RECT 1421.010 2642.720 1421.330 2642.780 ;
        RECT 1419.630 2642.580 1421.330 2642.720 ;
        RECT 1419.630 2642.520 1419.950 2642.580 ;
        RECT 1421.010 2642.520 1421.330 2642.580 ;
        RECT 1419.630 2594.780 1419.950 2594.840 ;
        RECT 1421.010 2594.780 1421.330 2594.840 ;
        RECT 1419.630 2594.640 1421.330 2594.780 ;
        RECT 1419.630 2594.580 1419.950 2594.640 ;
        RECT 1421.010 2594.580 1421.330 2594.640 ;
        RECT 1420.090 2546.160 1420.410 2546.220 ;
        RECT 1421.010 2546.160 1421.330 2546.220 ;
        RECT 1420.090 2546.020 1421.330 2546.160 ;
        RECT 1420.090 2545.960 1420.410 2546.020 ;
        RECT 1421.010 2545.960 1421.330 2546.020 ;
        RECT 1531.425 2518.620 1531.715 2518.665 ;
        RECT 1527.820 2518.480 1531.715 2518.620 ;
        RECT 1420.090 2518.280 1420.410 2518.340 ;
        RECT 1527.820 2518.280 1527.960 2518.480 ;
        RECT 1531.425 2518.435 1531.715 2518.480 ;
        RECT 1531.885 2518.620 1532.175 2518.665 ;
        RECT 1541.070 2518.620 1541.390 2518.680 ;
        RECT 1531.885 2518.480 1541.390 2518.620 ;
        RECT 1531.885 2518.435 1532.175 2518.480 ;
        RECT 1541.070 2518.420 1541.390 2518.480 ;
        RECT 1420.090 2518.140 1527.960 2518.280 ;
        RECT 1420.090 2518.080 1420.410 2518.140 ;
        RECT 1531.425 2517.600 1531.715 2517.645 ;
        RECT 1531.885 2517.600 1532.175 2517.645 ;
        RECT 1531.425 2517.460 1532.175 2517.600 ;
        RECT 1531.425 2517.415 1531.715 2517.460 ;
        RECT 1531.885 2517.415 1532.175 2517.460 ;
      LAYER via ;
        RECT 1418.740 3477.900 1419.000 3478.160 ;
        RECT 1419.660 3477.900 1419.920 3478.160 ;
        RECT 1419.660 3442.880 1419.920 3443.140 ;
        RECT 1420.580 3442.880 1420.840 3443.140 ;
        RECT 1420.580 3428.940 1420.840 3429.200 ;
        RECT 1420.120 3381.000 1420.380 3381.260 ;
        RECT 1420.120 3367.400 1420.380 3367.660 ;
        RECT 1421.040 3367.400 1421.300 3367.660 ;
        RECT 1420.120 3270.500 1420.380 3270.760 ;
        RECT 1421.040 3270.500 1421.300 3270.760 ;
        RECT 1419.660 3221.880 1419.920 3222.140 ;
        RECT 1421.040 3221.880 1421.300 3222.140 ;
        RECT 1419.660 3173.940 1419.920 3174.200 ;
        RECT 1421.040 3173.940 1421.300 3174.200 ;
        RECT 1419.660 3125.320 1419.920 3125.580 ;
        RECT 1421.040 3125.320 1421.300 3125.580 ;
        RECT 1419.660 3077.380 1419.920 3077.640 ;
        RECT 1421.040 3077.380 1421.300 3077.640 ;
        RECT 1419.660 3028.760 1419.920 3029.020 ;
        RECT 1421.040 3028.760 1421.300 3029.020 ;
        RECT 1419.660 2980.820 1419.920 2981.080 ;
        RECT 1421.040 2980.820 1421.300 2981.080 ;
        RECT 1419.660 2932.200 1419.920 2932.460 ;
        RECT 1421.040 2932.200 1421.300 2932.460 ;
        RECT 1419.660 2884.260 1419.920 2884.520 ;
        RECT 1421.040 2884.260 1421.300 2884.520 ;
        RECT 1419.660 2835.640 1419.920 2835.900 ;
        RECT 1421.040 2835.640 1421.300 2835.900 ;
        RECT 1419.660 2787.700 1419.920 2787.960 ;
        RECT 1421.040 2787.700 1421.300 2787.960 ;
        RECT 1419.660 2739.080 1419.920 2739.340 ;
        RECT 1421.040 2739.080 1421.300 2739.340 ;
        RECT 1419.660 2642.520 1419.920 2642.780 ;
        RECT 1421.040 2642.520 1421.300 2642.780 ;
        RECT 1419.660 2594.580 1419.920 2594.840 ;
        RECT 1421.040 2594.580 1421.300 2594.840 ;
        RECT 1420.120 2545.960 1420.380 2546.220 ;
        RECT 1421.040 2545.960 1421.300 2546.220 ;
        RECT 1420.120 2518.080 1420.380 2518.340 ;
        RECT 1541.100 2518.420 1541.360 2518.680 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1419.050 3519.700 1419.610 3524.800 ;
=======
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3517.370 1419.400 3517.600 ;
        RECT 1418.800 3517.230 1419.400 3517.370 ;
        RECT 1418.800 3478.190 1418.940 3517.230 ;
        RECT 1418.740 3477.870 1419.000 3478.190 ;
        RECT 1419.660 3477.870 1419.920 3478.190 ;
        RECT 1419.720 3443.170 1419.860 3477.870 ;
        RECT 1419.660 3442.850 1419.920 3443.170 ;
        RECT 1420.580 3442.850 1420.840 3443.170 ;
        RECT 1420.640 3429.230 1420.780 3442.850 ;
        RECT 1420.580 3428.910 1420.840 3429.230 ;
        RECT 1420.120 3380.970 1420.380 3381.290 ;
        RECT 1420.180 3367.690 1420.320 3380.970 ;
        RECT 1420.120 3367.370 1420.380 3367.690 ;
        RECT 1421.040 3367.370 1421.300 3367.690 ;
        RECT 1421.100 3318.810 1421.240 3367.370 ;
        RECT 1420.180 3318.670 1421.240 3318.810 ;
        RECT 1420.180 3270.790 1420.320 3318.670 ;
        RECT 1420.120 3270.470 1420.380 3270.790 ;
        RECT 1421.040 3270.470 1421.300 3270.790 ;
        RECT 1421.100 3222.170 1421.240 3270.470 ;
        RECT 1419.660 3221.850 1419.920 3222.170 ;
        RECT 1421.040 3221.850 1421.300 3222.170 ;
        RECT 1419.720 3174.230 1419.860 3221.850 ;
        RECT 1419.660 3173.910 1419.920 3174.230 ;
        RECT 1421.040 3173.910 1421.300 3174.230 ;
        RECT 1421.100 3125.610 1421.240 3173.910 ;
        RECT 1419.660 3125.290 1419.920 3125.610 ;
        RECT 1421.040 3125.290 1421.300 3125.610 ;
        RECT 1419.720 3077.670 1419.860 3125.290 ;
        RECT 1419.660 3077.350 1419.920 3077.670 ;
        RECT 1421.040 3077.350 1421.300 3077.670 ;
        RECT 1421.100 3029.050 1421.240 3077.350 ;
        RECT 1419.660 3028.730 1419.920 3029.050 ;
        RECT 1421.040 3028.730 1421.300 3029.050 ;
        RECT 1419.720 2981.110 1419.860 3028.730 ;
        RECT 1419.660 2980.790 1419.920 2981.110 ;
        RECT 1421.040 2980.790 1421.300 2981.110 ;
        RECT 1421.100 2932.490 1421.240 2980.790 ;
        RECT 1419.660 2932.170 1419.920 2932.490 ;
        RECT 1421.040 2932.170 1421.300 2932.490 ;
        RECT 1419.720 2884.550 1419.860 2932.170 ;
        RECT 1419.660 2884.230 1419.920 2884.550 ;
        RECT 1421.040 2884.230 1421.300 2884.550 ;
        RECT 1421.100 2835.930 1421.240 2884.230 ;
        RECT 1419.660 2835.610 1419.920 2835.930 ;
        RECT 1421.040 2835.610 1421.300 2835.930 ;
        RECT 1419.720 2787.990 1419.860 2835.610 ;
        RECT 1419.660 2787.670 1419.920 2787.990 ;
        RECT 1421.040 2787.670 1421.300 2787.990 ;
        RECT 1421.100 2739.370 1421.240 2787.670 ;
        RECT 1419.660 2739.050 1419.920 2739.370 ;
        RECT 1421.040 2739.050 1421.300 2739.370 ;
        RECT 1419.720 2691.285 1419.860 2739.050 ;
        RECT 1419.650 2690.915 1419.930 2691.285 ;
        RECT 1421.030 2690.915 1421.310 2691.285 ;
        RECT 1421.100 2642.810 1421.240 2690.915 ;
        RECT 1419.660 2642.490 1419.920 2642.810 ;
        RECT 1421.040 2642.490 1421.300 2642.810 ;
        RECT 1419.720 2594.870 1419.860 2642.490 ;
        RECT 1419.660 2594.550 1419.920 2594.870 ;
        RECT 1421.040 2594.550 1421.300 2594.870 ;
        RECT 1421.100 2546.250 1421.240 2594.550 ;
        RECT 1420.120 2545.930 1420.380 2546.250 ;
        RECT 1421.040 2545.930 1421.300 2546.250 ;
        RECT 1420.180 2518.370 1420.320 2545.930 ;
        RECT 1541.100 2518.390 1541.360 2518.710 ;
        RECT 1420.120 2518.050 1420.380 2518.370 ;
        RECT 1541.160 2499.410 1541.300 2518.390 ;
        RECT 1542.930 2499.410 1543.210 2500.000 ;
        RECT 1541.160 2499.270 1543.210 2499.410 ;
        RECT 1542.930 2496.000 1543.210 2499.270 ;
      LAYER via2 ;
        RECT 1419.650 2690.960 1419.930 2691.240 ;
        RECT 1421.030 2690.960 1421.310 2691.240 ;
      LAYER met3 ;
        RECT 1419.625 2691.250 1419.955 2691.265 ;
        RECT 1421.005 2691.250 1421.335 2691.265 ;
        RECT 1419.625 2690.950 1421.335 2691.250 ;
        RECT 1419.625 2690.935 1419.955 2690.950 ;
        RECT 1421.005 2690.935 1421.335 2690.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1399.850 381.040 1400.170 381.100 ;
        RECT 1405.830 381.040 1406.150 381.100 ;
        RECT 1399.850 380.900 1406.150 381.040 ;
        RECT 1399.850 380.840 1400.170 380.900 ;
        RECT 1405.830 380.840 1406.150 380.900 ;
        RECT 2090.310 380.700 2090.630 380.760 ;
        RECT 2124.810 380.700 2125.130 380.760 ;
        RECT 2090.310 380.560 2125.130 380.700 ;
        RECT 2090.310 380.500 2090.630 380.560 ;
        RECT 2124.810 380.500 2125.130 380.560 ;
        RECT 1702.070 380.360 1702.390 380.420 ;
        RECT 1711.730 380.360 1712.050 380.420 ;
        RECT 1702.070 380.220 1712.050 380.360 ;
        RECT 1702.070 380.160 1702.390 380.220 ;
        RECT 1711.730 380.160 1712.050 380.220 ;
        RECT 1798.670 380.360 1798.990 380.420 ;
        RECT 1801.890 380.360 1802.210 380.420 ;
        RECT 1798.670 380.220 1802.210 380.360 ;
        RECT 1798.670 380.160 1798.990 380.220 ;
        RECT 1801.890 380.160 1802.210 380.220 ;
        RECT 1932.070 380.020 1932.390 380.080 ;
        RECT 1946.330 380.020 1946.650 380.080 ;
        RECT 1932.070 379.880 1946.650 380.020 ;
        RECT 1932.070 379.820 1932.390 379.880 ;
        RECT 1946.330 379.820 1946.650 379.880 ;
      LAYER via ;
        RECT 1399.880 380.840 1400.140 381.100 ;
        RECT 1405.860 380.840 1406.120 381.100 ;
        RECT 2090.340 380.500 2090.600 380.760 ;
        RECT 2124.840 380.500 2125.100 380.760 ;
        RECT 1702.100 380.160 1702.360 380.420 ;
        RECT 1711.760 380.160 1712.020 380.420 ;
        RECT 1798.700 380.160 1798.960 380.420 ;
        RECT 1801.920 380.160 1802.180 380.420 ;
        RECT 1932.100 379.820 1932.360 380.080 ;
        RECT 1946.360 379.820 1946.620 380.080 ;
      LAYER met2 ;
        RECT 1185.970 2498.050 1186.250 2500.000 ;
        RECT 1186.430 2498.050 1186.710 2498.165 ;
        RECT 1185.970 2497.910 1186.710 2498.050 ;
        RECT 1185.970 2496.000 1186.250 2497.910 ;
        RECT 1186.430 2497.795 1186.710 2497.910 ;
        RECT 1200.230 404.075 1200.510 404.445 ;
        RECT 1200.300 380.645 1200.440 404.075 ;
        RECT 2028.230 382.315 2028.510 382.685 ;
        RECT 1296.830 380.955 1297.110 381.325 ;
        RECT 1399.870 380.955 1400.150 381.325 ;
        RECT 1405.850 380.955 1406.130 381.325 ;
        RECT 1593.070 380.955 1593.350 381.325 ;
        RECT 1946.350 380.955 1946.630 381.325 ;
        RECT 1200.230 380.275 1200.510 380.645 ;
        RECT 1296.900 379.965 1297.040 380.955 ;
        RECT 1399.880 380.810 1400.140 380.955 ;
        RECT 1405.860 380.810 1406.120 380.955 ;
        RECT 1593.140 379.965 1593.280 380.955 ;
        RECT 1702.090 380.275 1702.370 380.645 ;
        RECT 1711.750 380.275 1712.030 380.645 ;
        RECT 1798.690 380.275 1798.970 380.645 ;
        RECT 1801.910 380.275 1802.190 380.645 ;
        RECT 1895.290 380.275 1895.570 380.645 ;
        RECT 1702.100 380.130 1702.360 380.275 ;
        RECT 1711.760 380.130 1712.020 380.275 ;
        RECT 1798.700 380.130 1798.960 380.275 ;
        RECT 1801.920 380.130 1802.180 380.275 ;
        RECT 1296.830 379.595 1297.110 379.965 ;
        RECT 1593.070 379.595 1593.350 379.965 ;
        RECT 1895.360 378.605 1895.500 380.275 ;
        RECT 1946.420 380.110 1946.560 380.955 ;
        RECT 2028.300 380.645 2028.440 382.315 ;
        RECT 2052.610 381.635 2052.890 382.005 ;
        RECT 2028.230 380.275 2028.510 380.645 ;
        RECT 1932.100 379.965 1932.360 380.110 ;
        RECT 1932.090 379.595 1932.370 379.965 ;
        RECT 1946.360 379.790 1946.620 380.110 ;
        RECT 2052.680 379.965 2052.820 381.635 ;
        RECT 2124.830 380.955 2125.110 381.325 ;
        RECT 2124.900 380.790 2125.040 380.955 ;
        RECT 2090.340 380.645 2090.600 380.790 ;
        RECT 2090.330 380.275 2090.610 380.645 ;
        RECT 2124.840 380.470 2125.100 380.790 ;
        RECT 2052.610 379.595 2052.890 379.965 ;
        RECT 1895.290 378.235 1895.570 378.605 ;
      LAYER via2 ;
        RECT 1186.430 2497.840 1186.710 2498.120 ;
        RECT 1200.230 404.120 1200.510 404.400 ;
        RECT 2028.230 382.360 2028.510 382.640 ;
        RECT 1296.830 381.000 1297.110 381.280 ;
        RECT 1399.870 381.000 1400.150 381.280 ;
        RECT 1405.850 381.000 1406.130 381.280 ;
        RECT 1593.070 381.000 1593.350 381.280 ;
        RECT 1946.350 381.000 1946.630 381.280 ;
        RECT 1200.230 380.320 1200.510 380.600 ;
        RECT 1702.090 380.320 1702.370 380.600 ;
        RECT 1711.750 380.320 1712.030 380.600 ;
        RECT 1798.690 380.320 1798.970 380.600 ;
        RECT 1801.910 380.320 1802.190 380.600 ;
        RECT 1895.290 380.320 1895.570 380.600 ;
        RECT 1296.830 379.640 1297.110 379.920 ;
        RECT 1593.070 379.640 1593.350 379.920 ;
        RECT 2052.610 381.680 2052.890 381.960 ;
        RECT 2028.230 380.320 2028.510 380.600 ;
        RECT 1932.090 379.640 1932.370 379.920 ;
        RECT 2124.830 381.000 2125.110 381.280 ;
        RECT 2090.330 380.320 2090.610 380.600 ;
        RECT 2052.610 379.640 2052.890 379.920 ;
        RECT 1895.290 378.280 1895.570 378.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 380.540 2924.800 381.740 ;
=======
        RECT 1186.405 2498.140 1186.735 2498.145 ;
        RECT 1186.150 2498.130 1186.735 2498.140 ;
        RECT 1185.950 2497.830 1186.735 2498.130 ;
        RECT 1186.150 2497.820 1186.735 2497.830 ;
        RECT 1186.405 2497.815 1186.735 2497.820 ;
        RECT 1186.150 404.410 1186.530 404.420 ;
        RECT 1200.205 404.410 1200.535 404.425 ;
        RECT 1186.150 404.110 1200.535 404.410 ;
        RECT 1186.150 404.100 1186.530 404.110 ;
        RECT 1200.205 404.095 1200.535 404.110 ;
        RECT 1980.110 382.650 1980.490 382.660 ;
        RECT 2028.205 382.650 2028.535 382.665 ;
        RECT 1980.110 382.350 2028.535 382.650 ;
        RECT 1980.110 382.340 1980.490 382.350 ;
        RECT 2028.205 382.335 2028.535 382.350 ;
        RECT 2052.585 381.970 2052.915 381.985 ;
        RECT 2028.910 381.670 2052.915 381.970 ;
        RECT 1296.805 381.290 1297.135 381.305 ;
        RECT 1399.845 381.290 1400.175 381.305 ;
        RECT 1248.750 380.990 1297.135 381.290 ;
        RECT 1200.205 380.610 1200.535 380.625 ;
        RECT 1200.205 380.310 1225.130 380.610 ;
        RECT 1200.205 380.295 1200.535 380.310 ;
        RECT 1224.830 379.930 1225.130 380.310 ;
        RECT 1248.750 379.930 1249.050 380.990 ;
        RECT 1296.805 380.975 1297.135 380.990 ;
        RECT 1366.510 380.990 1400.175 381.290 ;
        RECT 1224.830 379.630 1249.050 379.930 ;
        RECT 1296.805 379.930 1297.135 379.945 ;
        RECT 1366.510 379.930 1366.810 380.990 ;
        RECT 1399.845 380.975 1400.175 380.990 ;
        RECT 1405.825 381.290 1406.155 381.305 ;
        RECT 1593.045 381.290 1593.375 381.305 ;
        RECT 1405.825 380.990 1593.375 381.290 ;
        RECT 1405.825 380.975 1406.155 380.990 ;
        RECT 1593.045 380.975 1593.375 380.990 ;
        RECT 1946.325 381.290 1946.655 381.305 ;
        RECT 1980.110 381.290 1980.490 381.300 ;
        RECT 1946.325 380.990 1980.490 381.290 ;
        RECT 1946.325 380.975 1946.655 380.990 ;
        RECT 1980.110 380.980 1980.490 380.990 ;
        RECT 1702.065 380.610 1702.395 380.625 ;
        RECT 1656.310 380.310 1702.395 380.610 ;
        RECT 1296.805 379.630 1366.810 379.930 ;
        RECT 1593.045 379.930 1593.375 379.945 ;
        RECT 1656.310 379.930 1656.610 380.310 ;
        RECT 1702.065 380.295 1702.395 380.310 ;
        RECT 1711.725 380.610 1712.055 380.625 ;
        RECT 1798.665 380.610 1798.995 380.625 ;
        RECT 1711.725 380.310 1738.490 380.610 ;
        RECT 1711.725 380.295 1712.055 380.310 ;
        RECT 1593.045 379.630 1656.610 379.930 ;
        RECT 1738.190 379.930 1738.490 380.310 ;
        RECT 1752.910 380.310 1798.995 380.610 ;
        RECT 1752.910 379.930 1753.210 380.310 ;
        RECT 1798.665 380.295 1798.995 380.310 ;
        RECT 1801.885 380.610 1802.215 380.625 ;
        RECT 1895.265 380.610 1895.595 380.625 ;
        RECT 1801.885 380.310 1835.090 380.610 ;
        RECT 1801.885 380.295 1802.215 380.310 ;
        RECT 1738.190 379.630 1753.210 379.930 ;
        RECT 1834.790 379.930 1835.090 380.310 ;
        RECT 1849.510 380.310 1895.595 380.610 ;
        RECT 1849.510 379.930 1849.810 380.310 ;
        RECT 1895.265 380.295 1895.595 380.310 ;
        RECT 2028.205 380.610 2028.535 380.625 ;
        RECT 2028.910 380.610 2029.210 381.670 ;
        RECT 2052.585 381.655 2052.915 381.670 ;
        RECT 2124.805 381.290 2125.135 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2124.805 380.990 2159.850 381.290 ;
        RECT 2124.805 380.975 2125.135 380.990 ;
        RECT 2090.305 380.610 2090.635 380.625 ;
        RECT 2028.205 380.310 2029.210 380.610 ;
        RECT 2076.750 380.310 2090.635 380.610 ;
        RECT 2159.550 380.610 2159.850 380.990 ;
        RECT 2208.310 380.990 2256.450 381.290 ;
        RECT 2159.550 380.310 2207.690 380.610 ;
        RECT 2028.205 380.295 2028.535 380.310 ;
        RECT 1932.065 379.930 1932.395 379.945 ;
        RECT 1834.790 379.630 1849.810 379.930 ;
        RECT 1931.390 379.630 1932.395 379.930 ;
        RECT 1296.805 379.615 1297.135 379.630 ;
        RECT 1593.045 379.615 1593.375 379.630 ;
        RECT 1895.265 378.570 1895.595 378.585 ;
        RECT 1931.390 378.570 1931.690 379.630 ;
        RECT 1932.065 379.615 1932.395 379.630 ;
        RECT 2052.585 379.930 2052.915 379.945 ;
        RECT 2076.750 379.930 2077.050 380.310 ;
        RECT 2090.305 380.295 2090.635 380.310 ;
        RECT 2052.585 379.630 2077.050 379.930 ;
        RECT 2207.390 379.930 2207.690 380.310 ;
        RECT 2208.310 379.930 2208.610 380.990 ;
        RECT 2256.150 380.610 2256.450 380.990 ;
        RECT 2304.910 380.990 2353.050 381.290 ;
        RECT 2256.150 380.310 2304.290 380.610 ;
        RECT 2207.390 379.630 2208.610 379.930 ;
        RECT 2303.990 379.930 2304.290 380.310 ;
        RECT 2304.910 379.930 2305.210 380.990 ;
        RECT 2352.750 380.610 2353.050 380.990 ;
        RECT 2401.510 380.990 2449.650 381.290 ;
        RECT 2352.750 380.310 2400.890 380.610 ;
        RECT 2303.990 379.630 2305.210 379.930 ;
        RECT 2400.590 379.930 2400.890 380.310 ;
        RECT 2401.510 379.930 2401.810 380.990 ;
        RECT 2449.350 380.610 2449.650 380.990 ;
        RECT 2498.110 380.990 2546.250 381.290 ;
        RECT 2449.350 380.310 2497.490 380.610 ;
        RECT 2400.590 379.630 2401.810 379.930 ;
        RECT 2497.190 379.930 2497.490 380.310 ;
        RECT 2498.110 379.930 2498.410 380.990 ;
        RECT 2545.950 380.610 2546.250 380.990 ;
        RECT 2594.710 380.990 2642.850 381.290 ;
        RECT 2545.950 380.310 2594.090 380.610 ;
        RECT 2497.190 379.630 2498.410 379.930 ;
        RECT 2593.790 379.930 2594.090 380.310 ;
        RECT 2594.710 379.930 2595.010 380.990 ;
        RECT 2642.550 380.610 2642.850 380.990 ;
        RECT 2691.310 380.990 2739.450 381.290 ;
        RECT 2642.550 380.310 2690.690 380.610 ;
        RECT 2593.790 379.630 2595.010 379.930 ;
        RECT 2690.390 379.930 2690.690 380.310 ;
        RECT 2691.310 379.930 2691.610 380.990 ;
        RECT 2739.150 380.610 2739.450 380.990 ;
        RECT 2787.910 380.990 2836.050 381.290 ;
        RECT 2739.150 380.310 2787.290 380.610 ;
        RECT 2690.390 379.630 2691.610 379.930 ;
        RECT 2786.990 379.930 2787.290 380.310 ;
        RECT 2787.910 379.930 2788.210 380.990 ;
        RECT 2835.750 380.610 2836.050 380.990 ;
        RECT 2916.710 380.990 2924.800 381.290 ;
        RECT 2916.710 380.610 2917.010 380.990 ;
        RECT 2835.750 380.310 2883.890 380.610 ;
        RECT 2786.990 379.630 2788.210 379.930 ;
        RECT 2883.590 379.930 2883.890 380.310 ;
        RECT 2884.510 380.310 2917.010 380.610 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2884.510 379.930 2884.810 380.310 ;
        RECT 2883.590 379.630 2884.810 379.930 ;
        RECT 2052.585 379.615 2052.915 379.630 ;
        RECT 1895.265 378.270 1931.690 378.570 ;
        RECT 1895.265 378.255 1895.595 378.270 ;
      LAYER via3 ;
        RECT 1186.180 2497.820 1186.500 2498.140 ;
        RECT 1186.180 404.100 1186.500 404.420 ;
        RECT 1980.140 382.340 1980.460 382.660 ;
        RECT 1980.140 380.980 1980.460 381.300 ;
      LAYER met4 ;
        RECT 1186.175 2497.815 1186.505 2498.145 ;
        RECT 1186.190 404.425 1186.490 2497.815 ;
        RECT 1186.175 404.095 1186.505 404.425 ;
        RECT 1980.135 382.335 1980.465 382.665 ;
        RECT 1980.150 381.305 1980.450 382.335 ;
        RECT 1980.135 380.975 1980.465 381.305 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1555.405 2517.785 1556.495 2517.955 ;
        RECT 1555.405 2517.445 1555.575 2517.785 ;
      LAYER mcon ;
        RECT 1556.325 2517.785 1556.495 2517.955 ;
      LAYER met1 ;
        RECT 1094.870 3500.540 1095.190 3500.600 ;
        RECT 1541.990 3500.540 1542.310 3500.600 ;
        RECT 1094.870 3500.400 1542.310 3500.540 ;
        RECT 1094.870 3500.340 1095.190 3500.400 ;
        RECT 1541.990 3500.340 1542.310 3500.400 ;
        RECT 1556.265 2517.940 1556.555 2517.985 ;
        RECT 1563.150 2517.940 1563.470 2518.000 ;
        RECT 1556.265 2517.800 1563.470 2517.940 ;
        RECT 1556.265 2517.755 1556.555 2517.800 ;
        RECT 1563.150 2517.740 1563.470 2517.800 ;
        RECT 1541.990 2517.600 1542.310 2517.660 ;
        RECT 1555.345 2517.600 1555.635 2517.645 ;
        RECT 1541.990 2517.460 1555.635 2517.600 ;
        RECT 1541.990 2517.400 1542.310 2517.460 ;
        RECT 1555.345 2517.415 1555.635 2517.460 ;
      LAYER via ;
        RECT 1094.900 3500.340 1095.160 3500.600 ;
        RECT 1542.020 3500.340 1542.280 3500.600 ;
        RECT 1563.180 2517.740 1563.440 2518.000 ;
        RECT 1542.020 2517.400 1542.280 2517.660 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1094.750 3519.700 1095.310 3524.800 ;
=======
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3500.630 1095.100 3517.600 ;
        RECT 1094.900 3500.310 1095.160 3500.630 ;
        RECT 1542.020 3500.310 1542.280 3500.630 ;
        RECT 1542.080 2517.690 1542.220 3500.310 ;
        RECT 1563.180 2517.710 1563.440 2518.030 ;
        RECT 1542.020 2517.370 1542.280 2517.690 ;
        RECT 1563.240 2500.000 1563.380 2517.710 ;
        RECT 1563.170 2496.000 1563.450 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 770.570 3504.620 770.890 3504.680 ;
        RECT 1562.690 3504.620 1563.010 3504.680 ;
        RECT 770.570 3504.480 1563.010 3504.620 ;
        RECT 770.570 3504.420 770.890 3504.480 ;
        RECT 1562.690 3504.420 1563.010 3504.480 ;
        RECT 1564.530 2518.280 1564.850 2518.340 ;
        RECT 1582.930 2518.280 1583.250 2518.340 ;
        RECT 1564.530 2518.140 1583.250 2518.280 ;
        RECT 1564.530 2518.080 1564.850 2518.140 ;
        RECT 1582.930 2518.080 1583.250 2518.140 ;
      LAYER via ;
        RECT 770.600 3504.420 770.860 3504.680 ;
        RECT 1562.720 3504.420 1562.980 3504.680 ;
        RECT 1564.560 2518.080 1564.820 2518.340 ;
        RECT 1582.960 2518.080 1583.220 2518.340 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 770.450 3519.700 771.010 3524.800 ;
=======
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3504.710 770.800 3517.600 ;
        RECT 770.600 3504.390 770.860 3504.710 ;
        RECT 1562.720 3504.390 1562.980 3504.710 ;
        RECT 1562.780 2518.450 1562.920 3504.390 ;
        RECT 1562.780 2518.310 1563.840 2518.450 ;
        RECT 1563.700 2517.770 1563.840 2518.310 ;
        RECT 1564.560 2518.050 1564.820 2518.370 ;
        RECT 1582.960 2518.050 1583.220 2518.370 ;
        RECT 1564.620 2517.770 1564.760 2518.050 ;
        RECT 1563.700 2517.630 1564.760 2517.770 ;
        RECT 1583.020 2500.000 1583.160 2518.050 ;
        RECT 1582.950 2496.000 1583.230 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.810 3502.920 446.130 3502.980 ;
        RECT 1583.390 3502.920 1583.710 3502.980 ;
        RECT 445.810 3502.780 1583.710 3502.920 ;
        RECT 445.810 3502.720 446.130 3502.780 ;
        RECT 1583.390 3502.720 1583.710 3502.780 ;
        RECT 1583.390 2518.280 1583.710 2518.340 ;
        RECT 1602.710 2518.280 1603.030 2518.340 ;
        RECT 1583.390 2518.140 1603.030 2518.280 ;
        RECT 1583.390 2518.080 1583.710 2518.140 ;
        RECT 1602.710 2518.080 1603.030 2518.140 ;
      LAYER via ;
        RECT 445.840 3502.720 446.100 3502.980 ;
        RECT 1583.420 3502.720 1583.680 3502.980 ;
        RECT 1583.420 2518.080 1583.680 2518.340 ;
        RECT 1602.740 2518.080 1603.000 2518.340 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 445.690 3519.700 446.250 3524.800 ;
=======
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3503.010 446.040 3517.600 ;
        RECT 445.840 3502.690 446.100 3503.010 ;
        RECT 1583.420 3502.690 1583.680 3503.010 ;
        RECT 1583.480 2518.370 1583.620 3502.690 ;
        RECT 1583.420 2518.050 1583.680 2518.370 ;
        RECT 1602.740 2518.050 1603.000 2518.370 ;
        RECT 1602.800 2500.000 1602.940 2518.050 ;
        RECT 1602.730 2496.000 1603.010 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1604.090 2518.280 1604.410 2518.340 ;
        RECT 1622.490 2518.280 1622.810 2518.340 ;
        RECT 1604.090 2518.140 1622.810 2518.280 ;
        RECT 1604.090 2518.080 1604.410 2518.140 ;
        RECT 1622.490 2518.080 1622.810 2518.140 ;
      LAYER via ;
        RECT 1604.120 2518.080 1604.380 2518.340 ;
        RECT 1622.520 2518.080 1622.780 2518.340 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 121.390 3519.700 121.950 3524.800 ;
=======
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3502.525 121.740 3517.600 ;
        RECT 121.530 3502.155 121.810 3502.525 ;
        RECT 1604.110 3502.155 1604.390 3502.525 ;
        RECT 1604.180 2518.370 1604.320 3502.155 ;
        RECT 1604.120 2518.050 1604.380 2518.370 ;
        RECT 1622.520 2518.050 1622.780 2518.370 ;
        RECT 1622.580 2500.000 1622.720 2518.050 ;
        RECT 1622.510 2496.000 1622.790 2500.000 ;
      LAYER via2 ;
        RECT 121.530 3502.200 121.810 3502.480 ;
        RECT 1604.110 3502.200 1604.390 3502.480 ;
      LAYER met3 ;
        RECT 121.505 3502.490 121.835 3502.505 ;
        RECT 1604.085 3502.490 1604.415 3502.505 ;
        RECT 121.505 3502.190 1604.415 3502.490 ;
        RECT 121.505 3502.175 121.835 3502.190 ;
        RECT 1604.085 3502.175 1604.415 3502.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 1642.270 3339.720 1642.590 3339.780 ;
        RECT 17.090 3339.580 1642.590 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 1642.270 3339.520 1642.590 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 1642.300 3339.520 1642.560 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 1642.300 3339.490 1642.560 3339.810 ;
        RECT 1642.360 2500.000 1642.500 3339.490 ;
        RECT 1642.290 2496.000 1642.570 2500.000 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3339.220 0.300 3340.420 ;
=======
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 1656.070 3050.040 1656.390 3050.100 ;
        RECT 17.090 3049.900 1656.390 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 1656.070 3049.840 1656.390 3049.900 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 1656.100 3049.840 1656.360 3050.100 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 1656.100 3049.810 1656.360 3050.130 ;
        RECT 1656.160 2502.130 1656.300 3049.810 ;
        RECT 1656.160 2501.990 1660.440 2502.130 ;
        RECT 1660.300 2499.410 1660.440 2501.990 ;
        RECT 1662.070 2499.410 1662.350 2500.000 ;
        RECT 1660.300 2499.270 1662.350 2499.410 ;
        RECT 1662.070 2496.000 1662.350 2499.270 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3051.580 0.300 3052.780 ;
=======
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2760.360 16.030 2760.420 ;
        RECT 1676.770 2760.360 1677.090 2760.420 ;
        RECT 15.710 2760.220 1677.090 2760.360 ;
        RECT 15.710 2760.160 16.030 2760.220 ;
        RECT 1676.770 2760.160 1677.090 2760.220 ;
      LAYER via ;
        RECT 15.740 2760.160 16.000 2760.420 ;
        RECT 1676.800 2760.160 1677.060 2760.420 ;
      LAYER met2 ;
        RECT 15.730 2765.035 16.010 2765.405 ;
        RECT 15.800 2760.450 15.940 2765.035 ;
        RECT 15.740 2760.130 16.000 2760.450 ;
        RECT 1676.800 2760.130 1677.060 2760.450 ;
        RECT 1676.860 2498.730 1677.000 2760.130 ;
        RECT 1681.850 2498.730 1682.130 2500.000 ;
        RECT 1676.860 2498.590 1682.130 2498.730 ;
        RECT 1681.850 2496.000 1682.130 2498.590 ;
      LAYER via2 ;
        RECT 15.730 2765.080 16.010 2765.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2764.620 0.300 2765.820 ;
=======
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 15.705 2765.370 16.035 2765.385 ;
        RECT -4.800 2765.070 16.035 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 15.705 2765.055 16.035 2765.070 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 21.690 2513.180 22.010 2513.240 ;
        RECT 1701.610 2513.180 1701.930 2513.240 ;
        RECT 21.690 2513.040 1701.930 2513.180 ;
        RECT 21.690 2512.980 22.010 2513.040 ;
        RECT 1701.610 2512.980 1701.930 2513.040 ;
        RECT 13.870 2477.820 14.190 2477.880 ;
        RECT 21.690 2477.820 22.010 2477.880 ;
        RECT 13.870 2477.680 22.010 2477.820 ;
        RECT 13.870 2477.620 14.190 2477.680 ;
        RECT 21.690 2477.620 22.010 2477.680 ;
      LAYER via ;
        RECT 21.720 2512.980 21.980 2513.240 ;
        RECT 1701.640 2512.980 1701.900 2513.240 ;
        RECT 13.900 2477.620 14.160 2477.880 ;
        RECT 21.720 2477.620 21.980 2477.880 ;
      LAYER met2 ;
        RECT 21.720 2512.950 21.980 2513.270 ;
        RECT 1701.640 2512.950 1701.900 2513.270 ;
        RECT 21.780 2477.910 21.920 2512.950 ;
        RECT 1701.700 2500.000 1701.840 2512.950 ;
        RECT 1701.630 2496.000 1701.910 2500.000 ;
        RECT 13.900 2477.765 14.160 2477.910 ;
        RECT 13.890 2477.395 14.170 2477.765 ;
        RECT 21.720 2477.590 21.980 2477.910 ;
      LAYER via2 ;
        RECT 13.890 2477.440 14.170 2477.720 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2476.980 0.300 2478.180 ;
=======
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 13.865 2477.730 14.195 2477.745 ;
        RECT -4.800 2477.430 14.195 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 13.865 2477.415 14.195 2477.430 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 22.610 2512.500 22.930 2512.560 ;
        RECT 1721.390 2512.500 1721.710 2512.560 ;
        RECT 22.610 2512.360 1721.710 2512.500 ;
        RECT 22.610 2512.300 22.930 2512.360 ;
        RECT 1721.390 2512.300 1721.710 2512.360 ;
        RECT 13.870 2190.180 14.190 2190.240 ;
        RECT 22.610 2190.180 22.930 2190.240 ;
        RECT 13.870 2190.040 22.930 2190.180 ;
        RECT 13.870 2189.980 14.190 2190.040 ;
        RECT 22.610 2189.980 22.930 2190.040 ;
      LAYER via ;
        RECT 22.640 2512.300 22.900 2512.560 ;
        RECT 1721.420 2512.300 1721.680 2512.560 ;
        RECT 13.900 2189.980 14.160 2190.240 ;
        RECT 22.640 2189.980 22.900 2190.240 ;
      LAYER met2 ;
        RECT 22.640 2512.270 22.900 2512.590 ;
        RECT 1721.420 2512.270 1721.680 2512.590 ;
        RECT 22.700 2190.270 22.840 2512.270 ;
        RECT 1721.480 2500.000 1721.620 2512.270 ;
        RECT 1721.410 2496.000 1721.690 2500.000 ;
        RECT 13.900 2190.125 14.160 2190.270 ;
        RECT 13.890 2189.755 14.170 2190.125 ;
        RECT 22.640 2189.950 22.900 2190.270 ;
      LAYER via2 ;
        RECT 13.890 2189.800 14.170 2190.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2189.340 0.300 2190.540 ;
=======
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 13.865 2190.090 14.195 2190.105 ;
        RECT -4.800 2189.790 14.195 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 13.865 2189.775 14.195 2189.790 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 2511.820 15.570 2511.880 ;
        RECT 1741.630 2511.820 1741.950 2511.880 ;
        RECT 15.250 2511.680 1741.950 2511.820 ;
        RECT 15.250 2511.620 15.570 2511.680 ;
        RECT 1741.630 2511.620 1741.950 2511.680 ;
      LAYER via ;
        RECT 15.280 2511.620 15.540 2511.880 ;
        RECT 1741.660 2511.620 1741.920 2511.880 ;
      LAYER met2 ;
        RECT 15.280 2511.590 15.540 2511.910 ;
        RECT 1741.660 2511.590 1741.920 2511.910 ;
        RECT 15.340 1903.165 15.480 2511.590 ;
        RECT 1741.720 2500.000 1741.860 2511.590 ;
        RECT 1741.650 2496.000 1741.930 2500.000 ;
        RECT 15.270 1902.795 15.550 1903.165 ;
      LAYER via2 ;
        RECT 15.270 1902.840 15.550 1903.120 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1902.380 0.300 1903.580 ;
=======
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 15.245 1903.130 15.575 1903.145 ;
        RECT -4.800 1902.830 15.575 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 15.245 1902.815 15.575 1902.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1352.010 615.640 1352.330 615.700 ;
        RECT 1386.510 615.640 1386.830 615.700 ;
        RECT 1352.010 615.500 1386.830 615.640 ;
        RECT 1352.010 615.440 1352.330 615.500 ;
        RECT 1386.510 615.440 1386.830 615.500 ;
        RECT 1593.970 615.300 1594.290 615.360 ;
        RECT 1607.770 615.300 1608.090 615.360 ;
        RECT 1593.970 615.160 1608.090 615.300 ;
        RECT 1593.970 615.100 1594.290 615.160 ;
        RECT 1607.770 615.100 1608.090 615.160 ;
        RECT 2090.310 615.300 2090.630 615.360 ;
        RECT 2124.810 615.300 2125.130 615.360 ;
        RECT 2090.310 615.160 2125.130 615.300 ;
        RECT 2090.310 615.100 2090.630 615.160 ;
        RECT 2124.810 615.100 2125.130 615.160 ;
        RECT 1702.070 614.960 1702.390 615.020 ;
        RECT 1711.730 614.960 1712.050 615.020 ;
        RECT 1702.070 614.820 1712.050 614.960 ;
        RECT 1702.070 614.760 1702.390 614.820 ;
        RECT 1711.730 614.760 1712.050 614.820 ;
        RECT 1798.670 614.960 1798.990 615.020 ;
        RECT 1801.890 614.960 1802.210 615.020 ;
        RECT 1798.670 614.820 1802.210 614.960 ;
        RECT 1798.670 614.760 1798.990 614.820 ;
        RECT 1801.890 614.760 1802.210 614.820 ;
        RECT 1932.070 614.620 1932.390 614.680 ;
        RECT 1946.330 614.620 1946.650 614.680 ;
        RECT 1932.070 614.480 1946.650 614.620 ;
        RECT 1932.070 614.420 1932.390 614.480 ;
        RECT 1946.330 614.420 1946.650 614.480 ;
      LAYER via ;
        RECT 1352.040 615.440 1352.300 615.700 ;
        RECT 1386.540 615.440 1386.800 615.700 ;
        RECT 1594.000 615.100 1594.260 615.360 ;
        RECT 1607.800 615.100 1608.060 615.360 ;
        RECT 2090.340 615.100 2090.600 615.360 ;
        RECT 2124.840 615.100 2125.100 615.360 ;
        RECT 1702.100 614.760 1702.360 615.020 ;
        RECT 1711.760 614.760 1712.020 615.020 ;
        RECT 1798.700 614.760 1798.960 615.020 ;
        RECT 1801.920 614.760 1802.180 615.020 ;
        RECT 1932.100 614.420 1932.360 614.680 ;
        RECT 1946.360 614.420 1946.620 614.680 ;
      LAYER met2 ;
        RECT 1205.750 2498.050 1206.030 2500.000 ;
        RECT 1206.210 2498.050 1206.490 2498.165 ;
        RECT 1205.750 2497.910 1206.490 2498.050 ;
        RECT 1205.750 2496.000 1206.030 2497.910 ;
        RECT 1206.210 2497.795 1206.490 2497.910 ;
        RECT 2028.230 616.915 2028.510 617.285 ;
        RECT 1352.030 615.555 1352.310 615.925 ;
        RECT 1352.040 615.410 1352.300 615.555 ;
        RECT 1386.540 615.410 1386.800 615.730 ;
        RECT 1946.350 615.555 1946.630 615.925 ;
        RECT 1386.600 615.245 1386.740 615.410 ;
        RECT 1594.000 615.245 1594.260 615.390 ;
        RECT 1607.800 615.245 1608.060 615.390 ;
        RECT 1386.530 614.875 1386.810 615.245 ;
        RECT 1593.990 614.875 1594.270 615.245 ;
        RECT 1607.790 614.875 1608.070 615.245 ;
        RECT 1702.090 614.875 1702.370 615.245 ;
        RECT 1711.750 614.875 1712.030 615.245 ;
        RECT 1798.690 614.875 1798.970 615.245 ;
        RECT 1801.910 614.875 1802.190 615.245 ;
        RECT 1895.290 614.875 1895.570 615.245 ;
        RECT 1702.100 614.730 1702.360 614.875 ;
        RECT 1711.760 614.730 1712.020 614.875 ;
        RECT 1798.700 614.730 1798.960 614.875 ;
        RECT 1801.920 614.730 1802.180 614.875 ;
        RECT 1895.360 613.205 1895.500 614.875 ;
        RECT 1946.420 614.710 1946.560 615.555 ;
        RECT 2028.300 615.245 2028.440 616.915 ;
        RECT 2052.610 616.235 2052.890 616.605 ;
        RECT 2028.230 614.875 2028.510 615.245 ;
        RECT 1932.100 614.565 1932.360 614.710 ;
        RECT 1932.090 614.195 1932.370 614.565 ;
        RECT 1946.360 614.390 1946.620 614.710 ;
        RECT 2052.680 614.565 2052.820 616.235 ;
        RECT 2124.830 615.555 2125.110 615.925 ;
        RECT 2124.900 615.390 2125.040 615.555 ;
        RECT 2090.340 615.245 2090.600 615.390 ;
        RECT 2090.330 614.875 2090.610 615.245 ;
        RECT 2124.840 615.070 2125.100 615.390 ;
        RECT 2052.610 614.195 2052.890 614.565 ;
        RECT 1895.290 612.835 1895.570 613.205 ;
      LAYER via2 ;
        RECT 1206.210 2497.840 1206.490 2498.120 ;
        RECT 2028.230 616.960 2028.510 617.240 ;
        RECT 1352.030 615.600 1352.310 615.880 ;
        RECT 1946.350 615.600 1946.630 615.880 ;
        RECT 1386.530 614.920 1386.810 615.200 ;
        RECT 1593.990 614.920 1594.270 615.200 ;
        RECT 1607.790 614.920 1608.070 615.200 ;
        RECT 1702.090 614.920 1702.370 615.200 ;
        RECT 1711.750 614.920 1712.030 615.200 ;
        RECT 1798.690 614.920 1798.970 615.200 ;
        RECT 1801.910 614.920 1802.190 615.200 ;
        RECT 1895.290 614.920 1895.570 615.200 ;
        RECT 2052.610 616.280 2052.890 616.560 ;
        RECT 2028.230 614.920 2028.510 615.200 ;
        RECT 1932.090 614.240 1932.370 614.520 ;
        RECT 2124.830 615.600 2125.110 615.880 ;
        RECT 2090.330 614.920 2090.610 615.200 ;
        RECT 2052.610 614.240 2052.890 614.520 ;
        RECT 1895.290 612.880 1895.570 613.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 615.140 2924.800 616.340 ;
=======
        RECT 1206.185 2498.140 1206.515 2498.145 ;
        RECT 1206.185 2498.130 1206.770 2498.140 ;
        RECT 1206.185 2497.830 1206.970 2498.130 ;
        RECT 1206.185 2497.820 1206.770 2497.830 ;
        RECT 1206.185 2497.815 1206.515 2497.820 ;
        RECT 1980.110 617.250 1980.490 617.260 ;
        RECT 2028.205 617.250 2028.535 617.265 ;
        RECT 1980.110 616.950 2028.535 617.250 ;
        RECT 1980.110 616.940 1980.490 616.950 ;
        RECT 2028.205 616.935 2028.535 616.950 ;
        RECT 2052.585 616.570 2052.915 616.585 ;
        RECT 2028.910 616.270 2052.915 616.570 ;
        RECT 1352.005 615.890 1352.335 615.905 ;
        RECT 1946.325 615.890 1946.655 615.905 ;
        RECT 1980.110 615.890 1980.490 615.900 ;
        RECT 1274.510 615.720 1296.890 615.890 ;
        RECT 1297.510 615.720 1317.130 615.890 ;
        RECT 1318.670 615.720 1352.335 615.890 ;
        RECT 1274.510 615.590 1352.335 615.720 ;
        RECT 1206.390 615.210 1206.770 615.220 ;
        RECT 1274.510 615.210 1274.810 615.590 ;
        RECT 1296.590 615.420 1297.810 615.590 ;
        RECT 1316.830 615.420 1318.970 615.590 ;
        RECT 1352.005 615.575 1352.335 615.590 ;
        RECT 1463.110 615.590 1511.250 615.890 ;
        RECT 1206.390 614.910 1274.810 615.210 ;
        RECT 1386.505 615.210 1386.835 615.225 ;
        RECT 1463.110 615.210 1463.410 615.590 ;
        RECT 1386.505 614.910 1463.410 615.210 ;
        RECT 1206.390 614.900 1206.770 614.910 ;
        RECT 1386.505 614.895 1386.835 614.910 ;
        RECT 1510.950 614.530 1511.250 615.590 ;
        RECT 1946.325 615.590 1980.490 615.890 ;
        RECT 1946.325 615.575 1946.655 615.590 ;
        RECT 1980.110 615.580 1980.490 615.590 ;
        RECT 1593.965 615.210 1594.295 615.225 ;
        RECT 1559.710 614.910 1594.295 615.210 ;
        RECT 1559.710 614.530 1560.010 614.910 ;
        RECT 1593.965 614.895 1594.295 614.910 ;
        RECT 1607.765 615.210 1608.095 615.225 ;
        RECT 1702.065 615.210 1702.395 615.225 ;
        RECT 1607.765 614.910 1641.890 615.210 ;
        RECT 1607.765 614.895 1608.095 614.910 ;
        RECT 1510.950 614.230 1560.010 614.530 ;
        RECT 1641.590 614.530 1641.890 614.910 ;
        RECT 1656.310 614.910 1702.395 615.210 ;
        RECT 1656.310 614.530 1656.610 614.910 ;
        RECT 1702.065 614.895 1702.395 614.910 ;
        RECT 1711.725 615.210 1712.055 615.225 ;
        RECT 1798.665 615.210 1798.995 615.225 ;
        RECT 1711.725 614.910 1738.490 615.210 ;
        RECT 1711.725 614.895 1712.055 614.910 ;
        RECT 1641.590 614.230 1656.610 614.530 ;
        RECT 1738.190 614.530 1738.490 614.910 ;
        RECT 1752.910 614.910 1798.995 615.210 ;
        RECT 1752.910 614.530 1753.210 614.910 ;
        RECT 1798.665 614.895 1798.995 614.910 ;
        RECT 1801.885 615.210 1802.215 615.225 ;
        RECT 1895.265 615.210 1895.595 615.225 ;
        RECT 1801.885 614.910 1835.090 615.210 ;
        RECT 1801.885 614.895 1802.215 614.910 ;
        RECT 1738.190 614.230 1753.210 614.530 ;
        RECT 1834.790 614.530 1835.090 614.910 ;
        RECT 1849.510 614.910 1895.595 615.210 ;
        RECT 1849.510 614.530 1849.810 614.910 ;
        RECT 1895.265 614.895 1895.595 614.910 ;
        RECT 2028.205 615.210 2028.535 615.225 ;
        RECT 2028.910 615.210 2029.210 616.270 ;
        RECT 2052.585 616.255 2052.915 616.270 ;
        RECT 2124.805 615.890 2125.135 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2124.805 615.590 2159.850 615.890 ;
        RECT 2124.805 615.575 2125.135 615.590 ;
        RECT 2090.305 615.210 2090.635 615.225 ;
        RECT 2028.205 614.910 2029.210 615.210 ;
        RECT 2076.750 614.910 2090.635 615.210 ;
        RECT 2159.550 615.210 2159.850 615.590 ;
        RECT 2208.310 615.590 2256.450 615.890 ;
        RECT 2159.550 614.910 2207.690 615.210 ;
        RECT 2028.205 614.895 2028.535 614.910 ;
        RECT 1932.065 614.530 1932.395 614.545 ;
        RECT 1834.790 614.230 1849.810 614.530 ;
        RECT 1931.390 614.230 1932.395 614.530 ;
        RECT 1895.265 613.170 1895.595 613.185 ;
        RECT 1931.390 613.170 1931.690 614.230 ;
        RECT 1932.065 614.215 1932.395 614.230 ;
        RECT 2052.585 614.530 2052.915 614.545 ;
        RECT 2076.750 614.530 2077.050 614.910 ;
        RECT 2090.305 614.895 2090.635 614.910 ;
        RECT 2052.585 614.230 2077.050 614.530 ;
        RECT 2207.390 614.530 2207.690 614.910 ;
        RECT 2208.310 614.530 2208.610 615.590 ;
        RECT 2256.150 615.210 2256.450 615.590 ;
        RECT 2304.910 615.590 2353.050 615.890 ;
        RECT 2256.150 614.910 2304.290 615.210 ;
        RECT 2207.390 614.230 2208.610 614.530 ;
        RECT 2303.990 614.530 2304.290 614.910 ;
        RECT 2304.910 614.530 2305.210 615.590 ;
        RECT 2352.750 615.210 2353.050 615.590 ;
        RECT 2401.510 615.590 2449.650 615.890 ;
        RECT 2352.750 614.910 2400.890 615.210 ;
        RECT 2303.990 614.230 2305.210 614.530 ;
        RECT 2400.590 614.530 2400.890 614.910 ;
        RECT 2401.510 614.530 2401.810 615.590 ;
        RECT 2449.350 615.210 2449.650 615.590 ;
        RECT 2498.110 615.590 2546.250 615.890 ;
        RECT 2449.350 614.910 2497.490 615.210 ;
        RECT 2400.590 614.230 2401.810 614.530 ;
        RECT 2497.190 614.530 2497.490 614.910 ;
        RECT 2498.110 614.530 2498.410 615.590 ;
        RECT 2545.950 615.210 2546.250 615.590 ;
        RECT 2594.710 615.590 2642.850 615.890 ;
        RECT 2545.950 614.910 2594.090 615.210 ;
        RECT 2497.190 614.230 2498.410 614.530 ;
        RECT 2593.790 614.530 2594.090 614.910 ;
        RECT 2594.710 614.530 2595.010 615.590 ;
        RECT 2642.550 615.210 2642.850 615.590 ;
        RECT 2691.310 615.590 2739.450 615.890 ;
        RECT 2642.550 614.910 2690.690 615.210 ;
        RECT 2593.790 614.230 2595.010 614.530 ;
        RECT 2690.390 614.530 2690.690 614.910 ;
        RECT 2691.310 614.530 2691.610 615.590 ;
        RECT 2739.150 615.210 2739.450 615.590 ;
        RECT 2787.910 615.590 2836.050 615.890 ;
        RECT 2739.150 614.910 2787.290 615.210 ;
        RECT 2690.390 614.230 2691.610 614.530 ;
        RECT 2786.990 614.530 2787.290 614.910 ;
        RECT 2787.910 614.530 2788.210 615.590 ;
        RECT 2835.750 615.210 2836.050 615.590 ;
        RECT 2916.710 615.590 2924.800 615.890 ;
        RECT 2916.710 615.210 2917.010 615.590 ;
        RECT 2835.750 614.910 2883.890 615.210 ;
        RECT 2786.990 614.230 2788.210 614.530 ;
        RECT 2883.590 614.530 2883.890 614.910 ;
        RECT 2884.510 614.910 2917.010 615.210 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
        RECT 2884.510 614.530 2884.810 614.910 ;
        RECT 2883.590 614.230 2884.810 614.530 ;
        RECT 2052.585 614.215 2052.915 614.230 ;
        RECT 1895.265 612.870 1931.690 613.170 ;
        RECT 1895.265 612.855 1895.595 612.870 ;
      LAYER via3 ;
        RECT 1206.420 2497.820 1206.740 2498.140 ;
        RECT 1980.140 616.940 1980.460 617.260 ;
        RECT 1206.420 614.900 1206.740 615.220 ;
        RECT 1980.140 615.580 1980.460 615.900 ;
      LAYER met4 ;
        RECT 1206.415 2497.815 1206.745 2498.145 ;
        RECT 1206.430 615.225 1206.730 2497.815 ;
        RECT 1980.135 616.935 1980.465 617.265 ;
        RECT 1980.150 615.905 1980.450 616.935 ;
        RECT 1980.135 615.575 1980.465 615.905 ;
        RECT 1206.415 614.895 1206.745 615.225 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23.530 2500.600 23.850 2500.660 ;
        RECT 1761.410 2500.600 1761.730 2500.660 ;
        RECT 23.530 2500.460 1761.730 2500.600 ;
        RECT 23.530 2500.400 23.850 2500.460 ;
        RECT 1761.410 2500.400 1761.730 2500.460 ;
        RECT 13.870 1621.020 14.190 1621.080 ;
        RECT 23.530 1621.020 23.850 1621.080 ;
        RECT 13.870 1620.880 23.850 1621.020 ;
        RECT 13.870 1620.820 14.190 1620.880 ;
        RECT 23.530 1620.820 23.850 1620.880 ;
      LAYER via ;
        RECT 23.560 2500.400 23.820 2500.660 ;
        RECT 1761.440 2500.400 1761.700 2500.660 ;
        RECT 13.900 1620.820 14.160 1621.080 ;
        RECT 23.560 1620.820 23.820 1621.080 ;
      LAYER met2 ;
        RECT 23.560 2500.370 23.820 2500.690 ;
        RECT 1761.440 2500.370 1761.700 2500.690 ;
        RECT 23.620 1621.110 23.760 2500.370 ;
        RECT 1761.500 2500.000 1761.640 2500.370 ;
        RECT 1761.430 2496.000 1761.710 2500.000 ;
        RECT 13.900 1620.790 14.160 1621.110 ;
        RECT 23.560 1620.790 23.820 1621.110 ;
        RECT 13.960 1615.525 14.100 1620.790 ;
        RECT 13.890 1615.155 14.170 1615.525 ;
      LAYER via2 ;
        RECT 13.890 1615.200 14.170 1615.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1614.740 0.300 1615.940 ;
=======
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 13.865 1615.490 14.195 1615.505 ;
        RECT -4.800 1615.190 14.195 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 13.865 1615.175 14.195 1615.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 27.210 2500.260 27.530 2500.320 ;
        RECT 1780.270 2500.260 1780.590 2500.320 ;
        RECT 27.210 2500.120 1780.590 2500.260 ;
        RECT 27.210 2500.060 27.530 2500.120 ;
        RECT 1780.270 2500.060 1780.590 2500.120 ;
        RECT 13.870 1400.700 14.190 1400.760 ;
        RECT 27.210 1400.700 27.530 1400.760 ;
        RECT 13.870 1400.560 27.530 1400.700 ;
        RECT 13.870 1400.500 14.190 1400.560 ;
        RECT 27.210 1400.500 27.530 1400.560 ;
      LAYER via ;
        RECT 27.240 2500.060 27.500 2500.320 ;
        RECT 1780.300 2500.060 1780.560 2500.320 ;
        RECT 13.900 1400.500 14.160 1400.760 ;
        RECT 27.240 1400.500 27.500 1400.760 ;
      LAYER met2 ;
        RECT 27.240 2500.030 27.500 2500.350 ;
        RECT 1780.300 2500.030 1780.560 2500.350 ;
        RECT 27.300 1400.790 27.440 2500.030 ;
        RECT 1780.360 2499.410 1780.500 2500.030 ;
        RECT 1781.210 2499.410 1781.490 2500.000 ;
        RECT 1780.360 2499.270 1781.490 2499.410 ;
        RECT 1781.210 2496.000 1781.490 2499.270 ;
        RECT 13.900 1400.645 14.160 1400.790 ;
        RECT 13.890 1400.275 14.170 1400.645 ;
        RECT 27.240 1400.470 27.500 1400.790 ;
      LAYER via2 ;
        RECT 13.890 1400.320 14.170 1400.600 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1399.860 0.300 1401.060 ;
=======
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 13.865 1400.610 14.195 1400.625 ;
        RECT -4.800 1400.310 14.195 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 13.865 1400.295 14.195 1400.310 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 26.290 2499.920 26.610 2499.980 ;
        RECT 1800.510 2499.920 1800.830 2499.980 ;
        RECT 26.290 2499.780 1800.830 2499.920 ;
        RECT 26.290 2499.720 26.610 2499.780 ;
        RECT 1800.510 2499.720 1800.830 2499.780 ;
        RECT 13.870 1186.500 14.190 1186.560 ;
        RECT 26.290 1186.500 26.610 1186.560 ;
        RECT 13.870 1186.360 26.610 1186.500 ;
        RECT 13.870 1186.300 14.190 1186.360 ;
        RECT 26.290 1186.300 26.610 1186.360 ;
      LAYER via ;
        RECT 26.320 2499.720 26.580 2499.980 ;
        RECT 1800.540 2499.720 1800.800 2499.980 ;
        RECT 13.900 1186.300 14.160 1186.560 ;
        RECT 26.320 1186.300 26.580 1186.560 ;
      LAYER met2 ;
        RECT 26.320 2499.690 26.580 2500.010 ;
        RECT 1800.540 2499.690 1800.800 2500.010 ;
        RECT 26.380 1186.590 26.520 2499.690 ;
        RECT 1800.600 2499.410 1800.740 2499.690 ;
        RECT 1800.990 2499.410 1801.270 2500.000 ;
        RECT 1800.600 2499.270 1801.270 2499.410 ;
        RECT 1800.990 2496.000 1801.270 2499.270 ;
        RECT 13.900 1186.270 14.160 1186.590 ;
        RECT 26.320 1186.270 26.580 1186.590 ;
        RECT 13.960 1185.085 14.100 1186.270 ;
        RECT 13.890 1184.715 14.170 1185.085 ;
      LAYER via2 ;
        RECT 13.890 1184.760 14.170 1185.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1184.300 0.300 1185.500 ;
=======
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 13.865 1185.050 14.195 1185.065 ;
        RECT -4.800 1184.750 14.195 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 13.865 1184.735 14.195 1184.750 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 31.810 2499.580 32.130 2499.640 ;
        RECT 1818.910 2499.580 1819.230 2499.640 ;
        RECT 31.810 2499.440 1819.230 2499.580 ;
        RECT 31.810 2499.380 32.130 2499.440 ;
        RECT 1818.910 2499.380 1819.230 2499.440 ;
        RECT 16.170 971.620 16.490 971.680 ;
        RECT 31.810 971.620 32.130 971.680 ;
        RECT 16.170 971.480 32.130 971.620 ;
        RECT 16.170 971.420 16.490 971.480 ;
        RECT 31.810 971.420 32.130 971.480 ;
      LAYER via ;
        RECT 31.840 2499.380 32.100 2499.640 ;
        RECT 1818.940 2499.380 1819.200 2499.640 ;
        RECT 16.200 971.420 16.460 971.680 ;
        RECT 31.840 971.420 32.100 971.680 ;
      LAYER met2 ;
        RECT 31.840 2499.350 32.100 2499.670 ;
        RECT 1818.940 2499.410 1819.200 2499.670 ;
        RECT 1820.770 2499.410 1821.050 2500.000 ;
        RECT 1818.940 2499.350 1821.050 2499.410 ;
        RECT 31.900 971.710 32.040 2499.350 ;
        RECT 1819.000 2499.270 1821.050 2499.350 ;
        RECT 1820.770 2496.000 1821.050 2499.270 ;
        RECT 16.200 971.390 16.460 971.710 ;
        RECT 31.840 971.390 32.100 971.710 ;
        RECT 16.260 969.525 16.400 971.390 ;
        RECT 16.190 969.155 16.470 969.525 ;
      LAYER via2 ;
        RECT 16.190 969.200 16.470 969.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 968.740 0.300 969.940 ;
=======
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 16.165 969.490 16.495 969.505 ;
        RECT -4.800 969.190 16.495 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 16.165 969.175 16.495 969.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.910 2499.240 25.230 2499.300 ;
        RECT 1839.150 2499.240 1839.470 2499.300 ;
        RECT 24.910 2499.100 1839.470 2499.240 ;
        RECT 24.910 2499.040 25.230 2499.100 ;
        RECT 1839.150 2499.040 1839.470 2499.100 ;
        RECT 13.870 756.060 14.190 756.120 ;
        RECT 24.910 756.060 25.230 756.120 ;
        RECT 13.870 755.920 25.230 756.060 ;
        RECT 13.870 755.860 14.190 755.920 ;
        RECT 24.910 755.860 25.230 755.920 ;
      LAYER via ;
        RECT 24.940 2499.040 25.200 2499.300 ;
        RECT 1839.180 2499.040 1839.440 2499.300 ;
        RECT 13.900 755.860 14.160 756.120 ;
        RECT 24.940 755.860 25.200 756.120 ;
      LAYER met2 ;
        RECT 1840.550 2499.410 1840.830 2500.000 ;
        RECT 1839.240 2499.330 1840.830 2499.410 ;
        RECT 24.940 2499.010 25.200 2499.330 ;
        RECT 1839.180 2499.270 1840.830 2499.330 ;
        RECT 1839.180 2499.010 1839.440 2499.270 ;
        RECT 25.000 756.150 25.140 2499.010 ;
        RECT 1840.550 2496.000 1840.830 2499.270 ;
        RECT 13.900 755.830 14.160 756.150 ;
        RECT 24.940 755.830 25.200 756.150 ;
        RECT 13.960 753.965 14.100 755.830 ;
        RECT 13.890 753.595 14.170 753.965 ;
      LAYER via2 ;
        RECT 13.890 753.640 14.170 753.920 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 753.180 0.300 754.380 ;
=======
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 13.865 753.930 14.195 753.945 ;
        RECT -4.800 753.630 14.195 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 13.865 753.615 14.195 753.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2498.900 17.870 2498.960 ;
        RECT 1858.470 2498.900 1858.790 2498.960 ;
        RECT 17.550 2498.760 1858.790 2498.900 ;
        RECT 17.550 2498.700 17.870 2498.760 ;
        RECT 1858.470 2498.700 1858.790 2498.760 ;
      LAYER via ;
        RECT 17.580 2498.700 17.840 2498.960 ;
        RECT 1858.500 2498.700 1858.760 2498.960 ;
      LAYER met2 ;
        RECT 17.580 2498.670 17.840 2498.990 ;
        RECT 1858.500 2498.730 1858.760 2498.990 ;
        RECT 1860.330 2498.730 1860.610 2500.000 ;
        RECT 1858.500 2498.670 1860.610 2498.730 ;
        RECT 17.640 538.405 17.780 2498.670 ;
        RECT 1858.560 2498.590 1860.610 2498.670 ;
        RECT 1860.330 2496.000 1860.610 2498.590 ;
        RECT 17.570 538.035 17.850 538.405 ;
      LAYER via2 ;
        RECT 17.570 538.080 17.850 538.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 537.620 0.300 538.820 ;
=======
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 17.545 538.370 17.875 538.385 ;
        RECT -4.800 538.070 17.875 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 17.545 538.055 17.875 538.070 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 31.350 2498.560 31.670 2498.620 ;
        RECT 1878.710 2498.560 1879.030 2498.620 ;
        RECT 31.350 2498.420 1879.030 2498.560 ;
        RECT 31.350 2498.360 31.670 2498.420 ;
        RECT 1878.710 2498.360 1879.030 2498.420 ;
        RECT 15.710 323.580 16.030 323.640 ;
        RECT 31.350 323.580 31.670 323.640 ;
        RECT 15.710 323.440 31.670 323.580 ;
        RECT 15.710 323.380 16.030 323.440 ;
        RECT 31.350 323.380 31.670 323.440 ;
      LAYER via ;
        RECT 31.380 2498.360 31.640 2498.620 ;
        RECT 1878.740 2498.360 1879.000 2498.620 ;
        RECT 15.740 323.380 16.000 323.640 ;
        RECT 31.380 323.380 31.640 323.640 ;
      LAYER met2 ;
        RECT 1880.110 2498.730 1880.390 2500.000 ;
        RECT 1878.800 2498.650 1880.390 2498.730 ;
        RECT 31.380 2498.330 31.640 2498.650 ;
        RECT 1878.740 2498.590 1880.390 2498.650 ;
        RECT 1878.740 2498.330 1879.000 2498.590 ;
        RECT 31.440 323.670 31.580 2498.330 ;
        RECT 1880.110 2496.000 1880.390 2498.590 ;
        RECT 15.740 323.350 16.000 323.670 ;
        RECT 31.380 323.350 31.640 323.670 ;
        RECT 15.800 322.845 15.940 323.350 ;
        RECT 15.730 322.475 16.010 322.845 ;
      LAYER via2 ;
        RECT 15.730 322.520 16.010 322.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 322.060 0.300 323.260 ;
=======
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 15.705 322.810 16.035 322.825 ;
        RECT -4.800 322.510 16.035 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 15.705 322.495 16.035 322.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.890 2497.880 31.210 2497.940 ;
        RECT 1898.950 2497.880 1899.270 2497.940 ;
        RECT 30.890 2497.740 1899.270 2497.880 ;
        RECT 30.890 2497.680 31.210 2497.740 ;
        RECT 1898.950 2497.680 1899.270 2497.740 ;
        RECT 14.790 109.040 15.110 109.100 ;
        RECT 30.890 109.040 31.210 109.100 ;
        RECT 14.790 108.900 31.210 109.040 ;
        RECT 14.790 108.840 15.110 108.900 ;
        RECT 30.890 108.840 31.210 108.900 ;
      LAYER via ;
        RECT 30.920 2497.680 31.180 2497.940 ;
        RECT 1898.980 2497.680 1899.240 2497.940 ;
        RECT 14.820 108.840 15.080 109.100 ;
        RECT 30.920 108.840 31.180 109.100 ;
      LAYER met2 ;
        RECT 1900.350 2498.050 1900.630 2500.000 ;
        RECT 1899.040 2497.970 1900.630 2498.050 ;
        RECT 30.920 2497.650 31.180 2497.970 ;
        RECT 1898.980 2497.910 1900.630 2497.970 ;
        RECT 1898.980 2497.650 1899.240 2497.910 ;
        RECT 30.980 109.130 31.120 2497.650 ;
        RECT 1900.350 2496.000 1900.630 2497.910 ;
        RECT 14.820 108.810 15.080 109.130 ;
        RECT 30.920 108.810 31.180 109.130 ;
        RECT 14.880 107.285 15.020 108.810 ;
        RECT 14.810 106.915 15.090 107.285 ;
      LAYER via2 ;
        RECT 14.810 106.960 15.090 107.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 106.500 0.300 107.700 ;
=======
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 14.785 107.250 15.115 107.265 ;
        RECT -4.800 106.950 15.115 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 14.785 106.935 15.115 106.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2090.310 849.900 2090.630 849.960 ;
        RECT 2124.810 849.900 2125.130 849.960 ;
        RECT 2090.310 849.760 2125.130 849.900 ;
        RECT 2090.310 849.700 2090.630 849.760 ;
        RECT 2124.810 849.700 2125.130 849.760 ;
        RECT 1606.390 849.560 1606.710 849.620 ;
        RECT 1607.770 849.560 1608.090 849.620 ;
        RECT 1606.390 849.420 1608.090 849.560 ;
        RECT 1606.390 849.360 1606.710 849.420 ;
        RECT 1607.770 849.360 1608.090 849.420 ;
        RECT 1702.070 849.560 1702.390 849.620 ;
        RECT 1711.730 849.560 1712.050 849.620 ;
        RECT 1702.070 849.420 1712.050 849.560 ;
        RECT 1702.070 849.360 1702.390 849.420 ;
        RECT 1711.730 849.360 1712.050 849.420 ;
        RECT 1798.670 849.560 1798.990 849.620 ;
        RECT 1801.890 849.560 1802.210 849.620 ;
        RECT 1798.670 849.420 1802.210 849.560 ;
        RECT 1798.670 849.360 1798.990 849.420 ;
        RECT 1801.890 849.360 1802.210 849.420 ;
        RECT 1932.070 849.220 1932.390 849.280 ;
        RECT 1946.330 849.220 1946.650 849.280 ;
        RECT 1932.070 849.080 1946.650 849.220 ;
        RECT 1932.070 849.020 1932.390 849.080 ;
        RECT 1946.330 849.020 1946.650 849.080 ;
      LAYER via ;
        RECT 2090.340 849.700 2090.600 849.960 ;
        RECT 2124.840 849.700 2125.100 849.960 ;
        RECT 1606.420 849.360 1606.680 849.620 ;
        RECT 1607.800 849.360 1608.060 849.620 ;
        RECT 1702.100 849.360 1702.360 849.620 ;
        RECT 1711.760 849.360 1712.020 849.620 ;
        RECT 1798.700 849.360 1798.960 849.620 ;
        RECT 1801.920 849.360 1802.180 849.620 ;
        RECT 1932.100 849.020 1932.360 849.280 ;
        RECT 1946.360 849.020 1946.620 849.280 ;
      LAYER met2 ;
        RECT 1225.990 2498.050 1226.270 2500.000 ;
        RECT 1226.450 2498.050 1226.730 2498.165 ;
        RECT 1225.990 2497.910 1226.730 2498.050 ;
        RECT 1225.990 2496.000 1226.270 2497.910 ;
        RECT 1226.450 2497.795 1226.730 2497.910 ;
        RECT 1255.430 859.675 1255.710 860.045 ;
        RECT 1255.500 849.845 1255.640 859.675 ;
        RECT 2028.230 851.515 2028.510 851.885 ;
        RECT 1325.350 850.835 1325.630 851.205 ;
        RECT 1490.030 850.835 1490.310 851.205 ;
        RECT 1325.420 849.845 1325.560 850.835 ;
        RECT 1255.430 849.475 1255.710 849.845 ;
        RECT 1325.350 849.475 1325.630 849.845 ;
        RECT 1490.100 849.165 1490.240 850.835 ;
        RECT 1496.930 850.155 1497.210 850.525 ;
        RECT 1946.350 850.155 1946.630 850.525 ;
        RECT 1497.000 849.165 1497.140 850.155 ;
        RECT 1606.410 849.475 1606.690 849.845 ;
        RECT 1607.790 849.475 1608.070 849.845 ;
        RECT 1702.090 849.475 1702.370 849.845 ;
        RECT 1711.750 849.475 1712.030 849.845 ;
        RECT 1798.690 849.475 1798.970 849.845 ;
        RECT 1801.910 849.475 1802.190 849.845 ;
        RECT 1895.290 849.475 1895.570 849.845 ;
        RECT 1606.420 849.330 1606.680 849.475 ;
        RECT 1607.800 849.330 1608.060 849.475 ;
        RECT 1702.100 849.330 1702.360 849.475 ;
        RECT 1711.760 849.330 1712.020 849.475 ;
        RECT 1798.700 849.330 1798.960 849.475 ;
        RECT 1801.920 849.330 1802.180 849.475 ;
        RECT 1490.030 848.795 1490.310 849.165 ;
        RECT 1496.930 848.795 1497.210 849.165 ;
        RECT 1895.360 847.805 1895.500 849.475 ;
        RECT 1946.420 849.310 1946.560 850.155 ;
        RECT 2028.300 849.845 2028.440 851.515 ;
        RECT 2052.610 850.835 2052.890 851.205 ;
        RECT 2028.230 849.475 2028.510 849.845 ;
        RECT 1932.100 849.165 1932.360 849.310 ;
        RECT 1932.090 848.795 1932.370 849.165 ;
        RECT 1946.360 848.990 1946.620 849.310 ;
        RECT 2052.680 849.165 2052.820 850.835 ;
        RECT 2124.830 850.155 2125.110 850.525 ;
        RECT 2124.900 849.990 2125.040 850.155 ;
        RECT 2090.340 849.845 2090.600 849.990 ;
        RECT 2090.330 849.475 2090.610 849.845 ;
        RECT 2124.840 849.670 2125.100 849.990 ;
        RECT 2052.610 848.795 2052.890 849.165 ;
        RECT 1895.290 847.435 1895.570 847.805 ;
      LAYER via2 ;
        RECT 1226.450 2497.840 1226.730 2498.120 ;
        RECT 1255.430 859.720 1255.710 860.000 ;
        RECT 2028.230 851.560 2028.510 851.840 ;
        RECT 1325.350 850.880 1325.630 851.160 ;
        RECT 1490.030 850.880 1490.310 851.160 ;
        RECT 1255.430 849.520 1255.710 849.800 ;
        RECT 1325.350 849.520 1325.630 849.800 ;
        RECT 1496.930 850.200 1497.210 850.480 ;
        RECT 1946.350 850.200 1946.630 850.480 ;
        RECT 1606.410 849.520 1606.690 849.800 ;
        RECT 1607.790 849.520 1608.070 849.800 ;
        RECT 1702.090 849.520 1702.370 849.800 ;
        RECT 1711.750 849.520 1712.030 849.800 ;
        RECT 1798.690 849.520 1798.970 849.800 ;
        RECT 1801.910 849.520 1802.190 849.800 ;
        RECT 1895.290 849.520 1895.570 849.800 ;
        RECT 1490.030 848.840 1490.310 849.120 ;
        RECT 1496.930 848.840 1497.210 849.120 ;
        RECT 2052.610 850.880 2052.890 851.160 ;
        RECT 2028.230 849.520 2028.510 849.800 ;
        RECT 1932.090 848.840 1932.370 849.120 ;
        RECT 2124.830 850.200 2125.110 850.480 ;
        RECT 2090.330 849.520 2090.610 849.800 ;
        RECT 2052.610 848.840 2052.890 849.120 ;
        RECT 1895.290 847.480 1895.570 847.760 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 849.740 2924.800 850.940 ;
=======
        RECT 1226.425 2498.140 1226.755 2498.145 ;
        RECT 1226.425 2498.130 1227.010 2498.140 ;
        RECT 1226.425 2497.830 1227.210 2498.130 ;
        RECT 1226.425 2497.820 1227.010 2497.830 ;
        RECT 1226.425 2497.815 1226.755 2497.820 ;
        RECT 1226.630 860.010 1227.010 860.020 ;
        RECT 1255.405 860.010 1255.735 860.025 ;
        RECT 1226.630 859.710 1255.735 860.010 ;
        RECT 1226.630 859.700 1227.010 859.710 ;
        RECT 1255.405 859.695 1255.735 859.710 ;
        RECT 1980.110 851.850 1980.490 851.860 ;
        RECT 2028.205 851.850 2028.535 851.865 ;
        RECT 1980.110 851.550 2028.535 851.850 ;
        RECT 1980.110 851.540 1980.490 851.550 ;
        RECT 2028.205 851.535 2028.535 851.550 ;
        RECT 1325.325 851.170 1325.655 851.185 ;
        RECT 1345.310 851.170 1345.690 851.180 ;
        RECT 1325.325 850.870 1345.690 851.170 ;
        RECT 1325.325 850.855 1325.655 850.870 ;
        RECT 1345.310 850.860 1345.690 850.870 ;
        RECT 1441.910 851.170 1442.290 851.180 ;
        RECT 1490.005 851.170 1490.335 851.185 ;
        RECT 2052.585 851.170 2052.915 851.185 ;
        RECT 1441.910 850.870 1490.335 851.170 ;
        RECT 1441.910 850.860 1442.290 850.870 ;
        RECT 1490.005 850.855 1490.335 850.870 ;
        RECT 2028.910 850.870 2052.915 851.170 ;
        RECT 1496.905 850.490 1497.235 850.505 ;
        RECT 1946.325 850.490 1946.655 850.505 ;
        RECT 1980.110 850.490 1980.490 850.500 ;
        RECT 1496.905 850.175 1497.450 850.490 ;
        RECT 1946.325 850.190 1980.490 850.490 ;
        RECT 1946.325 850.175 1946.655 850.190 ;
        RECT 1980.110 850.180 1980.490 850.190 ;
        RECT 1255.405 849.810 1255.735 849.825 ;
        RECT 1325.325 849.810 1325.655 849.825 ;
        RECT 1255.405 849.510 1325.655 849.810 ;
        RECT 1255.405 849.495 1255.735 849.510 ;
        RECT 1325.325 849.495 1325.655 849.510 ;
        RECT 1345.310 849.810 1345.690 849.820 ;
        RECT 1441.910 849.810 1442.290 849.820 ;
        RECT 1345.310 849.510 1442.290 849.810 ;
        RECT 1497.150 849.810 1497.450 850.175 ;
        RECT 1606.385 849.810 1606.715 849.825 ;
        RECT 1497.150 849.510 1545.290 849.810 ;
        RECT 1345.310 849.500 1345.690 849.510 ;
        RECT 1441.910 849.500 1442.290 849.510 ;
        RECT 1490.005 849.130 1490.335 849.145 ;
        RECT 1496.905 849.130 1497.235 849.145 ;
        RECT 1490.005 848.830 1497.235 849.130 ;
        RECT 1544.990 849.130 1545.290 849.510 ;
        RECT 1559.710 849.510 1606.715 849.810 ;
        RECT 1559.710 849.130 1560.010 849.510 ;
        RECT 1606.385 849.495 1606.715 849.510 ;
        RECT 1607.765 849.810 1608.095 849.825 ;
        RECT 1702.065 849.810 1702.395 849.825 ;
        RECT 1607.765 849.510 1641.890 849.810 ;
        RECT 1607.765 849.495 1608.095 849.510 ;
        RECT 1544.990 848.830 1560.010 849.130 ;
        RECT 1641.590 849.130 1641.890 849.510 ;
        RECT 1656.310 849.510 1702.395 849.810 ;
        RECT 1656.310 849.130 1656.610 849.510 ;
        RECT 1702.065 849.495 1702.395 849.510 ;
        RECT 1711.725 849.810 1712.055 849.825 ;
        RECT 1798.665 849.810 1798.995 849.825 ;
        RECT 1711.725 849.510 1738.490 849.810 ;
        RECT 1711.725 849.495 1712.055 849.510 ;
        RECT 1641.590 848.830 1656.610 849.130 ;
        RECT 1738.190 849.130 1738.490 849.510 ;
        RECT 1752.910 849.510 1798.995 849.810 ;
        RECT 1752.910 849.130 1753.210 849.510 ;
        RECT 1798.665 849.495 1798.995 849.510 ;
        RECT 1801.885 849.810 1802.215 849.825 ;
        RECT 1895.265 849.810 1895.595 849.825 ;
        RECT 1801.885 849.510 1835.090 849.810 ;
        RECT 1801.885 849.495 1802.215 849.510 ;
        RECT 1738.190 848.830 1753.210 849.130 ;
        RECT 1834.790 849.130 1835.090 849.510 ;
        RECT 1849.510 849.510 1895.595 849.810 ;
        RECT 1849.510 849.130 1849.810 849.510 ;
        RECT 1895.265 849.495 1895.595 849.510 ;
        RECT 2028.205 849.810 2028.535 849.825 ;
        RECT 2028.910 849.810 2029.210 850.870 ;
        RECT 2052.585 850.855 2052.915 850.870 ;
        RECT 2124.805 850.490 2125.135 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2124.805 850.190 2159.850 850.490 ;
        RECT 2124.805 850.175 2125.135 850.190 ;
        RECT 2090.305 849.810 2090.635 849.825 ;
        RECT 2028.205 849.510 2029.210 849.810 ;
        RECT 2076.750 849.510 2090.635 849.810 ;
        RECT 2159.550 849.810 2159.850 850.190 ;
        RECT 2208.310 850.190 2256.450 850.490 ;
        RECT 2159.550 849.510 2207.690 849.810 ;
        RECT 2028.205 849.495 2028.535 849.510 ;
        RECT 1932.065 849.130 1932.395 849.145 ;
        RECT 1834.790 848.830 1849.810 849.130 ;
        RECT 1931.390 848.830 1932.395 849.130 ;
        RECT 1490.005 848.815 1490.335 848.830 ;
        RECT 1496.905 848.815 1497.235 848.830 ;
        RECT 1895.265 847.770 1895.595 847.785 ;
        RECT 1931.390 847.770 1931.690 848.830 ;
        RECT 1932.065 848.815 1932.395 848.830 ;
        RECT 2052.585 849.130 2052.915 849.145 ;
        RECT 2076.750 849.130 2077.050 849.510 ;
        RECT 2090.305 849.495 2090.635 849.510 ;
        RECT 2052.585 848.830 2077.050 849.130 ;
        RECT 2207.390 849.130 2207.690 849.510 ;
        RECT 2208.310 849.130 2208.610 850.190 ;
        RECT 2256.150 849.810 2256.450 850.190 ;
        RECT 2304.910 850.190 2353.050 850.490 ;
        RECT 2256.150 849.510 2304.290 849.810 ;
        RECT 2207.390 848.830 2208.610 849.130 ;
        RECT 2303.990 849.130 2304.290 849.510 ;
        RECT 2304.910 849.130 2305.210 850.190 ;
        RECT 2352.750 849.810 2353.050 850.190 ;
        RECT 2401.510 850.190 2449.650 850.490 ;
        RECT 2352.750 849.510 2400.890 849.810 ;
        RECT 2303.990 848.830 2305.210 849.130 ;
        RECT 2400.590 849.130 2400.890 849.510 ;
        RECT 2401.510 849.130 2401.810 850.190 ;
        RECT 2449.350 849.810 2449.650 850.190 ;
        RECT 2498.110 850.190 2546.250 850.490 ;
        RECT 2449.350 849.510 2497.490 849.810 ;
        RECT 2400.590 848.830 2401.810 849.130 ;
        RECT 2497.190 849.130 2497.490 849.510 ;
        RECT 2498.110 849.130 2498.410 850.190 ;
        RECT 2545.950 849.810 2546.250 850.190 ;
        RECT 2594.710 850.190 2642.850 850.490 ;
        RECT 2545.950 849.510 2594.090 849.810 ;
        RECT 2497.190 848.830 2498.410 849.130 ;
        RECT 2593.790 849.130 2594.090 849.510 ;
        RECT 2594.710 849.130 2595.010 850.190 ;
        RECT 2642.550 849.810 2642.850 850.190 ;
        RECT 2691.310 850.190 2739.450 850.490 ;
        RECT 2642.550 849.510 2690.690 849.810 ;
        RECT 2593.790 848.830 2595.010 849.130 ;
        RECT 2690.390 849.130 2690.690 849.510 ;
        RECT 2691.310 849.130 2691.610 850.190 ;
        RECT 2739.150 849.810 2739.450 850.190 ;
        RECT 2787.910 850.190 2836.050 850.490 ;
        RECT 2739.150 849.510 2787.290 849.810 ;
        RECT 2690.390 848.830 2691.610 849.130 ;
        RECT 2786.990 849.130 2787.290 849.510 ;
        RECT 2787.910 849.130 2788.210 850.190 ;
        RECT 2835.750 849.810 2836.050 850.190 ;
        RECT 2916.710 850.190 2924.800 850.490 ;
        RECT 2916.710 849.810 2917.010 850.190 ;
        RECT 2835.750 849.510 2883.890 849.810 ;
        RECT 2786.990 848.830 2788.210 849.130 ;
        RECT 2883.590 849.130 2883.890 849.510 ;
        RECT 2884.510 849.510 2917.010 849.810 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
        RECT 2884.510 849.130 2884.810 849.510 ;
        RECT 2883.590 848.830 2884.810 849.130 ;
        RECT 2052.585 848.815 2052.915 848.830 ;
        RECT 1895.265 847.470 1931.690 847.770 ;
        RECT 1895.265 847.455 1895.595 847.470 ;
      LAYER via3 ;
        RECT 1226.660 2497.820 1226.980 2498.140 ;
        RECT 1226.660 859.700 1226.980 860.020 ;
        RECT 1980.140 851.540 1980.460 851.860 ;
        RECT 1345.340 850.860 1345.660 851.180 ;
        RECT 1441.940 850.860 1442.260 851.180 ;
        RECT 1980.140 850.180 1980.460 850.500 ;
        RECT 1345.340 849.500 1345.660 849.820 ;
        RECT 1441.940 849.500 1442.260 849.820 ;
      LAYER met4 ;
        RECT 1226.655 2497.815 1226.985 2498.145 ;
        RECT 1226.670 860.025 1226.970 2497.815 ;
        RECT 1226.655 859.695 1226.985 860.025 ;
        RECT 1980.135 851.535 1980.465 851.865 ;
        RECT 1345.335 850.855 1345.665 851.185 ;
        RECT 1441.935 850.855 1442.265 851.185 ;
        RECT 1345.350 849.825 1345.650 850.855 ;
        RECT 1441.950 849.825 1442.250 850.855 ;
        RECT 1980.150 850.505 1980.450 851.535 ;
        RECT 1980.135 850.175 1980.465 850.505 ;
        RECT 1345.335 849.495 1345.665 849.825 ;
        RECT 1441.935 849.495 1442.265 849.825 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2090.310 1084.500 2090.630 1084.560 ;
        RECT 2124.810 1084.500 2125.130 1084.560 ;
        RECT 2090.310 1084.360 2125.130 1084.500 ;
        RECT 2090.310 1084.300 2090.630 1084.360 ;
        RECT 2124.810 1084.300 2125.130 1084.360 ;
        RECT 1606.390 1084.160 1606.710 1084.220 ;
        RECT 1607.770 1084.160 1608.090 1084.220 ;
        RECT 1606.390 1084.020 1608.090 1084.160 ;
        RECT 1606.390 1083.960 1606.710 1084.020 ;
        RECT 1607.770 1083.960 1608.090 1084.020 ;
        RECT 1702.070 1084.160 1702.390 1084.220 ;
        RECT 1711.730 1084.160 1712.050 1084.220 ;
        RECT 1702.070 1084.020 1712.050 1084.160 ;
        RECT 1702.070 1083.960 1702.390 1084.020 ;
        RECT 1711.730 1083.960 1712.050 1084.020 ;
        RECT 1798.670 1084.160 1798.990 1084.220 ;
        RECT 1801.890 1084.160 1802.210 1084.220 ;
        RECT 1798.670 1084.020 1802.210 1084.160 ;
        RECT 1798.670 1083.960 1798.990 1084.020 ;
        RECT 1801.890 1083.960 1802.210 1084.020 ;
        RECT 1932.070 1083.820 1932.390 1083.880 ;
        RECT 1946.330 1083.820 1946.650 1083.880 ;
        RECT 1932.070 1083.680 1946.650 1083.820 ;
        RECT 1932.070 1083.620 1932.390 1083.680 ;
        RECT 1946.330 1083.620 1946.650 1083.680 ;
      LAYER via ;
        RECT 2090.340 1084.300 2090.600 1084.560 ;
        RECT 2124.840 1084.300 2125.100 1084.560 ;
        RECT 1606.420 1083.960 1606.680 1084.220 ;
        RECT 1607.800 1083.960 1608.060 1084.220 ;
        RECT 1702.100 1083.960 1702.360 1084.220 ;
        RECT 1711.760 1083.960 1712.020 1084.220 ;
        RECT 1798.700 1083.960 1798.960 1084.220 ;
        RECT 1801.920 1083.960 1802.180 1084.220 ;
        RECT 1932.100 1083.620 1932.360 1083.880 ;
        RECT 1946.360 1083.620 1946.620 1083.880 ;
      LAYER met2 ;
        RECT 1245.770 2498.050 1246.050 2500.000 ;
        RECT 1246.690 2498.050 1246.970 2498.165 ;
        RECT 1245.770 2497.910 1246.970 2498.050 ;
        RECT 1245.770 2496.000 1246.050 2497.910 ;
        RECT 1246.690 2497.795 1246.970 2497.910 ;
        RECT 1579.270 1086.115 1579.550 1086.485 ;
        RECT 2028.230 1086.115 2028.510 1086.485 ;
        RECT 1355.710 1084.755 1355.990 1085.125 ;
        RECT 1483.130 1084.755 1483.410 1085.125 ;
        RECT 1355.780 1083.085 1355.920 1084.755 ;
        RECT 1483.200 1084.445 1483.340 1084.755 ;
        RECT 1579.340 1084.445 1579.480 1086.115 ;
        RECT 1946.350 1084.755 1946.630 1085.125 ;
        RECT 1483.130 1084.075 1483.410 1084.445 ;
        RECT 1579.270 1084.075 1579.550 1084.445 ;
        RECT 1606.410 1084.075 1606.690 1084.445 ;
        RECT 1607.790 1084.075 1608.070 1084.445 ;
        RECT 1702.090 1084.075 1702.370 1084.445 ;
        RECT 1711.750 1084.075 1712.030 1084.445 ;
        RECT 1798.690 1084.075 1798.970 1084.445 ;
        RECT 1801.910 1084.075 1802.190 1084.445 ;
        RECT 1895.290 1084.075 1895.570 1084.445 ;
        RECT 1606.420 1083.930 1606.680 1084.075 ;
        RECT 1607.800 1083.930 1608.060 1084.075 ;
        RECT 1702.100 1083.930 1702.360 1084.075 ;
        RECT 1711.760 1083.930 1712.020 1084.075 ;
        RECT 1798.700 1083.930 1798.960 1084.075 ;
        RECT 1801.920 1083.930 1802.180 1084.075 ;
        RECT 1355.710 1082.715 1355.990 1083.085 ;
        RECT 1895.360 1082.405 1895.500 1084.075 ;
        RECT 1946.420 1083.910 1946.560 1084.755 ;
        RECT 2028.300 1084.445 2028.440 1086.115 ;
        RECT 2052.610 1085.435 2052.890 1085.805 ;
        RECT 2028.230 1084.075 2028.510 1084.445 ;
        RECT 1932.100 1083.765 1932.360 1083.910 ;
        RECT 1932.090 1083.395 1932.370 1083.765 ;
        RECT 1946.360 1083.590 1946.620 1083.910 ;
        RECT 2052.680 1083.765 2052.820 1085.435 ;
        RECT 2124.830 1084.755 2125.110 1085.125 ;
        RECT 2124.900 1084.590 2125.040 1084.755 ;
        RECT 2090.340 1084.445 2090.600 1084.590 ;
        RECT 2090.330 1084.075 2090.610 1084.445 ;
        RECT 2124.840 1084.270 2125.100 1084.590 ;
        RECT 2052.610 1083.395 2052.890 1083.765 ;
        RECT 1895.290 1082.035 1895.570 1082.405 ;
      LAYER via2 ;
        RECT 1246.690 2497.840 1246.970 2498.120 ;
        RECT 1579.270 1086.160 1579.550 1086.440 ;
        RECT 2028.230 1086.160 2028.510 1086.440 ;
        RECT 1355.710 1084.800 1355.990 1085.080 ;
        RECT 1483.130 1084.800 1483.410 1085.080 ;
        RECT 1946.350 1084.800 1946.630 1085.080 ;
        RECT 1483.130 1084.120 1483.410 1084.400 ;
        RECT 1579.270 1084.120 1579.550 1084.400 ;
        RECT 1606.410 1084.120 1606.690 1084.400 ;
        RECT 1607.790 1084.120 1608.070 1084.400 ;
        RECT 1702.090 1084.120 1702.370 1084.400 ;
        RECT 1711.750 1084.120 1712.030 1084.400 ;
        RECT 1798.690 1084.120 1798.970 1084.400 ;
        RECT 1801.910 1084.120 1802.190 1084.400 ;
        RECT 1895.290 1084.120 1895.570 1084.400 ;
        RECT 1355.710 1082.760 1355.990 1083.040 ;
        RECT 2052.610 1085.480 2052.890 1085.760 ;
        RECT 2028.230 1084.120 2028.510 1084.400 ;
        RECT 1932.090 1083.440 1932.370 1083.720 ;
        RECT 2124.830 1084.800 2125.110 1085.080 ;
        RECT 2090.330 1084.120 2090.610 1084.400 ;
        RECT 2052.610 1083.440 2052.890 1083.720 ;
        RECT 1895.290 1082.080 1895.570 1082.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1084.340 2924.800 1085.540 ;
=======
        RECT 1246.665 2498.140 1246.995 2498.145 ;
        RECT 1246.665 2498.130 1247.250 2498.140 ;
        RECT 1246.665 2497.830 1247.450 2498.130 ;
        RECT 1246.665 2497.820 1247.250 2497.830 ;
        RECT 1246.665 2497.815 1246.995 2497.820 ;
        RECT 1579.245 1086.450 1579.575 1086.465 ;
        RECT 1532.110 1086.150 1579.575 1086.450 ;
        RECT 1331.510 1085.090 1331.890 1085.100 ;
        RECT 1355.685 1085.090 1356.015 1085.105 ;
        RECT 1272.670 1084.790 1314.370 1085.090 ;
        RECT 1246.870 1084.410 1247.250 1084.420 ;
        RECT 1272.670 1084.410 1272.970 1084.790 ;
        RECT 1246.870 1084.110 1272.970 1084.410 ;
        RECT 1246.870 1084.100 1247.250 1084.110 ;
        RECT 1314.070 1083.730 1314.370 1084.790 ;
        RECT 1331.510 1084.790 1356.015 1085.090 ;
        RECT 1331.510 1084.780 1331.890 1084.790 ;
        RECT 1355.685 1084.775 1356.015 1084.790 ;
        RECT 1483.105 1085.090 1483.435 1085.105 ;
        RECT 1532.110 1085.090 1532.410 1086.150 ;
        RECT 1579.245 1086.135 1579.575 1086.150 ;
        RECT 1980.110 1086.450 1980.490 1086.460 ;
        RECT 2028.205 1086.450 2028.535 1086.465 ;
        RECT 1980.110 1086.150 2028.535 1086.450 ;
        RECT 1980.110 1086.140 1980.490 1086.150 ;
        RECT 2028.205 1086.135 2028.535 1086.150 ;
        RECT 2052.585 1085.770 2052.915 1085.785 ;
        RECT 2028.910 1085.470 2052.915 1085.770 ;
        RECT 1483.105 1084.790 1532.410 1085.090 ;
        RECT 1946.325 1085.090 1946.655 1085.105 ;
        RECT 1980.110 1085.090 1980.490 1085.100 ;
        RECT 1946.325 1084.790 1980.490 1085.090 ;
        RECT 1483.105 1084.775 1483.435 1084.790 ;
        RECT 1946.325 1084.775 1946.655 1084.790 ;
        RECT 1980.110 1084.780 1980.490 1084.790 ;
        RECT 1483.105 1084.410 1483.435 1084.425 ;
        RECT 1435.510 1084.110 1483.435 1084.410 ;
        RECT 1331.510 1083.730 1331.890 1083.740 ;
        RECT 1435.510 1083.730 1435.810 1084.110 ;
        RECT 1483.105 1084.095 1483.435 1084.110 ;
        RECT 1579.245 1084.410 1579.575 1084.425 ;
        RECT 1606.385 1084.410 1606.715 1084.425 ;
        RECT 1579.245 1084.110 1606.715 1084.410 ;
        RECT 1579.245 1084.095 1579.575 1084.110 ;
        RECT 1606.385 1084.095 1606.715 1084.110 ;
        RECT 1607.765 1084.410 1608.095 1084.425 ;
        RECT 1702.065 1084.410 1702.395 1084.425 ;
        RECT 1607.765 1084.110 1641.890 1084.410 ;
        RECT 1607.765 1084.095 1608.095 1084.110 ;
        RECT 1314.070 1083.430 1331.890 1083.730 ;
        RECT 1331.510 1083.420 1331.890 1083.430 ;
        RECT 1399.630 1083.430 1400.850 1083.730 ;
        RECT 1355.685 1083.050 1356.015 1083.065 ;
        RECT 1399.630 1083.050 1399.930 1083.430 ;
        RECT 1355.685 1082.750 1399.930 1083.050 ;
        RECT 1400.550 1083.050 1400.850 1083.430 ;
        RECT 1415.270 1083.430 1435.810 1083.730 ;
        RECT 1641.590 1083.730 1641.890 1084.110 ;
        RECT 1656.310 1084.110 1702.395 1084.410 ;
        RECT 1656.310 1083.730 1656.610 1084.110 ;
        RECT 1702.065 1084.095 1702.395 1084.110 ;
        RECT 1711.725 1084.410 1712.055 1084.425 ;
        RECT 1798.665 1084.410 1798.995 1084.425 ;
        RECT 1711.725 1084.110 1738.490 1084.410 ;
        RECT 1711.725 1084.095 1712.055 1084.110 ;
        RECT 1641.590 1083.430 1656.610 1083.730 ;
        RECT 1738.190 1083.730 1738.490 1084.110 ;
        RECT 1752.910 1084.110 1798.995 1084.410 ;
        RECT 1752.910 1083.730 1753.210 1084.110 ;
        RECT 1798.665 1084.095 1798.995 1084.110 ;
        RECT 1801.885 1084.410 1802.215 1084.425 ;
        RECT 1895.265 1084.410 1895.595 1084.425 ;
        RECT 1801.885 1084.110 1835.090 1084.410 ;
        RECT 1801.885 1084.095 1802.215 1084.110 ;
        RECT 1738.190 1083.430 1753.210 1083.730 ;
        RECT 1834.790 1083.730 1835.090 1084.110 ;
        RECT 1849.510 1084.110 1895.595 1084.410 ;
        RECT 1849.510 1083.730 1849.810 1084.110 ;
        RECT 1895.265 1084.095 1895.595 1084.110 ;
        RECT 2028.205 1084.410 2028.535 1084.425 ;
        RECT 2028.910 1084.410 2029.210 1085.470 ;
        RECT 2052.585 1085.455 2052.915 1085.470 ;
        RECT 2124.805 1085.090 2125.135 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2124.805 1084.790 2159.850 1085.090 ;
        RECT 2124.805 1084.775 2125.135 1084.790 ;
        RECT 2090.305 1084.410 2090.635 1084.425 ;
        RECT 2028.205 1084.110 2029.210 1084.410 ;
        RECT 2076.750 1084.110 2090.635 1084.410 ;
        RECT 2159.550 1084.410 2159.850 1084.790 ;
        RECT 2208.310 1084.790 2256.450 1085.090 ;
        RECT 2159.550 1084.110 2207.690 1084.410 ;
        RECT 2028.205 1084.095 2028.535 1084.110 ;
        RECT 1932.065 1083.730 1932.395 1083.745 ;
        RECT 1834.790 1083.430 1849.810 1083.730 ;
        RECT 1931.390 1083.430 1932.395 1083.730 ;
        RECT 1415.270 1083.050 1415.570 1083.430 ;
        RECT 1400.550 1082.750 1415.570 1083.050 ;
        RECT 1355.685 1082.735 1356.015 1082.750 ;
        RECT 1895.265 1082.370 1895.595 1082.385 ;
        RECT 1931.390 1082.370 1931.690 1083.430 ;
        RECT 1932.065 1083.415 1932.395 1083.430 ;
        RECT 2052.585 1083.730 2052.915 1083.745 ;
        RECT 2076.750 1083.730 2077.050 1084.110 ;
        RECT 2090.305 1084.095 2090.635 1084.110 ;
        RECT 2052.585 1083.430 2077.050 1083.730 ;
        RECT 2207.390 1083.730 2207.690 1084.110 ;
        RECT 2208.310 1083.730 2208.610 1084.790 ;
        RECT 2256.150 1084.410 2256.450 1084.790 ;
        RECT 2304.910 1084.790 2353.050 1085.090 ;
        RECT 2256.150 1084.110 2304.290 1084.410 ;
        RECT 2207.390 1083.430 2208.610 1083.730 ;
        RECT 2303.990 1083.730 2304.290 1084.110 ;
        RECT 2304.910 1083.730 2305.210 1084.790 ;
        RECT 2352.750 1084.410 2353.050 1084.790 ;
        RECT 2401.510 1084.790 2449.650 1085.090 ;
        RECT 2352.750 1084.110 2400.890 1084.410 ;
        RECT 2303.990 1083.430 2305.210 1083.730 ;
        RECT 2400.590 1083.730 2400.890 1084.110 ;
        RECT 2401.510 1083.730 2401.810 1084.790 ;
        RECT 2449.350 1084.410 2449.650 1084.790 ;
        RECT 2498.110 1084.790 2546.250 1085.090 ;
        RECT 2449.350 1084.110 2497.490 1084.410 ;
        RECT 2400.590 1083.430 2401.810 1083.730 ;
        RECT 2497.190 1083.730 2497.490 1084.110 ;
        RECT 2498.110 1083.730 2498.410 1084.790 ;
        RECT 2545.950 1084.410 2546.250 1084.790 ;
        RECT 2594.710 1084.790 2642.850 1085.090 ;
        RECT 2545.950 1084.110 2594.090 1084.410 ;
        RECT 2497.190 1083.430 2498.410 1083.730 ;
        RECT 2593.790 1083.730 2594.090 1084.110 ;
        RECT 2594.710 1083.730 2595.010 1084.790 ;
        RECT 2642.550 1084.410 2642.850 1084.790 ;
        RECT 2691.310 1084.790 2739.450 1085.090 ;
        RECT 2642.550 1084.110 2690.690 1084.410 ;
        RECT 2593.790 1083.430 2595.010 1083.730 ;
        RECT 2690.390 1083.730 2690.690 1084.110 ;
        RECT 2691.310 1083.730 2691.610 1084.790 ;
        RECT 2739.150 1084.410 2739.450 1084.790 ;
        RECT 2787.910 1084.790 2836.050 1085.090 ;
        RECT 2739.150 1084.110 2787.290 1084.410 ;
        RECT 2690.390 1083.430 2691.610 1083.730 ;
        RECT 2786.990 1083.730 2787.290 1084.110 ;
        RECT 2787.910 1083.730 2788.210 1084.790 ;
        RECT 2835.750 1084.410 2836.050 1084.790 ;
        RECT 2916.710 1084.790 2924.800 1085.090 ;
        RECT 2916.710 1084.410 2917.010 1084.790 ;
        RECT 2835.750 1084.110 2883.890 1084.410 ;
        RECT 2786.990 1083.430 2788.210 1083.730 ;
        RECT 2883.590 1083.730 2883.890 1084.110 ;
        RECT 2884.510 1084.110 2917.010 1084.410 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
        RECT 2884.510 1083.730 2884.810 1084.110 ;
        RECT 2883.590 1083.430 2884.810 1083.730 ;
        RECT 2052.585 1083.415 2052.915 1083.430 ;
        RECT 1895.265 1082.070 1931.690 1082.370 ;
        RECT 1895.265 1082.055 1895.595 1082.070 ;
      LAYER via3 ;
        RECT 1246.900 2497.820 1247.220 2498.140 ;
        RECT 1246.900 1084.100 1247.220 1084.420 ;
        RECT 1331.540 1084.780 1331.860 1085.100 ;
        RECT 1980.140 1086.140 1980.460 1086.460 ;
        RECT 1980.140 1084.780 1980.460 1085.100 ;
        RECT 1331.540 1083.420 1331.860 1083.740 ;
      LAYER met4 ;
        RECT 1246.895 2497.815 1247.225 2498.145 ;
        RECT 1246.910 1084.425 1247.210 2497.815 ;
        RECT 1980.135 1086.135 1980.465 1086.465 ;
        RECT 1980.150 1085.105 1980.450 1086.135 ;
        RECT 1331.535 1084.775 1331.865 1085.105 ;
        RECT 1980.135 1084.775 1980.465 1085.105 ;
        RECT 1246.895 1084.095 1247.225 1084.425 ;
        RECT 1331.550 1083.745 1331.850 1084.775 ;
        RECT 1331.535 1083.415 1331.865 1083.745 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2090.310 1319.100 2090.630 1319.160 ;
        RECT 2124.810 1319.100 2125.130 1319.160 ;
        RECT 2090.310 1318.960 2125.130 1319.100 ;
        RECT 2090.310 1318.900 2090.630 1318.960 ;
        RECT 2124.810 1318.900 2125.130 1318.960 ;
        RECT 1606.390 1318.760 1606.710 1318.820 ;
        RECT 1607.770 1318.760 1608.090 1318.820 ;
        RECT 1606.390 1318.620 1608.090 1318.760 ;
        RECT 1606.390 1318.560 1606.710 1318.620 ;
        RECT 1607.770 1318.560 1608.090 1318.620 ;
        RECT 1702.070 1318.760 1702.390 1318.820 ;
        RECT 1711.730 1318.760 1712.050 1318.820 ;
        RECT 1702.070 1318.620 1712.050 1318.760 ;
        RECT 1702.070 1318.560 1702.390 1318.620 ;
        RECT 1711.730 1318.560 1712.050 1318.620 ;
        RECT 1798.670 1318.760 1798.990 1318.820 ;
        RECT 1801.890 1318.760 1802.210 1318.820 ;
        RECT 1798.670 1318.620 1802.210 1318.760 ;
        RECT 1798.670 1318.560 1798.990 1318.620 ;
        RECT 1801.890 1318.560 1802.210 1318.620 ;
        RECT 1932.070 1318.420 1932.390 1318.480 ;
        RECT 1946.330 1318.420 1946.650 1318.480 ;
        RECT 1932.070 1318.280 1946.650 1318.420 ;
        RECT 1932.070 1318.220 1932.390 1318.280 ;
        RECT 1946.330 1318.220 1946.650 1318.280 ;
      LAYER via ;
        RECT 2090.340 1318.900 2090.600 1319.160 ;
        RECT 2124.840 1318.900 2125.100 1319.160 ;
        RECT 1606.420 1318.560 1606.680 1318.820 ;
        RECT 1607.800 1318.560 1608.060 1318.820 ;
        RECT 1702.100 1318.560 1702.360 1318.820 ;
        RECT 1711.760 1318.560 1712.020 1318.820 ;
        RECT 1798.700 1318.560 1798.960 1318.820 ;
        RECT 1801.920 1318.560 1802.180 1318.820 ;
        RECT 1932.100 1318.220 1932.360 1318.480 ;
        RECT 1946.360 1318.220 1946.620 1318.480 ;
      LAYER met2 ;
        RECT 1265.550 2498.050 1265.830 2500.000 ;
        RECT 1267.390 2498.050 1267.670 2498.165 ;
        RECT 1265.550 2497.910 1267.670 2498.050 ;
        RECT 1265.550 2496.000 1265.830 2497.910 ;
        RECT 1267.390 2497.795 1267.670 2497.910 ;
        RECT 2028.230 1320.715 2028.510 1321.085 ;
        RECT 1448.630 1319.355 1448.910 1319.725 ;
        RECT 1946.350 1319.355 1946.630 1319.725 ;
        RECT 1448.700 1319.045 1448.840 1319.355 ;
        RECT 1448.630 1318.675 1448.910 1319.045 ;
        RECT 1606.410 1318.675 1606.690 1319.045 ;
        RECT 1607.790 1318.675 1608.070 1319.045 ;
        RECT 1702.090 1318.675 1702.370 1319.045 ;
        RECT 1711.750 1318.675 1712.030 1319.045 ;
        RECT 1798.690 1318.675 1798.970 1319.045 ;
        RECT 1801.910 1318.675 1802.190 1319.045 ;
        RECT 1895.290 1318.675 1895.570 1319.045 ;
        RECT 1606.420 1318.530 1606.680 1318.675 ;
        RECT 1607.800 1318.530 1608.060 1318.675 ;
        RECT 1702.100 1318.530 1702.360 1318.675 ;
        RECT 1711.760 1318.530 1712.020 1318.675 ;
        RECT 1798.700 1318.530 1798.960 1318.675 ;
        RECT 1801.920 1318.530 1802.180 1318.675 ;
        RECT 1895.360 1317.005 1895.500 1318.675 ;
        RECT 1946.420 1318.510 1946.560 1319.355 ;
        RECT 2028.300 1319.045 2028.440 1320.715 ;
        RECT 2052.610 1320.035 2052.890 1320.405 ;
        RECT 2028.230 1318.675 2028.510 1319.045 ;
        RECT 1932.100 1318.365 1932.360 1318.510 ;
        RECT 1932.090 1317.995 1932.370 1318.365 ;
        RECT 1946.360 1318.190 1946.620 1318.510 ;
        RECT 2052.680 1318.365 2052.820 1320.035 ;
        RECT 2124.830 1319.355 2125.110 1319.725 ;
        RECT 2124.900 1319.190 2125.040 1319.355 ;
        RECT 2090.340 1319.045 2090.600 1319.190 ;
        RECT 2090.330 1318.675 2090.610 1319.045 ;
        RECT 2124.840 1318.870 2125.100 1319.190 ;
        RECT 2052.610 1317.995 2052.890 1318.365 ;
        RECT 1895.290 1316.635 1895.570 1317.005 ;
      LAYER via2 ;
        RECT 1267.390 2497.840 1267.670 2498.120 ;
        RECT 2028.230 1320.760 2028.510 1321.040 ;
        RECT 1448.630 1319.400 1448.910 1319.680 ;
        RECT 1946.350 1319.400 1946.630 1319.680 ;
        RECT 1448.630 1318.720 1448.910 1319.000 ;
        RECT 1606.410 1318.720 1606.690 1319.000 ;
        RECT 1607.790 1318.720 1608.070 1319.000 ;
        RECT 1702.090 1318.720 1702.370 1319.000 ;
        RECT 1711.750 1318.720 1712.030 1319.000 ;
        RECT 1798.690 1318.720 1798.970 1319.000 ;
        RECT 1801.910 1318.720 1802.190 1319.000 ;
        RECT 1895.290 1318.720 1895.570 1319.000 ;
        RECT 2052.610 1320.080 2052.890 1320.360 ;
        RECT 2028.230 1318.720 2028.510 1319.000 ;
        RECT 1932.090 1318.040 1932.370 1318.320 ;
        RECT 2124.830 1319.400 2125.110 1319.680 ;
        RECT 2090.330 1318.720 2090.610 1319.000 ;
        RECT 2052.610 1318.040 2052.890 1318.320 ;
        RECT 1895.290 1316.680 1895.570 1316.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1318.940 2924.800 1320.140 ;
=======
        RECT 1267.365 2498.130 1267.695 2498.145 ;
        RECT 1268.950 2498.130 1269.330 2498.140 ;
        RECT 1267.365 2497.830 1269.330 2498.130 ;
        RECT 1267.365 2497.815 1267.695 2497.830 ;
        RECT 1268.950 2497.820 1269.330 2497.830 ;
        RECT 1980.110 1321.050 1980.490 1321.060 ;
        RECT 2028.205 1321.050 2028.535 1321.065 ;
        RECT 1980.110 1320.750 2028.535 1321.050 ;
        RECT 1980.110 1320.740 1980.490 1320.750 ;
        RECT 2028.205 1320.735 2028.535 1320.750 ;
        RECT 1268.950 1320.370 1269.330 1320.380 ;
        RECT 2052.585 1320.370 2052.915 1320.385 ;
        RECT 1268.950 1320.070 1365.890 1320.370 ;
        RECT 1268.950 1320.060 1269.330 1320.070 ;
        RECT 1365.590 1319.010 1365.890 1320.070 ;
        RECT 2028.910 1320.070 2052.915 1320.370 ;
        RECT 1448.605 1319.690 1448.935 1319.705 ;
        RECT 1946.325 1319.690 1946.655 1319.705 ;
        RECT 1980.110 1319.690 1980.490 1319.700 ;
        RECT 1448.605 1319.390 1511.250 1319.690 ;
        RECT 1448.605 1319.375 1448.935 1319.390 ;
        RECT 1448.605 1319.010 1448.935 1319.025 ;
        RECT 1365.590 1318.710 1448.935 1319.010 ;
        RECT 1448.605 1318.695 1448.935 1318.710 ;
        RECT 1510.950 1318.330 1511.250 1319.390 ;
        RECT 1946.325 1319.390 1980.490 1319.690 ;
        RECT 1946.325 1319.375 1946.655 1319.390 ;
        RECT 1980.110 1319.380 1980.490 1319.390 ;
        RECT 1606.385 1319.010 1606.715 1319.025 ;
        RECT 1559.710 1318.710 1606.715 1319.010 ;
        RECT 1559.710 1318.330 1560.010 1318.710 ;
        RECT 1606.385 1318.695 1606.715 1318.710 ;
        RECT 1607.765 1319.010 1608.095 1319.025 ;
        RECT 1702.065 1319.010 1702.395 1319.025 ;
        RECT 1607.765 1318.710 1641.890 1319.010 ;
        RECT 1607.765 1318.695 1608.095 1318.710 ;
        RECT 1510.950 1318.030 1560.010 1318.330 ;
        RECT 1641.590 1318.330 1641.890 1318.710 ;
        RECT 1656.310 1318.710 1702.395 1319.010 ;
        RECT 1656.310 1318.330 1656.610 1318.710 ;
        RECT 1702.065 1318.695 1702.395 1318.710 ;
        RECT 1711.725 1319.010 1712.055 1319.025 ;
        RECT 1798.665 1319.010 1798.995 1319.025 ;
        RECT 1711.725 1318.710 1738.490 1319.010 ;
        RECT 1711.725 1318.695 1712.055 1318.710 ;
        RECT 1641.590 1318.030 1656.610 1318.330 ;
        RECT 1738.190 1318.330 1738.490 1318.710 ;
        RECT 1752.910 1318.710 1798.995 1319.010 ;
        RECT 1752.910 1318.330 1753.210 1318.710 ;
        RECT 1798.665 1318.695 1798.995 1318.710 ;
        RECT 1801.885 1319.010 1802.215 1319.025 ;
        RECT 1895.265 1319.010 1895.595 1319.025 ;
        RECT 1801.885 1318.710 1835.090 1319.010 ;
        RECT 1801.885 1318.695 1802.215 1318.710 ;
        RECT 1738.190 1318.030 1753.210 1318.330 ;
        RECT 1834.790 1318.330 1835.090 1318.710 ;
        RECT 1849.510 1318.710 1895.595 1319.010 ;
        RECT 1849.510 1318.330 1849.810 1318.710 ;
        RECT 1895.265 1318.695 1895.595 1318.710 ;
        RECT 2028.205 1319.010 2028.535 1319.025 ;
        RECT 2028.910 1319.010 2029.210 1320.070 ;
        RECT 2052.585 1320.055 2052.915 1320.070 ;
        RECT 2124.805 1319.690 2125.135 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2124.805 1319.390 2159.850 1319.690 ;
        RECT 2124.805 1319.375 2125.135 1319.390 ;
        RECT 2090.305 1319.010 2090.635 1319.025 ;
        RECT 2028.205 1318.710 2029.210 1319.010 ;
        RECT 2076.750 1318.710 2090.635 1319.010 ;
        RECT 2159.550 1319.010 2159.850 1319.390 ;
        RECT 2208.310 1319.390 2256.450 1319.690 ;
        RECT 2159.550 1318.710 2207.690 1319.010 ;
        RECT 2028.205 1318.695 2028.535 1318.710 ;
        RECT 1932.065 1318.330 1932.395 1318.345 ;
        RECT 1834.790 1318.030 1849.810 1318.330 ;
        RECT 1931.390 1318.030 1932.395 1318.330 ;
        RECT 1895.265 1316.970 1895.595 1316.985 ;
        RECT 1931.390 1316.970 1931.690 1318.030 ;
        RECT 1932.065 1318.015 1932.395 1318.030 ;
        RECT 2052.585 1318.330 2052.915 1318.345 ;
        RECT 2076.750 1318.330 2077.050 1318.710 ;
        RECT 2090.305 1318.695 2090.635 1318.710 ;
        RECT 2052.585 1318.030 2077.050 1318.330 ;
        RECT 2207.390 1318.330 2207.690 1318.710 ;
        RECT 2208.310 1318.330 2208.610 1319.390 ;
        RECT 2256.150 1319.010 2256.450 1319.390 ;
        RECT 2304.910 1319.390 2353.050 1319.690 ;
        RECT 2256.150 1318.710 2304.290 1319.010 ;
        RECT 2207.390 1318.030 2208.610 1318.330 ;
        RECT 2303.990 1318.330 2304.290 1318.710 ;
        RECT 2304.910 1318.330 2305.210 1319.390 ;
        RECT 2352.750 1319.010 2353.050 1319.390 ;
        RECT 2401.510 1319.390 2449.650 1319.690 ;
        RECT 2352.750 1318.710 2400.890 1319.010 ;
        RECT 2303.990 1318.030 2305.210 1318.330 ;
        RECT 2400.590 1318.330 2400.890 1318.710 ;
        RECT 2401.510 1318.330 2401.810 1319.390 ;
        RECT 2449.350 1319.010 2449.650 1319.390 ;
        RECT 2498.110 1319.390 2546.250 1319.690 ;
        RECT 2449.350 1318.710 2497.490 1319.010 ;
        RECT 2400.590 1318.030 2401.810 1318.330 ;
        RECT 2497.190 1318.330 2497.490 1318.710 ;
        RECT 2498.110 1318.330 2498.410 1319.390 ;
        RECT 2545.950 1319.010 2546.250 1319.390 ;
        RECT 2594.710 1319.390 2642.850 1319.690 ;
        RECT 2545.950 1318.710 2594.090 1319.010 ;
        RECT 2497.190 1318.030 2498.410 1318.330 ;
        RECT 2593.790 1318.330 2594.090 1318.710 ;
        RECT 2594.710 1318.330 2595.010 1319.390 ;
        RECT 2642.550 1319.010 2642.850 1319.390 ;
        RECT 2691.310 1319.390 2739.450 1319.690 ;
        RECT 2642.550 1318.710 2690.690 1319.010 ;
        RECT 2593.790 1318.030 2595.010 1318.330 ;
        RECT 2690.390 1318.330 2690.690 1318.710 ;
        RECT 2691.310 1318.330 2691.610 1319.390 ;
        RECT 2739.150 1319.010 2739.450 1319.390 ;
        RECT 2787.910 1319.390 2836.050 1319.690 ;
        RECT 2739.150 1318.710 2787.290 1319.010 ;
        RECT 2690.390 1318.030 2691.610 1318.330 ;
        RECT 2786.990 1318.330 2787.290 1318.710 ;
        RECT 2787.910 1318.330 2788.210 1319.390 ;
        RECT 2835.750 1319.010 2836.050 1319.390 ;
        RECT 2916.710 1319.390 2924.800 1319.690 ;
        RECT 2916.710 1319.010 2917.010 1319.390 ;
        RECT 2835.750 1318.710 2883.890 1319.010 ;
        RECT 2786.990 1318.030 2788.210 1318.330 ;
        RECT 2883.590 1318.330 2883.890 1318.710 ;
        RECT 2884.510 1318.710 2917.010 1319.010 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT 2884.510 1318.330 2884.810 1318.710 ;
        RECT 2883.590 1318.030 2884.810 1318.330 ;
        RECT 2052.585 1318.015 2052.915 1318.030 ;
        RECT 1895.265 1316.670 1931.690 1316.970 ;
        RECT 1895.265 1316.655 1895.595 1316.670 ;
      LAYER via3 ;
        RECT 1268.980 2497.820 1269.300 2498.140 ;
        RECT 1980.140 1320.740 1980.460 1321.060 ;
        RECT 1268.980 1320.060 1269.300 1320.380 ;
        RECT 1980.140 1319.380 1980.460 1319.700 ;
      LAYER met4 ;
        RECT 1268.975 2497.815 1269.305 2498.145 ;
        RECT 1268.990 1320.385 1269.290 2497.815 ;
        RECT 1980.135 1320.735 1980.465 1321.065 ;
        RECT 1268.975 1320.055 1269.305 1320.385 ;
        RECT 1980.150 1319.705 1980.450 1320.735 ;
        RECT 1980.135 1319.375 1980.465 1319.705 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1285.310 2513.860 1285.630 2513.920 ;
        RECT 2639.090 2513.860 2639.410 2513.920 ;
        RECT 1285.310 2513.720 2639.410 2513.860 ;
        RECT 1285.310 2513.660 1285.630 2513.720 ;
        RECT 2639.090 2513.660 2639.410 2513.720 ;
        RECT 2639.090 1559.140 2639.410 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2639.090 1559.000 2901.150 1559.140 ;
        RECT 2639.090 1558.940 2639.410 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 1285.340 2513.660 1285.600 2513.920 ;
        RECT 2639.120 2513.660 2639.380 2513.920 ;
        RECT 2639.120 1558.940 2639.380 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 1285.340 2513.630 1285.600 2513.950 ;
        RECT 2639.120 2513.630 2639.380 2513.950 ;
        RECT 1285.400 2500.000 1285.540 2513.630 ;
        RECT 1285.330 2496.000 1285.610 2500.000 ;
        RECT 2639.180 1559.230 2639.320 2513.630 ;
        RECT 2639.120 1558.910 2639.380 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1553.540 2924.800 1554.740 ;
=======
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1926.165 2513.365 1926.335 2514.555 ;
      LAYER mcon ;
        RECT 1926.165 2514.385 1926.335 2514.555 ;
      LAYER met1 ;
        RECT 1305.090 2514.540 1305.410 2514.600 ;
        RECT 1926.105 2514.540 1926.395 2514.585 ;
        RECT 1305.090 2514.400 1926.395 2514.540 ;
        RECT 1305.090 2514.340 1305.410 2514.400 ;
        RECT 1926.105 2514.355 1926.395 2514.400 ;
        RECT 1926.105 2513.520 1926.395 2513.565 ;
        RECT 1949.090 2513.520 1949.410 2513.580 ;
        RECT 1926.105 2513.380 1949.410 2513.520 ;
        RECT 1926.105 2513.335 1926.395 2513.380 ;
        RECT 1949.090 2513.320 1949.410 2513.380 ;
        RECT 1949.090 1793.740 1949.410 1793.800 ;
        RECT 2900.830 1793.740 2901.150 1793.800 ;
        RECT 1949.090 1793.600 2901.150 1793.740 ;
        RECT 1949.090 1793.540 1949.410 1793.600 ;
        RECT 2900.830 1793.540 2901.150 1793.600 ;
      LAYER via ;
        RECT 1305.120 2514.340 1305.380 2514.600 ;
        RECT 1949.120 2513.320 1949.380 2513.580 ;
        RECT 1949.120 1793.540 1949.380 1793.800 ;
        RECT 2900.860 1793.540 2901.120 1793.800 ;
      LAYER met2 ;
        RECT 1305.120 2514.310 1305.380 2514.630 ;
        RECT 1305.180 2500.000 1305.320 2514.310 ;
        RECT 1949.120 2513.290 1949.380 2513.610 ;
        RECT 1305.110 2496.000 1305.390 2500.000 ;
        RECT 1949.180 1793.830 1949.320 2513.290 ;
        RECT 1949.120 1793.510 1949.380 1793.830 ;
        RECT 2900.860 1793.510 2901.120 1793.830 ;
        RECT 2900.920 1789.605 2901.060 1793.510 ;
        RECT 2900.850 1789.235 2901.130 1789.605 ;
      LAYER via2 ;
        RECT 2900.850 1789.280 2901.130 1789.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1788.820 2924.800 1790.020 ;
=======
        RECT 2900.825 1789.570 2901.155 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.825 1789.270 2924.800 1789.570 ;
        RECT 2900.825 1789.255 2901.155 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1950.470 2516.580 1950.790 2516.640 ;
        RECT 1932.620 2516.440 1950.790 2516.580 ;
        RECT 1324.870 2516.240 1325.190 2516.300 ;
        RECT 1932.620 2516.240 1932.760 2516.440 ;
        RECT 1950.470 2516.380 1950.790 2516.440 ;
        RECT 1324.870 2516.100 1932.760 2516.240 ;
        RECT 1324.870 2516.040 1325.190 2516.100 ;
        RECT 1950.470 2028.340 1950.790 2028.400 ;
        RECT 2900.830 2028.340 2901.150 2028.400 ;
        RECT 1950.470 2028.200 2901.150 2028.340 ;
        RECT 1950.470 2028.140 1950.790 2028.200 ;
        RECT 2900.830 2028.140 2901.150 2028.200 ;
      LAYER via ;
        RECT 1324.900 2516.040 1325.160 2516.300 ;
        RECT 1950.500 2516.380 1950.760 2516.640 ;
        RECT 1950.500 2028.140 1950.760 2028.400 ;
        RECT 2900.860 2028.140 2901.120 2028.400 ;
      LAYER met2 ;
        RECT 1950.500 2516.350 1950.760 2516.670 ;
        RECT 1324.900 2516.010 1325.160 2516.330 ;
        RECT 1324.960 2500.000 1325.100 2516.010 ;
        RECT 1324.890 2496.000 1325.170 2500.000 ;
        RECT 1950.560 2028.430 1950.700 2516.350 ;
        RECT 1950.500 2028.110 1950.760 2028.430 ;
        RECT 2900.860 2028.110 2901.120 2028.430 ;
        RECT 2900.920 2024.205 2901.060 2028.110 ;
        RECT 2900.850 2023.835 2901.130 2024.205 ;
      LAYER via2 ;
        RECT 2900.850 2023.880 2901.130 2024.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2023.420 2924.800 2024.620 ;
=======
        RECT 2900.825 2024.170 2901.155 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.825 2023.870 2924.800 2024.170 ;
        RECT 2900.825 2023.855 2901.155 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1931.685 2517.105 1931.855 2518.295 ;
      LAYER mcon ;
        RECT 1931.685 2518.125 1931.855 2518.295 ;
      LAYER met1 ;
        RECT 1931.625 2518.280 1931.915 2518.325 ;
        RECT 1952.310 2518.280 1952.630 2518.340 ;
        RECT 1931.625 2518.140 1952.630 2518.280 ;
        RECT 1931.625 2518.095 1931.915 2518.140 ;
        RECT 1952.310 2518.080 1952.630 2518.140 ;
        RECT 1344.650 2517.260 1344.970 2517.320 ;
        RECT 1931.625 2517.260 1931.915 2517.305 ;
        RECT 1344.650 2517.120 1931.915 2517.260 ;
        RECT 1344.650 2517.060 1344.970 2517.120 ;
        RECT 1931.625 2517.075 1931.915 2517.120 ;
        RECT 1952.310 2262.940 1952.630 2263.000 ;
        RECT 2900.830 2262.940 2901.150 2263.000 ;
        RECT 1952.310 2262.800 2901.150 2262.940 ;
        RECT 1952.310 2262.740 1952.630 2262.800 ;
        RECT 2900.830 2262.740 2901.150 2262.800 ;
      LAYER via ;
        RECT 1952.340 2518.080 1952.600 2518.340 ;
        RECT 1344.680 2517.060 1344.940 2517.320 ;
        RECT 1952.340 2262.740 1952.600 2263.000 ;
        RECT 2900.860 2262.740 2901.120 2263.000 ;
      LAYER met2 ;
        RECT 1952.340 2518.050 1952.600 2518.370 ;
        RECT 1344.680 2517.030 1344.940 2517.350 ;
        RECT 1344.740 2500.000 1344.880 2517.030 ;
        RECT 1344.670 2496.000 1344.950 2500.000 ;
        RECT 1952.400 2263.030 1952.540 2518.050 ;
        RECT 1952.340 2262.710 1952.600 2263.030 ;
        RECT 2900.860 2262.710 2901.120 2263.030 ;
        RECT 2900.920 2258.805 2901.060 2262.710 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2258.020 2924.800 2259.220 ;
=======
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 0.300 ;
=======
      LAYER met1 ;
        RECT 634.410 54.300 634.730 54.360 ;
        RECT 1319.350 54.300 1319.670 54.360 ;
        RECT 634.410 54.160 1319.670 54.300 ;
        RECT 634.410 54.100 634.730 54.160 ;
        RECT 1319.350 54.100 1319.670 54.160 ;
      LAYER via ;
        RECT 634.440 54.100 634.700 54.360 ;
        RECT 1319.380 54.100 1319.640 54.360 ;
      LAYER met2 ;
        RECT 1320.750 1700.410 1321.030 1704.000 ;
        RECT 1319.440 1700.270 1321.030 1700.410 ;
        RECT 1319.440 54.390 1319.580 1700.270 ;
        RECT 1320.750 1700.000 1321.030 1700.270 ;
        RECT 634.440 54.070 634.700 54.390 ;
        RECT 1319.380 54.070 1319.640 54.390 ;
        RECT 634.500 17.410 634.640 54.070 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1802.350 1683.920 1802.670 1683.980 ;
        RECT 1806.950 1683.920 1807.270 1683.980 ;
        RECT 1802.350 1683.780 1807.270 1683.920 ;
        RECT 1802.350 1683.720 1802.670 1683.780 ;
        RECT 1806.950 1683.720 1807.270 1683.780 ;
        RECT 1806.950 44.780 1807.270 44.840 ;
        RECT 2417.370 44.780 2417.690 44.840 ;
        RECT 1806.950 44.640 2417.690 44.780 ;
        RECT 1806.950 44.580 1807.270 44.640 ;
        RECT 2417.370 44.580 2417.690 44.640 ;
      LAYER via ;
        RECT 1802.380 1683.720 1802.640 1683.980 ;
        RECT 1806.980 1683.720 1807.240 1683.980 ;
        RECT 1806.980 44.580 1807.240 44.840 ;
        RECT 2417.400 44.580 2417.660 44.840 ;
      LAYER met2 ;
        RECT 1802.370 1700.000 1802.650 1704.000 ;
        RECT 1802.440 1684.010 1802.580 1700.000 ;
        RECT 1802.380 1683.690 1802.640 1684.010 ;
        RECT 1806.980 1683.690 1807.240 1684.010 ;
        RECT 1807.040 44.870 1807.180 1683.690 ;
        RECT 1806.980 44.550 1807.240 44.870 ;
        RECT 2417.400 44.550 2417.660 44.870 ;
        RECT 2417.460 2.400 2417.600 44.550 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2434.730 -4.800 2435.290 0.300 ;
=======
        RECT 1807.430 1700.410 1807.710 1704.000 ;
        RECT 1806.580 1700.270 1807.710 1700.410 ;
        RECT 1806.580 48.125 1806.720 1700.270 ;
        RECT 1807.430 1700.000 1807.710 1700.270 ;
        RECT 1806.510 47.755 1806.790 48.125 ;
        RECT 2434.870 47.755 2435.150 48.125 ;
        RECT 2434.940 2.400 2435.080 47.755 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
      LAYER via2 ;
        RECT 1806.510 47.800 1806.790 48.080 ;
        RECT 2434.870 47.800 2435.150 48.080 ;
      LAYER met3 ;
        RECT 1806.485 48.090 1806.815 48.105 ;
        RECT 2434.845 48.090 2435.175 48.105 ;
        RECT 1806.485 47.790 2435.175 48.090 ;
        RECT 1806.485 47.775 1806.815 47.790 ;
        RECT 2434.845 47.775 2435.175 47.790 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2452.670 -4.800 2453.230 0.300 ;
=======
        RECT 1812.030 1700.410 1812.310 1704.000 ;
        RECT 1812.030 1700.270 1813.620 1700.410 ;
        RECT 1812.030 1700.000 1812.310 1700.270 ;
        RECT 1813.480 47.445 1813.620 1700.270 ;
        RECT 1813.410 47.075 1813.690 47.445 ;
        RECT 2452.810 47.075 2453.090 47.445 ;
        RECT 2452.880 2.400 2453.020 47.075 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
      LAYER via2 ;
        RECT 1813.410 47.120 1813.690 47.400 ;
        RECT 2452.810 47.120 2453.090 47.400 ;
      LAYER met3 ;
        RECT 1813.385 47.410 1813.715 47.425 ;
        RECT 2452.785 47.410 2453.115 47.425 ;
        RECT 1813.385 47.110 2453.115 47.410 ;
        RECT 1813.385 47.095 1813.715 47.110 ;
        RECT 2452.785 47.095 2453.115 47.110 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1817.070 1684.260 1817.390 1684.320 ;
        RECT 1820.750 1684.260 1821.070 1684.320 ;
        RECT 1817.070 1684.120 1821.070 1684.260 ;
        RECT 1817.070 1684.060 1817.390 1684.120 ;
        RECT 1820.750 1684.060 1821.070 1684.120 ;
        RECT 1820.750 20.980 1821.070 21.040 ;
        RECT 2470.730 20.980 2471.050 21.040 ;
        RECT 1820.750 20.840 2471.050 20.980 ;
        RECT 1820.750 20.780 1821.070 20.840 ;
        RECT 2470.730 20.780 2471.050 20.840 ;
      LAYER via ;
        RECT 1817.100 1684.060 1817.360 1684.320 ;
        RECT 1820.780 1684.060 1821.040 1684.320 ;
        RECT 1820.780 20.780 1821.040 21.040 ;
        RECT 2470.760 20.780 2471.020 21.040 ;
      LAYER met2 ;
        RECT 1817.090 1700.000 1817.370 1704.000 ;
        RECT 1817.160 1684.350 1817.300 1700.000 ;
        RECT 1817.100 1684.030 1817.360 1684.350 ;
        RECT 1820.780 1684.030 1821.040 1684.350 ;
        RECT 1820.840 21.070 1820.980 1684.030 ;
        RECT 1820.780 20.750 1821.040 21.070 ;
        RECT 2470.760 20.750 2471.020 21.070 ;
        RECT 2470.820 2.400 2470.960 20.750 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 0.300 ;
=======
      LAYER li1 ;
        RECT 1873.725 21.165 1873.895 23.715 ;
      LAYER mcon ;
        RECT 1873.725 23.545 1873.895 23.715 ;
      LAYER met1 ;
        RECT 1823.050 1677.460 1823.370 1677.520 ;
        RECT 1827.650 1677.460 1827.970 1677.520 ;
        RECT 1823.050 1677.320 1827.970 1677.460 ;
        RECT 1823.050 1677.260 1823.370 1677.320 ;
        RECT 1827.650 1677.260 1827.970 1677.320 ;
        RECT 1873.665 23.700 1873.955 23.745 ;
        RECT 1833.260 23.560 1873.955 23.700 ;
        RECT 1827.650 23.360 1827.970 23.420 ;
        RECT 1833.260 23.360 1833.400 23.560 ;
        RECT 1873.665 23.515 1873.955 23.560 ;
        RECT 1827.650 23.220 1833.400 23.360 ;
        RECT 1827.650 23.160 1827.970 23.220 ;
        RECT 1873.665 21.320 1873.955 21.365 ;
        RECT 2488.670 21.320 2488.990 21.380 ;
        RECT 1873.665 21.180 2488.990 21.320 ;
        RECT 1873.665 21.135 1873.955 21.180 ;
        RECT 2488.670 21.120 2488.990 21.180 ;
      LAYER via ;
        RECT 1823.080 1677.260 1823.340 1677.520 ;
        RECT 1827.680 1677.260 1827.940 1677.520 ;
        RECT 1827.680 23.160 1827.940 23.420 ;
        RECT 2488.700 21.120 2488.960 21.380 ;
      LAYER met2 ;
        RECT 1821.690 1700.410 1821.970 1704.000 ;
        RECT 1821.690 1700.270 1823.280 1700.410 ;
        RECT 1821.690 1700.000 1821.970 1700.270 ;
        RECT 1823.140 1677.550 1823.280 1700.270 ;
        RECT 1823.080 1677.230 1823.340 1677.550 ;
        RECT 1827.680 1677.230 1827.940 1677.550 ;
        RECT 1827.740 23.450 1827.880 1677.230 ;
        RECT 1827.680 23.130 1827.940 23.450 ;
        RECT 2488.700 21.090 2488.960 21.410 ;
        RECT 2488.760 2.400 2488.900 21.090 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 0.300 ;
=======
      LAYER met1 ;
        RECT 2506.150 21.660 2506.470 21.720 ;
        RECT 1873.280 21.520 2506.470 21.660 ;
        RECT 1827.190 21.320 1827.510 21.380 ;
        RECT 1873.280 21.320 1873.420 21.520 ;
        RECT 2506.150 21.460 2506.470 21.520 ;
        RECT 1827.190 21.180 1873.420 21.320 ;
        RECT 1827.190 21.120 1827.510 21.180 ;
      LAYER via ;
        RECT 1827.220 21.120 1827.480 21.380 ;
        RECT 2506.180 21.460 2506.440 21.720 ;
      LAYER met2 ;
        RECT 1826.750 1700.410 1827.030 1704.000 ;
        RECT 1826.750 1700.270 1827.420 1700.410 ;
        RECT 1826.750 1700.000 1827.030 1700.270 ;
        RECT 1827.280 21.410 1827.420 1700.270 ;
        RECT 2506.180 21.430 2506.440 21.750 ;
        RECT 1827.220 21.090 1827.480 21.410 ;
        RECT 2506.240 2.400 2506.380 21.430 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1831.330 1683.920 1831.650 1683.980 ;
        RECT 1834.550 1683.920 1834.870 1683.980 ;
        RECT 1831.330 1683.780 1834.870 1683.920 ;
        RECT 1831.330 1683.720 1831.650 1683.780 ;
        RECT 1834.550 1683.720 1834.870 1683.780 ;
        RECT 2524.090 22.000 2524.410 22.060 ;
        RECT 1870.520 21.860 2524.410 22.000 ;
        RECT 1833.170 21.660 1833.490 21.720 ;
        RECT 1870.520 21.660 1870.660 21.860 ;
        RECT 2524.090 21.800 2524.410 21.860 ;
        RECT 1833.170 21.520 1870.660 21.660 ;
        RECT 1833.170 21.460 1833.490 21.520 ;
      LAYER via ;
        RECT 1831.360 1683.720 1831.620 1683.980 ;
        RECT 1834.580 1683.720 1834.840 1683.980 ;
        RECT 1833.200 21.460 1833.460 21.720 ;
        RECT 2524.120 21.800 2524.380 22.060 ;
      LAYER met2 ;
        RECT 1831.350 1700.000 1831.630 1704.000 ;
        RECT 1831.420 1684.010 1831.560 1700.000 ;
        RECT 1831.360 1683.690 1831.620 1684.010 ;
        RECT 1834.580 1683.690 1834.840 1684.010 ;
        RECT 1834.640 109.890 1834.780 1683.690 ;
        RECT 1833.260 109.750 1834.780 109.890 ;
        RECT 1833.260 21.750 1833.400 109.750 ;
        RECT 2524.120 21.770 2524.380 22.090 ;
        RECT 1833.200 21.430 1833.460 21.750 ;
        RECT 2524.180 2.400 2524.320 21.770 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 0.300 ;
=======
      LAYER li1 ;
        RECT 1873.265 22.185 1873.435 27.115 ;
      LAYER mcon ;
        RECT 1873.265 26.945 1873.435 27.115 ;
      LAYER met1 ;
        RECT 1836.390 1683.920 1836.710 1683.980 ;
        RECT 1841.910 1683.920 1842.230 1683.980 ;
        RECT 1836.390 1683.780 1842.230 1683.920 ;
        RECT 1836.390 1683.720 1836.710 1683.780 ;
        RECT 1841.910 1683.720 1842.230 1683.780 ;
        RECT 1841.910 27.100 1842.230 27.160 ;
        RECT 1873.205 27.100 1873.495 27.145 ;
        RECT 1841.910 26.960 1873.495 27.100 ;
        RECT 1841.910 26.900 1842.230 26.960 ;
        RECT 1873.205 26.915 1873.495 26.960 ;
        RECT 1873.205 22.340 1873.495 22.385 ;
        RECT 2542.030 22.340 2542.350 22.400 ;
        RECT 1873.205 22.200 2542.350 22.340 ;
        RECT 1873.205 22.155 1873.495 22.200 ;
        RECT 2542.030 22.140 2542.350 22.200 ;
      LAYER via ;
        RECT 1836.420 1683.720 1836.680 1683.980 ;
        RECT 1841.940 1683.720 1842.200 1683.980 ;
        RECT 1841.940 26.900 1842.200 27.160 ;
        RECT 2542.060 22.140 2542.320 22.400 ;
      LAYER met2 ;
        RECT 1836.410 1700.000 1836.690 1704.000 ;
        RECT 1836.480 1684.010 1836.620 1700.000 ;
        RECT 1836.420 1683.690 1836.680 1684.010 ;
        RECT 1841.940 1683.690 1842.200 1684.010 ;
        RECT 1842.000 27.190 1842.140 1683.690 ;
        RECT 1841.940 26.870 1842.200 27.190 ;
        RECT 2542.060 22.110 2542.320 22.430 ;
        RECT 2542.120 2.400 2542.260 22.110 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 0.300 ;
=======
      LAYER met1 ;
        RECT 2559.970 22.680 2560.290 22.740 ;
        RECT 1870.060 22.540 2560.290 22.680 ;
        RECT 1841.450 22.000 1841.770 22.060 ;
        RECT 1870.060 22.000 1870.200 22.540 ;
        RECT 2559.970 22.480 2560.290 22.540 ;
        RECT 1841.450 21.860 1870.200 22.000 ;
        RECT 1841.450 21.800 1841.770 21.860 ;
      LAYER via ;
        RECT 1841.480 21.800 1841.740 22.060 ;
        RECT 2560.000 22.480 2560.260 22.740 ;
      LAYER met2 ;
        RECT 1841.010 1700.410 1841.290 1704.000 ;
        RECT 1841.010 1700.270 1841.680 1700.410 ;
        RECT 1841.010 1700.000 1841.290 1700.270 ;
        RECT 1841.540 22.090 1841.680 1700.270 ;
        RECT 2560.000 22.450 2560.260 22.770 ;
        RECT 1841.480 21.770 1841.740 22.090 ;
        RECT 2560.060 2.400 2560.200 22.450 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1846.050 1685.280 1846.370 1685.340 ;
        RECT 1848.810 1685.280 1849.130 1685.340 ;
        RECT 1846.050 1685.140 1849.130 1685.280 ;
        RECT 1846.050 1685.080 1846.370 1685.140 ;
        RECT 1848.810 1685.080 1849.130 1685.140 ;
        RECT 2577.910 23.020 2578.230 23.080 ;
        RECT 1869.600 22.880 2578.230 23.020 ;
        RECT 1848.810 22.340 1849.130 22.400 ;
        RECT 1869.600 22.340 1869.740 22.880 ;
        RECT 2577.910 22.820 2578.230 22.880 ;
        RECT 1848.810 22.200 1869.740 22.340 ;
        RECT 1848.810 22.140 1849.130 22.200 ;
      LAYER via ;
        RECT 1846.080 1685.080 1846.340 1685.340 ;
        RECT 1848.840 1685.080 1849.100 1685.340 ;
        RECT 1848.840 22.140 1849.100 22.400 ;
        RECT 2577.940 22.820 2578.200 23.080 ;
      LAYER met2 ;
        RECT 1846.070 1700.000 1846.350 1704.000 ;
        RECT 1846.140 1685.370 1846.280 1700.000 ;
        RECT 1846.080 1685.050 1846.340 1685.370 ;
        RECT 1848.840 1685.050 1849.100 1685.370 ;
        RECT 1848.900 22.430 1849.040 1685.050 ;
        RECT 2577.940 22.790 2578.200 23.110 ;
        RECT 1848.840 22.110 1849.100 22.430 ;
        RECT 2578.000 2.400 2578.140 22.790 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 0.300 ;
=======
      LAYER met1 ;
        RECT 813.810 50.560 814.130 50.620 ;
        RECT 1367.650 50.560 1367.970 50.620 ;
        RECT 813.810 50.420 1367.970 50.560 ;
        RECT 813.810 50.360 814.130 50.420 ;
        RECT 1367.650 50.360 1367.970 50.420 ;
      LAYER via ;
        RECT 813.840 50.360 814.100 50.620 ;
        RECT 1367.680 50.360 1367.940 50.620 ;
      LAYER met2 ;
        RECT 1368.590 1700.410 1368.870 1704.000 ;
        RECT 1367.740 1700.270 1368.870 1700.410 ;
        RECT 1367.740 50.650 1367.880 1700.270 ;
        RECT 1368.590 1700.000 1368.870 1700.270 ;
        RECT 813.840 50.330 814.100 50.650 ;
        RECT 1367.680 50.330 1367.940 50.650 ;
        RECT 813.900 3.130 814.040 50.330 ;
        RECT 811.600 2.990 814.040 3.130 ;
        RECT 811.600 2.400 811.740 2.990 ;
        RECT 811.390 -4.800 811.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 0.300 ;
=======
      LAYER li1 ;
        RECT 1869.125 22.355 1869.295 22.695 ;
        RECT 1869.125 22.185 1870.675 22.355 ;
      LAYER mcon ;
        RECT 1869.125 22.525 1869.295 22.695 ;
        RECT 1870.505 22.185 1870.675 22.355 ;
      LAYER met1 ;
        RECT 1850.650 1685.620 1850.970 1685.680 ;
        RECT 1854.790 1685.620 1855.110 1685.680 ;
        RECT 1850.650 1685.480 1855.110 1685.620 ;
        RECT 1850.650 1685.420 1850.970 1685.480 ;
        RECT 1854.790 1685.420 1855.110 1685.480 ;
        RECT 1874.570 23.360 1874.890 23.420 ;
        RECT 2595.390 23.360 2595.710 23.420 ;
        RECT 1874.570 23.220 2595.710 23.360 ;
        RECT 1874.570 23.160 1874.890 23.220 ;
        RECT 2595.390 23.160 2595.710 23.220 ;
        RECT 1854.790 22.680 1855.110 22.740 ;
        RECT 1869.065 22.680 1869.355 22.725 ;
        RECT 1854.790 22.540 1869.355 22.680 ;
        RECT 1854.790 22.480 1855.110 22.540 ;
        RECT 1869.065 22.495 1869.355 22.540 ;
        RECT 1870.445 22.340 1870.735 22.385 ;
        RECT 1872.730 22.340 1873.050 22.400 ;
        RECT 1870.445 22.200 1873.050 22.340 ;
        RECT 1870.445 22.155 1870.735 22.200 ;
        RECT 1872.730 22.140 1873.050 22.200 ;
      LAYER via ;
        RECT 1850.680 1685.420 1850.940 1685.680 ;
        RECT 1854.820 1685.420 1855.080 1685.680 ;
        RECT 1874.600 23.160 1874.860 23.420 ;
        RECT 2595.420 23.160 2595.680 23.420 ;
        RECT 1854.820 22.480 1855.080 22.740 ;
        RECT 1872.760 22.140 1873.020 22.400 ;
      LAYER met2 ;
        RECT 1850.670 1700.000 1850.950 1704.000 ;
        RECT 1850.740 1685.710 1850.880 1700.000 ;
        RECT 1850.680 1685.390 1850.940 1685.710 ;
        RECT 1854.820 1685.390 1855.080 1685.710 ;
        RECT 1854.880 22.770 1855.020 1685.390 ;
        RECT 1874.600 23.130 1874.860 23.450 ;
        RECT 2595.420 23.130 2595.680 23.450 ;
        RECT 1874.660 22.850 1874.800 23.130 ;
        RECT 1854.820 22.450 1855.080 22.770 ;
        RECT 1872.820 22.710 1874.800 22.850 ;
        RECT 1872.820 22.430 1872.960 22.710 ;
        RECT 1872.760 22.110 1873.020 22.430 ;
        RECT 2595.480 2.400 2595.620 23.130 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 0.300 ;
=======
      LAYER met1 ;
        RECT 2613.330 23.700 2613.650 23.760 ;
        RECT 1874.200 23.560 2613.650 23.700 ;
        RECT 1855.250 23.360 1855.570 23.420 ;
        RECT 1874.200 23.360 1874.340 23.560 ;
        RECT 2613.330 23.500 2613.650 23.560 ;
        RECT 1855.250 23.220 1874.340 23.360 ;
        RECT 1855.250 23.160 1855.570 23.220 ;
      LAYER via ;
        RECT 1855.280 23.160 1855.540 23.420 ;
        RECT 2613.360 23.500 2613.620 23.760 ;
      LAYER met2 ;
        RECT 1855.270 1700.000 1855.550 1704.000 ;
        RECT 1855.340 23.450 1855.480 1700.000 ;
        RECT 2613.360 23.470 2613.620 23.790 ;
        RECT 1855.280 23.130 1855.540 23.450 ;
        RECT 2613.420 2.400 2613.560 23.470 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 0.300 ;
=======
      LAYER li1 ;
        RECT 1880.625 27.285 1881.715 27.455 ;
        RECT 1880.625 26.945 1880.795 27.285 ;
      LAYER mcon ;
        RECT 1881.545 27.285 1881.715 27.455 ;
      LAYER met1 ;
        RECT 1860.310 1686.640 1860.630 1686.700 ;
        RECT 1862.610 1686.640 1862.930 1686.700 ;
        RECT 1860.310 1686.500 1862.930 1686.640 ;
        RECT 1860.310 1686.440 1860.630 1686.500 ;
        RECT 1862.610 1686.440 1862.930 1686.500 ;
        RECT 1881.485 27.440 1881.775 27.485 ;
        RECT 2631.270 27.440 2631.590 27.500 ;
        RECT 1881.485 27.300 2631.590 27.440 ;
        RECT 1881.485 27.255 1881.775 27.300 ;
        RECT 2631.270 27.240 2631.590 27.300 ;
        RECT 1880.565 27.100 1880.855 27.145 ;
        RECT 1873.740 26.960 1880.855 27.100 ;
        RECT 1862.610 26.760 1862.930 26.820 ;
        RECT 1873.740 26.760 1873.880 26.960 ;
        RECT 1880.565 26.915 1880.855 26.960 ;
        RECT 1862.610 26.620 1873.880 26.760 ;
        RECT 1862.610 26.560 1862.930 26.620 ;
      LAYER via ;
        RECT 1860.340 1686.440 1860.600 1686.700 ;
        RECT 1862.640 1686.440 1862.900 1686.700 ;
        RECT 2631.300 27.240 2631.560 27.500 ;
        RECT 1862.640 26.560 1862.900 26.820 ;
      LAYER met2 ;
        RECT 1860.330 1700.000 1860.610 1704.000 ;
        RECT 1860.400 1686.730 1860.540 1700.000 ;
        RECT 1860.340 1686.410 1860.600 1686.730 ;
        RECT 1862.640 1686.410 1862.900 1686.730 ;
        RECT 1862.700 26.850 1862.840 1686.410 ;
        RECT 2631.300 27.210 2631.560 27.530 ;
        RECT 1862.640 26.530 1862.900 26.850 ;
        RECT 2631.360 2.400 2631.500 27.210 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1864.910 1685.620 1865.230 1685.680 ;
        RECT 1869.510 1685.620 1869.830 1685.680 ;
        RECT 1864.910 1685.480 1869.830 1685.620 ;
        RECT 1864.910 1685.420 1865.230 1685.480 ;
        RECT 1869.510 1685.420 1869.830 1685.480 ;
        RECT 1869.510 27.440 1869.830 27.500 ;
        RECT 1869.510 27.300 1881.240 27.440 ;
        RECT 1869.510 27.240 1869.830 27.300 ;
        RECT 1881.100 27.100 1881.240 27.300 ;
        RECT 2649.210 27.100 2649.530 27.160 ;
        RECT 1881.100 26.960 2649.530 27.100 ;
        RECT 2649.210 26.900 2649.530 26.960 ;
      LAYER via ;
        RECT 1864.940 1685.420 1865.200 1685.680 ;
        RECT 1869.540 1685.420 1869.800 1685.680 ;
        RECT 1869.540 27.240 1869.800 27.500 ;
        RECT 2649.240 26.900 2649.500 27.160 ;
      LAYER met2 ;
        RECT 1864.930 1700.000 1865.210 1704.000 ;
        RECT 1865.000 1685.710 1865.140 1700.000 ;
        RECT 1864.940 1685.390 1865.200 1685.710 ;
        RECT 1869.540 1685.390 1869.800 1685.710 ;
        RECT 1869.600 27.530 1869.740 1685.390 ;
        RECT 1869.540 27.210 1869.800 27.530 ;
        RECT 2649.240 26.870 2649.500 27.190 ;
        RECT 2649.300 2.400 2649.440 26.870 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1870.890 1685.280 1871.210 1685.340 ;
        RECT 1875.490 1685.280 1875.810 1685.340 ;
        RECT 1870.890 1685.140 1875.810 1685.280 ;
        RECT 1870.890 1685.080 1871.210 1685.140 ;
        RECT 1875.490 1685.080 1875.810 1685.140 ;
        RECT 1875.490 26.760 1875.810 26.820 ;
        RECT 2667.150 26.760 2667.470 26.820 ;
        RECT 1875.490 26.620 2667.470 26.760 ;
        RECT 1875.490 26.560 1875.810 26.620 ;
        RECT 2667.150 26.560 2667.470 26.620 ;
      LAYER via ;
        RECT 1870.920 1685.080 1871.180 1685.340 ;
        RECT 1875.520 1685.080 1875.780 1685.340 ;
        RECT 1875.520 26.560 1875.780 26.820 ;
        RECT 2667.180 26.560 2667.440 26.820 ;
      LAYER met2 ;
        RECT 1869.990 1700.410 1870.270 1704.000 ;
        RECT 1869.990 1700.270 1871.120 1700.410 ;
        RECT 1869.990 1700.000 1870.270 1700.270 ;
        RECT 1870.980 1685.370 1871.120 1700.270 ;
        RECT 1870.920 1685.050 1871.180 1685.370 ;
        RECT 1875.520 1685.050 1875.780 1685.370 ;
        RECT 1875.580 26.850 1875.720 1685.050 ;
        RECT 1875.520 26.530 1875.780 26.850 ;
        RECT 2667.180 26.530 2667.440 26.850 ;
        RECT 2667.240 2.400 2667.380 26.530 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 0.300 ;
=======
      LAYER li1 ;
        RECT 1916.965 26.265 1918.055 26.435 ;
        RECT 1916.965 25.245 1917.135 26.265 ;
      LAYER mcon ;
        RECT 1917.885 26.265 1918.055 26.435 ;
      LAYER met1 ;
        RECT 1917.825 26.420 1918.115 26.465 ;
        RECT 2684.630 26.420 2684.950 26.480 ;
        RECT 1917.825 26.280 2684.950 26.420 ;
        RECT 1917.825 26.235 1918.115 26.280 ;
        RECT 2684.630 26.220 2684.950 26.280 ;
        RECT 1875.950 25.400 1876.270 25.460 ;
        RECT 1916.905 25.400 1917.195 25.445 ;
        RECT 1875.950 25.260 1917.195 25.400 ;
        RECT 1875.950 25.200 1876.270 25.260 ;
        RECT 1916.905 25.215 1917.195 25.260 ;
      LAYER via ;
        RECT 2684.660 26.220 2684.920 26.480 ;
        RECT 1875.980 25.200 1876.240 25.460 ;
      LAYER met2 ;
        RECT 1874.590 1700.410 1874.870 1704.000 ;
        RECT 1874.590 1700.270 1876.180 1700.410 ;
        RECT 1874.590 1700.000 1874.870 1700.270 ;
        RECT 1876.040 25.490 1876.180 1700.270 ;
        RECT 2684.660 26.190 2684.920 26.510 ;
        RECT 1875.980 25.170 1876.240 25.490 ;
        RECT 2684.720 2.400 2684.860 26.190 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1879.630 1686.640 1879.950 1686.700 ;
        RECT 1882.850 1686.640 1883.170 1686.700 ;
        RECT 1879.630 1686.500 1883.170 1686.640 ;
        RECT 1879.630 1686.440 1879.950 1686.500 ;
        RECT 1882.850 1686.440 1883.170 1686.500 ;
        RECT 1882.850 1608.920 1883.170 1609.180 ;
        RECT 1882.940 1608.160 1883.080 1608.920 ;
        RECT 1882.850 1607.900 1883.170 1608.160 ;
        RECT 1882.850 26.420 1883.170 26.480 ;
        RECT 1882.850 26.280 1917.580 26.420 ;
        RECT 1882.850 26.220 1883.170 26.280 ;
        RECT 1917.440 26.080 1917.580 26.280 ;
        RECT 2702.570 26.080 2702.890 26.140 ;
        RECT 1917.440 25.940 2702.890 26.080 ;
        RECT 2702.570 25.880 2702.890 25.940 ;
      LAYER via ;
        RECT 1879.660 1686.440 1879.920 1686.700 ;
        RECT 1882.880 1686.440 1883.140 1686.700 ;
        RECT 1882.880 1608.920 1883.140 1609.180 ;
        RECT 1882.880 1607.900 1883.140 1608.160 ;
        RECT 1882.880 26.220 1883.140 26.480 ;
        RECT 2702.600 25.880 2702.860 26.140 ;
      LAYER met2 ;
        RECT 1879.650 1700.000 1879.930 1704.000 ;
        RECT 1879.720 1686.730 1879.860 1700.000 ;
        RECT 1879.660 1686.410 1879.920 1686.730 ;
        RECT 1882.880 1686.410 1883.140 1686.730 ;
        RECT 1882.940 1609.210 1883.080 1686.410 ;
        RECT 1882.880 1608.890 1883.140 1609.210 ;
        RECT 1882.880 1607.870 1883.140 1608.190 ;
        RECT 1882.940 26.510 1883.080 1607.870 ;
        RECT 1882.880 26.190 1883.140 26.510 ;
        RECT 2702.600 25.850 2702.860 26.170 ;
        RECT 2702.660 2.400 2702.800 25.850 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 0.300 ;
=======
      LAYER li1 ;
        RECT 1916.505 25.075 1916.675 26.095 ;
        RECT 1917.425 25.585 1918.975 25.755 ;
        RECT 1917.425 25.075 1917.595 25.585 ;
        RECT 1916.505 24.905 1917.595 25.075 ;
      LAYER mcon ;
        RECT 1916.505 25.925 1916.675 26.095 ;
        RECT 1918.805 25.585 1918.975 25.755 ;
      LAYER met1 ;
        RECT 1884.230 1685.280 1884.550 1685.340 ;
        RECT 1890.210 1685.280 1890.530 1685.340 ;
        RECT 1884.230 1685.140 1890.530 1685.280 ;
        RECT 1884.230 1685.080 1884.550 1685.140 ;
        RECT 1890.210 1685.080 1890.530 1685.140 ;
        RECT 1890.210 26.080 1890.530 26.140 ;
        RECT 1916.445 26.080 1916.735 26.125 ;
        RECT 1890.210 25.940 1916.735 26.080 ;
        RECT 1890.210 25.880 1890.530 25.940 ;
        RECT 1916.445 25.895 1916.735 25.940 ;
        RECT 1918.745 25.740 1919.035 25.785 ;
        RECT 2720.510 25.740 2720.830 25.800 ;
        RECT 1918.745 25.600 2720.830 25.740 ;
        RECT 1918.745 25.555 1919.035 25.600 ;
        RECT 2720.510 25.540 2720.830 25.600 ;
      LAYER via ;
        RECT 1884.260 1685.080 1884.520 1685.340 ;
        RECT 1890.240 1685.080 1890.500 1685.340 ;
        RECT 1890.240 25.880 1890.500 26.140 ;
        RECT 2720.540 25.540 2720.800 25.800 ;
      LAYER met2 ;
        RECT 1884.250 1700.000 1884.530 1704.000 ;
        RECT 1884.320 1685.370 1884.460 1700.000 ;
        RECT 1884.260 1685.050 1884.520 1685.370 ;
        RECT 1890.240 1685.050 1890.500 1685.370 ;
        RECT 1890.300 26.170 1890.440 1685.050 ;
        RECT 1890.240 25.850 1890.500 26.170 ;
        RECT 2720.540 25.510 2720.800 25.830 ;
        RECT 2720.600 2.400 2720.740 25.510 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 0.300 ;
=======
      LAYER met1 ;
        RECT 1883.770 1685.620 1884.090 1685.680 ;
        RECT 1887.910 1685.620 1888.230 1685.680 ;
        RECT 1883.770 1685.480 1888.230 1685.620 ;
        RECT 1883.770 1685.420 1884.090 1685.480 ;
        RECT 1887.910 1685.420 1888.230 1685.480 ;
        RECT 1883.770 1631.900 1884.090 1631.960 ;
        RECT 1889.750 1631.900 1890.070 1631.960 ;
        RECT 1883.770 1631.760 1890.070 1631.900 ;
        RECT 1883.770 1631.700 1884.090 1631.760 ;
        RECT 1889.750 1631.700 1890.070 1631.760 ;
      LAYER via ;
        RECT 1883.800 1685.420 1884.060 1685.680 ;
        RECT 1887.940 1685.420 1888.200 1685.680 ;
        RECT 1883.800 1631.700 1884.060 1631.960 ;
        RECT 1889.780 1631.700 1890.040 1631.960 ;
      LAYER met2 ;
        RECT 1889.310 1700.410 1889.590 1704.000 ;
        RECT 1888.000 1700.270 1889.590 1700.410 ;
        RECT 1888.000 1685.710 1888.140 1700.270 ;
        RECT 1889.310 1700.000 1889.590 1700.270 ;
        RECT 1883.800 1685.390 1884.060 1685.710 ;
        RECT 1887.940 1685.390 1888.200 1685.710 ;
        RECT 1883.860 1631.990 1884.000 1685.390 ;
        RECT 1883.800 1631.670 1884.060 1631.990 ;
        RECT 1889.780 1631.670 1890.040 1631.990 ;
        RECT 1889.840 27.045 1889.980 1631.670 ;
        RECT 1889.770 26.675 1890.050 27.045 ;
        RECT 2738.470 26.675 2738.750 27.045 ;
        RECT 2738.540 2.400 2738.680 26.675 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
      LAYER via2 ;
        RECT 1889.770 26.720 1890.050 27.000 ;
        RECT 2738.470 26.720 2738.750 27.000 ;
      LAYER met3 ;
        RECT 1889.745 27.010 1890.075 27.025 ;
        RECT 2738.445 27.010 2738.775 27.025 ;
        RECT 1889.745 26.710 2738.775 27.010 ;
        RECT 1889.745 26.695 1890.075 26.710 ;
        RECT 2738.445 26.695 2738.775 26.710 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 0.300 ;
=======
      LAYER met1 ;
        RECT 1891.130 1632.240 1891.450 1632.300 ;
        RECT 1897.110 1632.240 1897.430 1632.300 ;
        RECT 1891.130 1632.100 1897.430 1632.240 ;
        RECT 1891.130 1632.040 1891.450 1632.100 ;
        RECT 1897.110 1632.040 1897.430 1632.100 ;
      LAYER via ;
        RECT 1891.160 1632.040 1891.420 1632.300 ;
        RECT 1897.140 1632.040 1897.400 1632.300 ;
      LAYER met2 ;
        RECT 1893.910 1700.410 1894.190 1704.000 ;
        RECT 1893.060 1700.270 1894.190 1700.410 ;
        RECT 1893.060 1688.850 1893.200 1700.270 ;
        RECT 1893.910 1700.000 1894.190 1700.270 ;
        RECT 1891.220 1688.710 1893.200 1688.850 ;
        RECT 1891.220 1632.330 1891.360 1688.710 ;
        RECT 1891.160 1632.010 1891.420 1632.330 ;
        RECT 1897.140 1632.010 1897.400 1632.330 ;
        RECT 1897.200 26.365 1897.340 1632.010 ;
        RECT 1897.130 25.995 1897.410 26.365 ;
        RECT 2755.950 25.995 2756.230 26.365 ;
        RECT 2756.020 2.400 2756.160 25.995 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
      LAYER via2 ;
        RECT 1897.130 26.040 1897.410 26.320 ;
        RECT 2755.950 26.040 2756.230 26.320 ;
      LAYER met3 ;
        RECT 1897.105 26.330 1897.435 26.345 ;
        RECT 2755.925 26.330 2756.255 26.345 ;
        RECT 1897.105 26.030 2756.255 26.330 ;
        RECT 1897.105 26.015 1897.435 26.030 ;
        RECT 2755.925 26.015 2756.255 26.030 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 0.300 ;
=======
      LAYER met1 ;
        RECT 834.510 50.220 834.830 50.280 ;
        RECT 1374.550 50.220 1374.870 50.280 ;
        RECT 834.510 50.080 1374.870 50.220 ;
        RECT 834.510 50.020 834.830 50.080 ;
        RECT 1374.550 50.020 1374.870 50.080 ;
        RECT 829.450 2.960 829.770 3.020 ;
        RECT 834.510 2.960 834.830 3.020 ;
        RECT 829.450 2.820 834.830 2.960 ;
        RECT 829.450 2.760 829.770 2.820 ;
        RECT 834.510 2.760 834.830 2.820 ;
      LAYER via ;
        RECT 834.540 50.020 834.800 50.280 ;
        RECT 1374.580 50.020 1374.840 50.280 ;
        RECT 829.480 2.760 829.740 3.020 ;
        RECT 834.540 2.760 834.800 3.020 ;
      LAYER met2 ;
        RECT 1373.650 1700.410 1373.930 1704.000 ;
        RECT 1373.650 1700.270 1374.780 1700.410 ;
        RECT 1373.650 1700.000 1373.930 1700.270 ;
        RECT 1374.640 50.310 1374.780 1700.270 ;
        RECT 834.540 49.990 834.800 50.310 ;
        RECT 1374.580 49.990 1374.840 50.310 ;
        RECT 834.600 3.050 834.740 49.990 ;
        RECT 829.480 2.730 829.740 3.050 ;
        RECT 834.540 2.730 834.800 3.050 ;
        RECT 829.540 2.400 829.680 2.730 ;
        RECT 829.330 -4.800 829.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1899.870 1685.620 1900.190 1685.680 ;
        RECT 1903.090 1685.620 1903.410 1685.680 ;
        RECT 1899.870 1685.480 1903.410 1685.620 ;
        RECT 1899.870 1685.420 1900.190 1685.480 ;
        RECT 1903.090 1685.420 1903.410 1685.480 ;
        RECT 2773.870 25.400 2774.190 25.460 ;
        RECT 1942.280 25.260 2774.190 25.400 ;
        RECT 1903.090 25.060 1903.410 25.120 ;
        RECT 1942.280 25.060 1942.420 25.260 ;
        RECT 2773.870 25.200 2774.190 25.260 ;
        RECT 1903.090 24.920 1942.420 25.060 ;
        RECT 1903.090 24.860 1903.410 24.920 ;
      LAYER via ;
        RECT 1899.900 1685.420 1900.160 1685.680 ;
        RECT 1903.120 1685.420 1903.380 1685.680 ;
        RECT 1903.120 24.860 1903.380 25.120 ;
        RECT 2773.900 25.200 2774.160 25.460 ;
      LAYER met2 ;
        RECT 1898.970 1700.410 1899.250 1704.000 ;
        RECT 1898.970 1700.270 1900.100 1700.410 ;
        RECT 1898.970 1700.000 1899.250 1700.270 ;
        RECT 1899.960 1685.710 1900.100 1700.270 ;
        RECT 1899.900 1685.390 1900.160 1685.710 ;
        RECT 1903.120 1685.390 1903.380 1685.710 ;
        RECT 1903.180 25.150 1903.320 1685.390 ;
        RECT 2773.900 25.170 2774.160 25.490 ;
        RECT 1903.120 24.830 1903.380 25.150 ;
        RECT 2773.960 2.400 2774.100 25.170 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1898.030 1686.300 1898.350 1686.360 ;
        RECT 1903.550 1686.300 1903.870 1686.360 ;
        RECT 1898.030 1686.160 1903.870 1686.300 ;
        RECT 1898.030 1686.100 1898.350 1686.160 ;
        RECT 1903.550 1686.100 1903.870 1686.160 ;
        RECT 1897.570 1631.900 1897.890 1631.960 ;
        RECT 1903.550 1631.900 1903.870 1631.960 ;
        RECT 1897.570 1631.760 1903.870 1631.900 ;
        RECT 1897.570 1631.700 1897.890 1631.760 ;
        RECT 1903.550 1631.700 1903.870 1631.760 ;
      LAYER via ;
        RECT 1898.060 1686.100 1898.320 1686.360 ;
        RECT 1903.580 1686.100 1903.840 1686.360 ;
        RECT 1897.600 1631.700 1897.860 1631.960 ;
        RECT 1903.580 1631.700 1903.840 1631.960 ;
      LAYER met2 ;
        RECT 1903.570 1700.000 1903.850 1704.000 ;
        RECT 1903.640 1686.390 1903.780 1700.000 ;
        RECT 1898.060 1686.070 1898.320 1686.390 ;
        RECT 1903.580 1686.070 1903.840 1686.390 ;
        RECT 1898.120 1684.770 1898.260 1686.070 ;
        RECT 1897.660 1684.630 1898.260 1684.770 ;
        RECT 1897.660 1631.990 1897.800 1684.630 ;
        RECT 1897.600 1631.670 1897.860 1631.990 ;
        RECT 1903.580 1631.670 1903.840 1631.990 ;
        RECT 1903.640 25.685 1903.780 1631.670 ;
        RECT 1903.570 25.315 1903.850 25.685 ;
        RECT 2791.830 25.315 2792.110 25.685 ;
        RECT 2791.900 2.400 2792.040 25.315 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
      LAYER via2 ;
        RECT 1903.570 25.360 1903.850 25.640 ;
        RECT 2791.830 25.360 2792.110 25.640 ;
      LAYER met3 ;
        RECT 1903.545 25.650 1903.875 25.665 ;
        RECT 2791.805 25.650 2792.135 25.665 ;
        RECT 1903.545 25.350 2792.135 25.650 ;
        RECT 1903.545 25.335 1903.875 25.350 ;
        RECT 2791.805 25.335 2792.135 25.350 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1908.610 1684.260 1908.930 1684.320 ;
        RECT 1910.910 1684.260 1911.230 1684.320 ;
        RECT 1908.610 1684.120 1911.230 1684.260 ;
        RECT 1908.610 1684.060 1908.930 1684.120 ;
        RECT 1910.910 1684.060 1911.230 1684.120 ;
        RECT 1910.910 25.740 1911.230 25.800 ;
        RECT 1918.270 25.740 1918.590 25.800 ;
        RECT 1910.910 25.600 1918.590 25.740 ;
        RECT 1910.910 25.540 1911.230 25.600 ;
        RECT 1918.270 25.540 1918.590 25.600 ;
        RECT 2809.750 25.060 2810.070 25.120 ;
        RECT 1942.740 24.920 2810.070 25.060 ;
        RECT 1919.650 24.380 1919.970 24.440 ;
        RECT 1942.740 24.380 1942.880 24.920 ;
        RECT 2809.750 24.860 2810.070 24.920 ;
        RECT 1919.650 24.240 1942.880 24.380 ;
        RECT 1919.650 24.180 1919.970 24.240 ;
      LAYER via ;
        RECT 1908.640 1684.060 1908.900 1684.320 ;
        RECT 1910.940 1684.060 1911.200 1684.320 ;
        RECT 1910.940 25.540 1911.200 25.800 ;
        RECT 1918.300 25.540 1918.560 25.800 ;
        RECT 1919.680 24.180 1919.940 24.440 ;
        RECT 2809.780 24.860 2810.040 25.120 ;
      LAYER met2 ;
        RECT 1908.630 1700.000 1908.910 1704.000 ;
        RECT 1908.700 1684.350 1908.840 1700.000 ;
        RECT 1908.640 1684.030 1908.900 1684.350 ;
        RECT 1910.940 1684.030 1911.200 1684.350 ;
        RECT 1911.000 25.830 1911.140 1684.030 ;
        RECT 1910.940 25.510 1911.200 25.830 ;
        RECT 1918.300 25.510 1918.560 25.830 ;
        RECT 1918.360 24.890 1918.500 25.510 ;
        RECT 1918.360 24.750 1919.880 24.890 ;
        RECT 2809.780 24.830 2810.040 25.150 ;
        RECT 1919.740 24.470 1919.880 24.750 ;
        RECT 1919.680 24.150 1919.940 24.470 ;
        RECT 2809.840 2.400 2809.980 24.830 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 0.300 ;
=======
      LAYER li1 ;
        RECT 1941.805 24.735 1941.975 25.415 ;
        RECT 1941.805 24.565 1943.815 24.735 ;
      LAYER mcon ;
        RECT 1941.805 25.245 1941.975 25.415 ;
        RECT 1943.645 24.565 1943.815 24.735 ;
      LAYER met1 ;
        RECT 1913.210 1685.620 1913.530 1685.680 ;
        RECT 1917.810 1685.620 1918.130 1685.680 ;
        RECT 1913.210 1685.480 1918.130 1685.620 ;
        RECT 1913.210 1685.420 1913.530 1685.480 ;
        RECT 1917.810 1685.420 1918.130 1685.480 ;
        RECT 1917.810 25.400 1918.130 25.460 ;
        RECT 1941.745 25.400 1942.035 25.445 ;
        RECT 1917.810 25.260 1942.035 25.400 ;
        RECT 1917.810 25.200 1918.130 25.260 ;
        RECT 1941.745 25.215 1942.035 25.260 ;
        RECT 1943.585 24.720 1943.875 24.765 ;
        RECT 2827.690 24.720 2828.010 24.780 ;
        RECT 1943.585 24.580 2828.010 24.720 ;
        RECT 1943.585 24.535 1943.875 24.580 ;
        RECT 2827.690 24.520 2828.010 24.580 ;
      LAYER via ;
        RECT 1913.240 1685.420 1913.500 1685.680 ;
        RECT 1917.840 1685.420 1918.100 1685.680 ;
        RECT 1917.840 25.200 1918.100 25.460 ;
        RECT 2827.720 24.520 2827.980 24.780 ;
      LAYER met2 ;
        RECT 1913.230 1700.000 1913.510 1704.000 ;
        RECT 1913.300 1685.710 1913.440 1700.000 ;
        RECT 1913.240 1685.390 1913.500 1685.710 ;
        RECT 1917.840 1685.390 1918.100 1685.710 ;
        RECT 1917.900 25.490 1918.040 1685.390 ;
        RECT 1917.840 25.170 1918.100 25.490 ;
        RECT 2827.720 24.490 2827.980 24.810 ;
        RECT 2827.780 2.400 2827.920 24.490 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 0.300 ;
=======
      LAYER li1 ;
        RECT 1935.825 23.885 1935.995 24.735 ;
        RECT 1941.345 24.395 1941.515 24.735 ;
        RECT 1941.345 24.225 1943.355 24.395 ;
      LAYER mcon ;
        RECT 1935.825 24.565 1935.995 24.735 ;
        RECT 1941.345 24.565 1941.515 24.735 ;
        RECT 1943.185 24.225 1943.355 24.395 ;
      LAYER met1 ;
        RECT 1918.270 1686.300 1918.590 1686.360 ;
        RECT 1924.250 1686.300 1924.570 1686.360 ;
        RECT 1918.270 1686.160 1924.570 1686.300 ;
        RECT 1918.270 1686.100 1918.590 1686.160 ;
        RECT 1924.250 1686.100 1924.570 1686.160 ;
        RECT 1935.765 24.720 1936.055 24.765 ;
        RECT 1941.285 24.720 1941.575 24.765 ;
        RECT 1935.765 24.580 1941.575 24.720 ;
        RECT 1935.765 24.535 1936.055 24.580 ;
        RECT 1941.285 24.535 1941.575 24.580 ;
        RECT 1943.125 24.380 1943.415 24.425 ;
        RECT 2845.170 24.380 2845.490 24.440 ;
        RECT 1943.125 24.240 2845.490 24.380 ;
        RECT 1943.125 24.195 1943.415 24.240 ;
        RECT 2845.170 24.180 2845.490 24.240 ;
        RECT 1924.250 24.040 1924.570 24.100 ;
        RECT 1935.765 24.040 1936.055 24.085 ;
        RECT 1924.250 23.900 1936.055 24.040 ;
        RECT 1924.250 23.840 1924.570 23.900 ;
        RECT 1935.765 23.855 1936.055 23.900 ;
      LAYER via ;
        RECT 1918.300 1686.100 1918.560 1686.360 ;
        RECT 1924.280 1686.100 1924.540 1686.360 ;
        RECT 2845.200 24.180 2845.460 24.440 ;
        RECT 1924.280 23.840 1924.540 24.100 ;
      LAYER met2 ;
        RECT 1918.290 1700.000 1918.570 1704.000 ;
        RECT 1918.360 1686.390 1918.500 1700.000 ;
        RECT 1918.300 1686.070 1918.560 1686.390 ;
        RECT 1924.280 1686.070 1924.540 1686.390 ;
        RECT 1924.340 24.130 1924.480 1686.070 ;
        RECT 2845.200 24.150 2845.460 24.470 ;
        RECT 1924.280 23.810 1924.540 24.130 ;
        RECT 2845.260 2.400 2845.400 24.150 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1919.190 1684.260 1919.510 1684.320 ;
        RECT 1922.870 1684.260 1923.190 1684.320 ;
        RECT 1919.190 1684.120 1923.190 1684.260 ;
        RECT 1919.190 1684.060 1919.510 1684.120 ;
        RECT 1922.870 1684.060 1923.190 1684.120 ;
        RECT 1919.190 1631.900 1919.510 1631.960 ;
        RECT 1923.790 1631.900 1924.110 1631.960 ;
        RECT 1919.190 1631.760 1924.110 1631.900 ;
        RECT 1919.190 1631.700 1919.510 1631.760 ;
        RECT 1923.790 1631.700 1924.110 1631.760 ;
      LAYER via ;
        RECT 1919.220 1684.060 1919.480 1684.320 ;
        RECT 1922.900 1684.060 1923.160 1684.320 ;
        RECT 1919.220 1631.700 1919.480 1631.960 ;
        RECT 1923.820 1631.700 1924.080 1631.960 ;
      LAYER met2 ;
        RECT 1922.890 1700.000 1923.170 1704.000 ;
        RECT 1922.960 1684.350 1923.100 1700.000 ;
        RECT 1919.220 1684.030 1919.480 1684.350 ;
        RECT 1922.900 1684.030 1923.160 1684.350 ;
        RECT 1919.280 1631.990 1919.420 1684.030 ;
        RECT 1919.220 1631.670 1919.480 1631.990 ;
        RECT 1923.820 1631.670 1924.080 1631.990 ;
        RECT 1923.880 25.005 1924.020 1631.670 ;
        RECT 1923.810 24.635 1924.090 25.005 ;
        RECT 2863.130 24.635 2863.410 25.005 ;
        RECT 2863.200 2.400 2863.340 24.635 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
      LAYER via2 ;
        RECT 1923.810 24.680 1924.090 24.960 ;
        RECT 2863.130 24.680 2863.410 24.960 ;
      LAYER met3 ;
        RECT 1923.785 24.970 1924.115 24.985 ;
        RECT 2863.105 24.970 2863.435 24.985 ;
        RECT 1923.785 24.670 2863.435 24.970 ;
        RECT 1923.785 24.655 1924.115 24.670 ;
        RECT 2863.105 24.655 2863.435 24.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1927.930 1684.260 1928.250 1684.320 ;
        RECT 1931.150 1684.260 1931.470 1684.320 ;
        RECT 1927.930 1684.120 1931.470 1684.260 ;
        RECT 1927.930 1684.060 1928.250 1684.120 ;
        RECT 1931.150 1684.060 1931.470 1684.120 ;
      LAYER via ;
        RECT 1927.960 1684.060 1928.220 1684.320 ;
        RECT 1931.180 1684.060 1931.440 1684.320 ;
      LAYER met2 ;
        RECT 1927.950 1700.000 1928.230 1704.000 ;
        RECT 1928.020 1684.350 1928.160 1700.000 ;
        RECT 1927.960 1684.030 1928.220 1684.350 ;
        RECT 1931.180 1684.030 1931.440 1684.350 ;
        RECT 1931.240 24.325 1931.380 1684.030 ;
        RECT 1931.170 23.955 1931.450 24.325 ;
        RECT 2881.070 23.955 2881.350 24.325 ;
        RECT 2881.140 2.400 2881.280 23.955 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
      LAYER via2 ;
        RECT 1931.170 24.000 1931.450 24.280 ;
        RECT 2881.070 24.000 2881.350 24.280 ;
      LAYER met3 ;
        RECT 1931.145 24.290 1931.475 24.305 ;
        RECT 2881.045 24.290 2881.375 24.305 ;
        RECT 1931.145 23.990 2881.375 24.290 ;
        RECT 1931.145 23.975 1931.475 23.990 ;
        RECT 2881.045 23.975 2881.375 23.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1932.530 1685.620 1932.850 1685.680 ;
        RECT 1938.510 1685.620 1938.830 1685.680 ;
        RECT 1932.530 1685.480 1938.830 1685.620 ;
        RECT 1932.530 1685.420 1932.850 1685.480 ;
        RECT 1938.510 1685.420 1938.830 1685.480 ;
        RECT 1938.510 24.040 1938.830 24.100 ;
        RECT 2898.990 24.040 2899.310 24.100 ;
        RECT 1938.510 23.900 2899.310 24.040 ;
        RECT 1938.510 23.840 1938.830 23.900 ;
        RECT 2898.990 23.840 2899.310 23.900 ;
      LAYER via ;
        RECT 1932.560 1685.420 1932.820 1685.680 ;
        RECT 1938.540 1685.420 1938.800 1685.680 ;
        RECT 1938.540 23.840 1938.800 24.100 ;
        RECT 2899.020 23.840 2899.280 24.100 ;
      LAYER met2 ;
        RECT 1932.550 1700.000 1932.830 1704.000 ;
        RECT 1932.620 1685.710 1932.760 1700.000 ;
        RECT 1932.560 1685.390 1932.820 1685.710 ;
        RECT 1938.540 1685.390 1938.800 1685.710 ;
        RECT 1938.600 24.130 1938.740 1685.390 ;
        RECT 1938.540 23.810 1938.800 24.130 ;
        RECT 2899.020 23.810 2899.280 24.130 ;
        RECT 2899.080 2.400 2899.220 23.810 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 0.300 ;
=======
      LAYER met1 ;
        RECT 1373.170 1678.480 1373.490 1678.540 ;
        RECT 1377.310 1678.480 1377.630 1678.540 ;
        RECT 1373.170 1678.340 1377.630 1678.480 ;
        RECT 1373.170 1678.280 1373.490 1678.340 ;
        RECT 1377.310 1678.280 1377.630 1678.340 ;
      LAYER via ;
        RECT 1373.200 1678.280 1373.460 1678.540 ;
        RECT 1377.340 1678.280 1377.600 1678.540 ;
      LAYER met2 ;
        RECT 1378.250 1700.410 1378.530 1704.000 ;
        RECT 1377.400 1700.270 1378.530 1700.410 ;
        RECT 1377.400 1678.570 1377.540 1700.270 ;
        RECT 1378.250 1700.000 1378.530 1700.270 ;
        RECT 1373.200 1678.250 1373.460 1678.570 ;
        RECT 1377.340 1678.250 1377.600 1678.570 ;
        RECT 1373.260 26.365 1373.400 1678.250 ;
        RECT 846.950 25.995 847.230 26.365 ;
        RECT 1373.190 25.995 1373.470 26.365 ;
        RECT 847.020 2.400 847.160 25.995 ;
        RECT 846.810 -4.800 847.370 2.400 ;
      LAYER via2 ;
        RECT 846.950 26.040 847.230 26.320 ;
        RECT 1373.190 26.040 1373.470 26.320 ;
      LAYER met3 ;
        RECT 846.925 26.330 847.255 26.345 ;
        RECT 1373.165 26.330 1373.495 26.345 ;
        RECT 846.925 26.030 1373.495 26.330 ;
        RECT 846.925 26.015 847.255 26.030 ;
        RECT 1373.165 26.015 1373.495 26.030 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 864.750 -4.800 865.310 0.300 ;
=======
        RECT 1383.310 1700.410 1383.590 1704.000 ;
        RECT 1382.460 1700.270 1383.590 1700.410 ;
        RECT 1382.460 27.045 1382.600 1700.270 ;
        RECT 1383.310 1700.000 1383.590 1700.270 ;
        RECT 864.890 26.675 865.170 27.045 ;
        RECT 1382.390 26.675 1382.670 27.045 ;
        RECT 864.960 2.400 865.100 26.675 ;
        RECT 864.750 -4.800 865.310 2.400 ;
      LAYER via2 ;
        RECT 864.890 26.720 865.170 27.000 ;
        RECT 1382.390 26.720 1382.670 27.000 ;
      LAYER met3 ;
        RECT 864.865 27.010 865.195 27.025 ;
        RECT 1382.365 27.010 1382.695 27.025 ;
        RECT 864.865 26.710 1382.695 27.010 ;
        RECT 864.865 26.695 865.195 26.710 ;
        RECT 1382.365 26.695 1382.695 26.710 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 882.690 -4.800 883.250 0.300 ;
=======
        RECT 1387.910 1700.410 1388.190 1704.000 ;
        RECT 1387.060 1700.270 1388.190 1700.410 ;
        RECT 1387.060 27.725 1387.200 1700.270 ;
        RECT 1387.910 1700.000 1388.190 1700.270 ;
        RECT 882.830 27.355 883.110 27.725 ;
        RECT 1386.990 27.355 1387.270 27.725 ;
        RECT 882.900 2.400 883.040 27.355 ;
        RECT 882.690 -4.800 883.250 2.400 ;
      LAYER via2 ;
        RECT 882.830 27.400 883.110 27.680 ;
        RECT 1386.990 27.400 1387.270 27.680 ;
      LAYER met3 ;
        RECT 882.805 27.690 883.135 27.705 ;
        RECT 1386.965 27.690 1387.295 27.705 ;
        RECT 882.805 27.390 1387.295 27.690 ;
        RECT 882.805 27.375 883.135 27.390 ;
        RECT 1386.965 27.375 1387.295 27.390 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1387.430 1678.480 1387.750 1678.540 ;
        RECT 1391.570 1678.480 1391.890 1678.540 ;
        RECT 1387.430 1678.340 1391.890 1678.480 ;
        RECT 1387.430 1678.280 1387.750 1678.340 ;
        RECT 1391.570 1678.280 1391.890 1678.340 ;
        RECT 900.750 26.420 901.070 26.480 ;
        RECT 1387.430 26.420 1387.750 26.480 ;
        RECT 900.750 26.280 1387.750 26.420 ;
        RECT 900.750 26.220 901.070 26.280 ;
        RECT 1387.430 26.220 1387.750 26.280 ;
      LAYER via ;
        RECT 1387.460 1678.280 1387.720 1678.540 ;
        RECT 1391.600 1678.280 1391.860 1678.540 ;
        RECT 900.780 26.220 901.040 26.480 ;
        RECT 1387.460 26.220 1387.720 26.480 ;
      LAYER met2 ;
        RECT 1392.970 1700.410 1393.250 1704.000 ;
        RECT 1391.660 1700.270 1393.250 1700.410 ;
        RECT 1391.660 1678.570 1391.800 1700.270 ;
        RECT 1392.970 1700.000 1393.250 1700.270 ;
        RECT 1387.460 1678.250 1387.720 1678.570 ;
        RECT 1391.600 1678.250 1391.860 1678.570 ;
        RECT 1387.520 26.510 1387.660 1678.250 ;
        RECT 900.780 26.190 901.040 26.510 ;
        RECT 1387.460 26.190 1387.720 26.510 ;
        RECT 900.840 2.400 900.980 26.190 ;
        RECT 900.630 -4.800 901.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 0.300 ;
=======
      LAYER met1 ;
        RECT 1393.870 1678.480 1394.190 1678.540 ;
        RECT 1396.630 1678.480 1396.950 1678.540 ;
        RECT 1393.870 1678.340 1396.950 1678.480 ;
        RECT 1393.870 1678.280 1394.190 1678.340 ;
        RECT 1396.630 1678.280 1396.950 1678.340 ;
        RECT 918.690 26.760 919.010 26.820 ;
        RECT 1393.870 26.760 1394.190 26.820 ;
        RECT 918.690 26.620 1394.190 26.760 ;
        RECT 918.690 26.560 919.010 26.620 ;
        RECT 1393.870 26.560 1394.190 26.620 ;
      LAYER via ;
        RECT 1393.900 1678.280 1394.160 1678.540 ;
        RECT 1396.660 1678.280 1396.920 1678.540 ;
        RECT 918.720 26.560 918.980 26.820 ;
        RECT 1393.900 26.560 1394.160 26.820 ;
      LAYER met2 ;
        RECT 1397.570 1700.410 1397.850 1704.000 ;
        RECT 1396.720 1700.270 1397.850 1700.410 ;
        RECT 1396.720 1678.570 1396.860 1700.270 ;
        RECT 1397.570 1700.000 1397.850 1700.270 ;
        RECT 1393.900 1678.250 1394.160 1678.570 ;
        RECT 1396.660 1678.250 1396.920 1678.570 ;
        RECT 1393.960 26.850 1394.100 1678.250 ;
        RECT 918.720 26.530 918.980 26.850 ;
        RECT 1393.900 26.530 1394.160 26.850 ;
        RECT 918.780 2.400 918.920 26.530 ;
        RECT 918.570 -4.800 919.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 0.300 ;
=======
      LAYER met1 ;
        RECT 938.010 49.880 938.330 49.940 ;
        RECT 1402.610 49.880 1402.930 49.940 ;
        RECT 938.010 49.740 1402.930 49.880 ;
        RECT 938.010 49.680 938.330 49.740 ;
        RECT 1402.610 49.680 1402.930 49.740 ;
      LAYER via ;
        RECT 938.040 49.680 938.300 49.940 ;
        RECT 1402.640 49.680 1402.900 49.940 ;
      LAYER met2 ;
        RECT 1402.630 1700.000 1402.910 1704.000 ;
        RECT 1402.700 49.970 1402.840 1700.000 ;
        RECT 938.040 49.650 938.300 49.970 ;
        RECT 1402.640 49.650 1402.900 49.970 ;
        RECT 938.100 17.410 938.240 49.650 ;
        RECT 936.260 17.270 938.240 17.410 ;
        RECT 936.260 2.400 936.400 17.270 ;
        RECT 936.050 -4.800 936.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 0.300 ;
=======
      LAYER li1 ;
        RECT 1403.605 1490.645 1403.775 1568.675 ;
        RECT 1404.065 1248.905 1404.235 1297.015 ;
        RECT 1403.145 1048.985 1403.315 1097.095 ;
        RECT 1403.145 993.565 1403.315 1041.675 ;
        RECT 1403.605 234.685 1403.775 255.935 ;
      LAYER mcon ;
        RECT 1403.605 1568.505 1403.775 1568.675 ;
        RECT 1404.065 1296.845 1404.235 1297.015 ;
        RECT 1403.145 1096.925 1403.315 1097.095 ;
        RECT 1403.145 1041.505 1403.315 1041.675 ;
        RECT 1403.605 255.765 1403.775 255.935 ;
      LAYER met1 ;
        RECT 1403.530 1686.640 1403.850 1686.700 ;
        RECT 1407.210 1686.640 1407.530 1686.700 ;
        RECT 1403.530 1686.500 1407.530 1686.640 ;
        RECT 1403.530 1686.440 1403.850 1686.500 ;
        RECT 1407.210 1686.440 1407.530 1686.500 ;
        RECT 1403.070 1593.820 1403.390 1593.880 ;
        RECT 1403.530 1593.820 1403.850 1593.880 ;
        RECT 1403.070 1593.680 1403.850 1593.820 ;
        RECT 1403.070 1593.620 1403.390 1593.680 ;
        RECT 1403.530 1593.620 1403.850 1593.680 ;
        RECT 1403.070 1568.660 1403.390 1568.720 ;
        RECT 1403.545 1568.660 1403.835 1568.705 ;
        RECT 1403.070 1568.520 1403.835 1568.660 ;
        RECT 1403.070 1568.460 1403.390 1568.520 ;
        RECT 1403.545 1568.475 1403.835 1568.520 ;
        RECT 1403.530 1490.800 1403.850 1490.860 ;
        RECT 1403.335 1490.660 1403.850 1490.800 ;
        RECT 1403.530 1490.600 1403.850 1490.660 ;
        RECT 1403.530 1463.060 1403.850 1463.320 ;
        RECT 1403.620 1462.640 1403.760 1463.060 ;
        RECT 1403.530 1462.380 1403.850 1462.640 ;
        RECT 1403.530 1327.600 1403.850 1327.660 ;
        RECT 1403.990 1327.600 1404.310 1327.660 ;
        RECT 1403.530 1327.460 1404.310 1327.600 ;
        RECT 1403.530 1327.400 1403.850 1327.460 ;
        RECT 1403.990 1327.400 1404.310 1327.460 ;
        RECT 1403.990 1297.000 1404.310 1297.060 ;
        RECT 1403.795 1296.860 1404.310 1297.000 ;
        RECT 1403.990 1296.800 1404.310 1296.860 ;
        RECT 1404.005 1249.060 1404.295 1249.105 ;
        RECT 1404.450 1249.060 1404.770 1249.120 ;
        RECT 1404.005 1248.920 1404.770 1249.060 ;
        RECT 1404.005 1248.875 1404.295 1248.920 ;
        RECT 1404.450 1248.860 1404.770 1248.920 ;
        RECT 1403.530 1159.100 1403.850 1159.360 ;
        RECT 1403.620 1158.680 1403.760 1159.100 ;
        RECT 1403.530 1158.420 1403.850 1158.680 ;
        RECT 1403.530 1135.300 1403.850 1135.560 ;
        RECT 1403.620 1134.880 1403.760 1135.300 ;
        RECT 1403.530 1134.620 1403.850 1134.880 ;
        RECT 1403.085 1097.080 1403.375 1097.125 ;
        RECT 1403.530 1097.080 1403.850 1097.140 ;
        RECT 1403.085 1096.940 1403.850 1097.080 ;
        RECT 1403.085 1096.895 1403.375 1096.940 ;
        RECT 1403.530 1096.880 1403.850 1096.940 ;
        RECT 1403.070 1049.140 1403.390 1049.200 ;
        RECT 1402.875 1049.000 1403.390 1049.140 ;
        RECT 1403.070 1048.940 1403.390 1049.000 ;
        RECT 1403.070 1041.660 1403.390 1041.720 ;
        RECT 1402.875 1041.520 1403.390 1041.660 ;
        RECT 1403.070 1041.460 1403.390 1041.520 ;
        RECT 1403.085 993.720 1403.375 993.765 ;
        RECT 1403.530 993.720 1403.850 993.780 ;
        RECT 1403.085 993.580 1403.850 993.720 ;
        RECT 1403.085 993.535 1403.375 993.580 ;
        RECT 1403.530 993.520 1403.850 993.580 ;
        RECT 1403.530 966.520 1403.850 966.580 ;
        RECT 1403.160 966.380 1403.850 966.520 ;
        RECT 1403.160 965.900 1403.300 966.380 ;
        RECT 1403.530 966.320 1403.850 966.380 ;
        RECT 1403.070 965.640 1403.390 965.900 ;
        RECT 1403.070 917.900 1403.390 917.960 ;
        RECT 1403.530 917.900 1403.850 917.960 ;
        RECT 1403.070 917.760 1403.850 917.900 ;
        RECT 1403.070 917.700 1403.390 917.760 ;
        RECT 1403.530 917.700 1403.850 917.760 ;
        RECT 1403.070 724.440 1403.390 724.500 ;
        RECT 1403.990 724.440 1404.310 724.500 ;
        RECT 1403.070 724.300 1404.310 724.440 ;
        RECT 1403.070 724.240 1403.390 724.300 ;
        RECT 1403.990 724.240 1404.310 724.300 ;
        RECT 1403.070 579.600 1403.390 579.660 ;
        RECT 1403.990 579.600 1404.310 579.660 ;
        RECT 1403.070 579.460 1404.310 579.600 ;
        RECT 1403.070 579.400 1403.390 579.460 ;
        RECT 1403.990 579.400 1404.310 579.460 ;
        RECT 1403.530 255.920 1403.850 255.980 ;
        RECT 1403.335 255.780 1403.850 255.920 ;
        RECT 1403.530 255.720 1403.850 255.780 ;
        RECT 1403.530 234.840 1403.850 234.900 ;
        RECT 1403.335 234.700 1403.850 234.840 ;
        RECT 1403.530 234.640 1403.850 234.700 ;
        RECT 1403.530 137.740 1403.850 138.000 ;
        RECT 1403.620 137.320 1403.760 137.740 ;
        RECT 1403.530 137.060 1403.850 137.320 ;
        RECT 954.110 27.100 954.430 27.160 ;
        RECT 1402.610 27.100 1402.930 27.160 ;
        RECT 954.110 26.960 1402.930 27.100 ;
        RECT 954.110 26.900 954.430 26.960 ;
        RECT 1402.610 26.900 1402.930 26.960 ;
      LAYER via ;
        RECT 1403.560 1686.440 1403.820 1686.700 ;
        RECT 1407.240 1686.440 1407.500 1686.700 ;
        RECT 1403.100 1593.620 1403.360 1593.880 ;
        RECT 1403.560 1593.620 1403.820 1593.880 ;
        RECT 1403.100 1568.460 1403.360 1568.720 ;
        RECT 1403.560 1490.600 1403.820 1490.860 ;
        RECT 1403.560 1463.060 1403.820 1463.320 ;
        RECT 1403.560 1462.380 1403.820 1462.640 ;
        RECT 1403.560 1327.400 1403.820 1327.660 ;
        RECT 1404.020 1327.400 1404.280 1327.660 ;
        RECT 1404.020 1296.800 1404.280 1297.060 ;
        RECT 1404.480 1248.860 1404.740 1249.120 ;
        RECT 1403.560 1159.100 1403.820 1159.360 ;
        RECT 1403.560 1158.420 1403.820 1158.680 ;
        RECT 1403.560 1135.300 1403.820 1135.560 ;
        RECT 1403.560 1134.620 1403.820 1134.880 ;
        RECT 1403.560 1096.880 1403.820 1097.140 ;
        RECT 1403.100 1048.940 1403.360 1049.200 ;
        RECT 1403.100 1041.460 1403.360 1041.720 ;
        RECT 1403.560 993.520 1403.820 993.780 ;
        RECT 1403.560 966.320 1403.820 966.580 ;
        RECT 1403.100 965.640 1403.360 965.900 ;
        RECT 1403.100 917.700 1403.360 917.960 ;
        RECT 1403.560 917.700 1403.820 917.960 ;
        RECT 1403.100 724.240 1403.360 724.500 ;
        RECT 1404.020 724.240 1404.280 724.500 ;
        RECT 1403.100 579.400 1403.360 579.660 ;
        RECT 1404.020 579.400 1404.280 579.660 ;
        RECT 1403.560 255.720 1403.820 255.980 ;
        RECT 1403.560 234.640 1403.820 234.900 ;
        RECT 1403.560 137.740 1403.820 138.000 ;
        RECT 1403.560 137.060 1403.820 137.320 ;
        RECT 954.140 26.900 954.400 27.160 ;
        RECT 1402.640 26.900 1402.900 27.160 ;
      LAYER met2 ;
        RECT 1407.230 1700.000 1407.510 1704.000 ;
        RECT 1407.300 1686.730 1407.440 1700.000 ;
        RECT 1403.560 1686.410 1403.820 1686.730 ;
        RECT 1407.240 1686.410 1407.500 1686.730 ;
        RECT 1403.620 1593.910 1403.760 1686.410 ;
        RECT 1403.100 1593.590 1403.360 1593.910 ;
        RECT 1403.560 1593.590 1403.820 1593.910 ;
        RECT 1403.160 1568.750 1403.300 1593.590 ;
        RECT 1403.100 1568.430 1403.360 1568.750 ;
        RECT 1403.560 1490.570 1403.820 1490.890 ;
        RECT 1403.620 1463.350 1403.760 1490.570 ;
        RECT 1403.560 1463.030 1403.820 1463.350 ;
        RECT 1403.560 1462.350 1403.820 1462.670 ;
        RECT 1403.620 1327.690 1403.760 1462.350 ;
        RECT 1403.560 1327.370 1403.820 1327.690 ;
        RECT 1404.020 1327.370 1404.280 1327.690 ;
        RECT 1404.080 1297.090 1404.220 1327.370 ;
        RECT 1404.020 1296.770 1404.280 1297.090 ;
        RECT 1404.480 1248.830 1404.740 1249.150 ;
        RECT 1404.540 1208.090 1404.680 1248.830 ;
        RECT 1404.080 1207.950 1404.680 1208.090 ;
        RECT 1404.080 1200.610 1404.220 1207.950 ;
        RECT 1403.620 1200.470 1404.220 1200.610 ;
        RECT 1403.620 1159.390 1403.760 1200.470 ;
        RECT 1403.560 1159.070 1403.820 1159.390 ;
        RECT 1403.560 1158.390 1403.820 1158.710 ;
        RECT 1403.620 1135.590 1403.760 1158.390 ;
        RECT 1403.560 1135.270 1403.820 1135.590 ;
        RECT 1403.560 1134.590 1403.820 1134.910 ;
        RECT 1403.620 1097.170 1403.760 1134.590 ;
        RECT 1403.560 1096.850 1403.820 1097.170 ;
        RECT 1403.100 1048.910 1403.360 1049.230 ;
        RECT 1403.160 1041.750 1403.300 1048.910 ;
        RECT 1403.100 1041.430 1403.360 1041.750 ;
        RECT 1403.560 993.490 1403.820 993.810 ;
        RECT 1403.620 966.610 1403.760 993.490 ;
        RECT 1403.560 966.290 1403.820 966.610 ;
        RECT 1403.100 965.610 1403.360 965.930 ;
        RECT 1403.160 917.990 1403.300 965.610 ;
        RECT 1403.100 917.670 1403.360 917.990 ;
        RECT 1403.560 917.670 1403.820 917.990 ;
        RECT 1403.620 835.450 1403.760 917.670 ;
        RECT 1403.160 835.310 1403.760 835.450 ;
        RECT 1403.160 834.770 1403.300 835.310 ;
        RECT 1403.160 834.630 1403.760 834.770 ;
        RECT 1403.620 738.890 1403.760 834.630 ;
        RECT 1403.620 738.750 1404.220 738.890 ;
        RECT 1404.080 724.725 1404.220 738.750 ;
        RECT 1403.090 724.355 1403.370 724.725 ;
        RECT 1404.010 724.355 1404.290 724.725 ;
        RECT 1403.100 724.210 1403.360 724.355 ;
        RECT 1404.020 724.210 1404.280 724.355 ;
        RECT 1404.080 688.570 1404.220 724.210 ;
        RECT 1403.620 688.430 1404.220 688.570 ;
        RECT 1403.620 580.565 1403.760 688.430 ;
        RECT 1403.550 580.195 1403.830 580.565 ;
        RECT 1403.090 579.515 1403.370 579.885 ;
        RECT 1403.100 579.370 1403.360 579.515 ;
        RECT 1404.020 579.370 1404.280 579.690 ;
        RECT 1404.080 531.490 1404.220 579.370 ;
        RECT 1403.620 531.350 1404.220 531.490 ;
        RECT 1403.620 256.010 1403.760 531.350 ;
        RECT 1403.560 255.690 1403.820 256.010 ;
        RECT 1403.560 234.610 1403.820 234.930 ;
        RECT 1403.620 211.210 1403.760 234.610 ;
        RECT 1403.620 211.070 1404.220 211.210 ;
        RECT 1404.080 138.450 1404.220 211.070 ;
        RECT 1403.620 138.310 1404.220 138.450 ;
        RECT 1403.620 138.030 1403.760 138.310 ;
        RECT 1403.560 137.710 1403.820 138.030 ;
        RECT 1403.560 137.030 1403.820 137.350 ;
        RECT 1403.620 49.370 1403.760 137.030 ;
        RECT 1402.700 49.230 1403.760 49.370 ;
        RECT 1402.700 27.190 1402.840 49.230 ;
        RECT 954.140 26.870 954.400 27.190 ;
        RECT 1402.640 26.870 1402.900 27.190 ;
        RECT 954.200 2.400 954.340 26.870 ;
        RECT 953.990 -4.800 954.550 2.400 ;
      LAYER via2 ;
        RECT 1403.090 724.400 1403.370 724.680 ;
        RECT 1404.010 724.400 1404.290 724.680 ;
        RECT 1403.550 580.240 1403.830 580.520 ;
        RECT 1403.090 579.560 1403.370 579.840 ;
      LAYER met3 ;
        RECT 1403.065 724.690 1403.395 724.705 ;
        RECT 1403.985 724.690 1404.315 724.705 ;
        RECT 1403.065 724.390 1404.315 724.690 ;
        RECT 1403.065 724.375 1403.395 724.390 ;
        RECT 1403.985 724.375 1404.315 724.390 ;
        RECT 1403.525 580.530 1403.855 580.545 ;
        RECT 1402.390 580.230 1403.855 580.530 ;
        RECT 1402.390 579.850 1402.690 580.230 ;
        RECT 1403.525 580.215 1403.855 580.230 ;
        RECT 1403.065 579.850 1403.395 579.865 ;
        RECT 1402.390 579.550 1403.395 579.850 ;
        RECT 1403.065 579.535 1403.395 579.550 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1407.670 1678.480 1407.990 1678.540 ;
        RECT 1410.890 1678.480 1411.210 1678.540 ;
        RECT 1407.670 1678.340 1411.210 1678.480 ;
        RECT 1407.670 1678.280 1407.990 1678.340 ;
        RECT 1410.890 1678.280 1411.210 1678.340 ;
        RECT 972.050 27.440 972.370 27.500 ;
        RECT 1407.670 27.440 1407.990 27.500 ;
        RECT 972.050 27.300 1407.990 27.440 ;
        RECT 972.050 27.240 972.370 27.300 ;
        RECT 1407.670 27.240 1407.990 27.300 ;
      LAYER via ;
        RECT 1407.700 1678.280 1407.960 1678.540 ;
        RECT 1410.920 1678.280 1411.180 1678.540 ;
        RECT 972.080 27.240 972.340 27.500 ;
        RECT 1407.700 27.240 1407.960 27.500 ;
      LAYER met2 ;
        RECT 1412.290 1700.410 1412.570 1704.000 ;
        RECT 1410.980 1700.270 1412.570 1700.410 ;
        RECT 1410.980 1678.570 1411.120 1700.270 ;
        RECT 1412.290 1700.000 1412.570 1700.270 ;
        RECT 1407.700 1678.250 1407.960 1678.570 ;
        RECT 1410.920 1678.250 1411.180 1678.570 ;
        RECT 1407.760 27.530 1407.900 1678.250 ;
        RECT 972.080 27.210 972.340 27.530 ;
        RECT 1407.700 27.210 1407.960 27.530 ;
        RECT 972.140 2.400 972.280 27.210 ;
        RECT 971.930 -4.800 972.490 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 650.850 -4.800 651.410 0.300 ;
=======
        RECT 1325.350 1700.410 1325.630 1704.000 ;
        RECT 1324.960 1700.270 1325.630 1700.410 ;
        RECT 1324.960 25.685 1325.100 1700.270 ;
        RECT 1325.350 1700.000 1325.630 1700.270 ;
        RECT 650.990 25.315 651.270 25.685 ;
        RECT 1324.890 25.315 1325.170 25.685 ;
        RECT 651.060 2.400 651.200 25.315 ;
        RECT 650.850 -4.800 651.410 2.400 ;
      LAYER via2 ;
        RECT 650.990 25.360 651.270 25.640 ;
        RECT 1324.890 25.360 1325.170 25.640 ;
      LAYER met3 ;
        RECT 650.965 25.650 651.295 25.665 ;
        RECT 1324.865 25.650 1325.195 25.665 ;
        RECT 650.965 25.350 1325.195 25.650 ;
        RECT 650.965 25.335 651.295 25.350 ;
        RECT 1324.865 25.335 1325.195 25.350 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1414.570 1678.140 1414.890 1678.200 ;
        RECT 1415.950 1678.140 1416.270 1678.200 ;
        RECT 1414.570 1678.000 1416.270 1678.140 ;
        RECT 1414.570 1677.940 1414.890 1678.000 ;
        RECT 1415.950 1677.940 1416.270 1678.000 ;
        RECT 989.990 23.700 990.310 23.760 ;
        RECT 1414.570 23.700 1414.890 23.760 ;
        RECT 989.990 23.560 1414.890 23.700 ;
        RECT 989.990 23.500 990.310 23.560 ;
        RECT 1414.570 23.500 1414.890 23.560 ;
      LAYER via ;
        RECT 1414.600 1677.940 1414.860 1678.200 ;
        RECT 1415.980 1677.940 1416.240 1678.200 ;
        RECT 990.020 23.500 990.280 23.760 ;
        RECT 1414.600 23.500 1414.860 23.760 ;
      LAYER met2 ;
        RECT 1416.890 1700.410 1417.170 1704.000 ;
        RECT 1416.040 1700.270 1417.170 1700.410 ;
        RECT 1416.040 1678.230 1416.180 1700.270 ;
        RECT 1416.890 1700.000 1417.170 1700.270 ;
        RECT 1414.600 1677.910 1414.860 1678.230 ;
        RECT 1415.980 1677.910 1416.240 1678.230 ;
        RECT 1414.660 23.790 1414.800 1677.910 ;
        RECT 990.020 23.470 990.280 23.790 ;
        RECT 1414.600 23.470 1414.860 23.790 ;
        RECT 990.080 2.400 990.220 23.470 ;
        RECT 989.870 -4.800 990.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1007.470 23.360 1007.790 23.420 ;
        RECT 1421.930 23.360 1422.250 23.420 ;
        RECT 1007.470 23.220 1422.250 23.360 ;
        RECT 1007.470 23.160 1007.790 23.220 ;
        RECT 1421.930 23.160 1422.250 23.220 ;
      LAYER via ;
        RECT 1007.500 23.160 1007.760 23.420 ;
        RECT 1421.960 23.160 1422.220 23.420 ;
      LAYER met2 ;
        RECT 1421.950 1700.000 1422.230 1704.000 ;
        RECT 1422.020 23.450 1422.160 1700.000 ;
        RECT 1007.500 23.130 1007.760 23.450 ;
        RECT 1421.960 23.130 1422.220 23.450 ;
        RECT 1007.560 2.400 1007.700 23.130 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1421.470 1678.140 1421.790 1678.200 ;
        RECT 1425.610 1678.140 1425.930 1678.200 ;
        RECT 1421.470 1678.000 1425.930 1678.140 ;
        RECT 1421.470 1677.940 1421.790 1678.000 ;
        RECT 1425.610 1677.940 1425.930 1678.000 ;
        RECT 1025.410 23.020 1025.730 23.080 ;
        RECT 1421.470 23.020 1421.790 23.080 ;
        RECT 1025.410 22.880 1421.790 23.020 ;
        RECT 1025.410 22.820 1025.730 22.880 ;
        RECT 1421.470 22.820 1421.790 22.880 ;
      LAYER via ;
        RECT 1421.500 1677.940 1421.760 1678.200 ;
        RECT 1425.640 1677.940 1425.900 1678.200 ;
        RECT 1025.440 22.820 1025.700 23.080 ;
        RECT 1421.500 22.820 1421.760 23.080 ;
      LAYER met2 ;
        RECT 1426.550 1700.410 1426.830 1704.000 ;
        RECT 1425.700 1700.270 1426.830 1700.410 ;
        RECT 1425.700 1678.230 1425.840 1700.270 ;
        RECT 1426.550 1700.000 1426.830 1700.270 ;
        RECT 1421.500 1677.910 1421.760 1678.230 ;
        RECT 1425.640 1677.910 1425.900 1678.230 ;
        RECT 1421.560 23.110 1421.700 1677.910 ;
        RECT 1025.440 22.790 1025.700 23.110 ;
        RECT 1421.500 22.790 1421.760 23.110 ;
        RECT 1025.500 2.400 1025.640 22.790 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 0.300 ;
=======
      LAYER met1 ;
        RECT 1043.350 22.680 1043.670 22.740 ;
        RECT 1430.670 22.680 1430.990 22.740 ;
        RECT 1043.350 22.540 1430.990 22.680 ;
        RECT 1043.350 22.480 1043.670 22.540 ;
        RECT 1430.670 22.480 1430.990 22.540 ;
      LAYER via ;
        RECT 1043.380 22.480 1043.640 22.740 ;
        RECT 1430.700 22.480 1430.960 22.740 ;
      LAYER met2 ;
        RECT 1431.610 1700.410 1431.890 1704.000 ;
        RECT 1430.760 1700.270 1431.890 1700.410 ;
        RECT 1430.760 22.770 1430.900 1700.270 ;
        RECT 1431.610 1700.000 1431.890 1700.270 ;
        RECT 1043.380 22.450 1043.640 22.770 ;
        RECT 1430.700 22.450 1430.960 22.770 ;
        RECT 1043.440 2.400 1043.580 22.450 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1061.290 22.340 1061.610 22.400 ;
        RECT 1435.270 22.340 1435.590 22.400 ;
        RECT 1061.290 22.200 1435.590 22.340 ;
        RECT 1061.290 22.140 1061.610 22.200 ;
        RECT 1435.270 22.140 1435.590 22.200 ;
      LAYER via ;
        RECT 1061.320 22.140 1061.580 22.400 ;
        RECT 1435.300 22.140 1435.560 22.400 ;
      LAYER met2 ;
        RECT 1436.210 1700.410 1436.490 1704.000 ;
        RECT 1435.360 1700.270 1436.490 1700.410 ;
        RECT 1435.360 22.430 1435.500 1700.270 ;
        RECT 1436.210 1700.000 1436.490 1700.270 ;
        RECT 1061.320 22.110 1061.580 22.430 ;
        RECT 1435.300 22.110 1435.560 22.430 ;
        RECT 1061.380 2.400 1061.520 22.110 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1435.730 1678.140 1436.050 1678.200 ;
        RECT 1439.870 1678.140 1440.190 1678.200 ;
        RECT 1435.730 1678.000 1440.190 1678.140 ;
        RECT 1435.730 1677.940 1436.050 1678.000 ;
        RECT 1439.870 1677.940 1440.190 1678.000 ;
        RECT 1079.230 22.000 1079.550 22.060 ;
        RECT 1435.730 22.000 1436.050 22.060 ;
        RECT 1079.230 21.860 1436.050 22.000 ;
        RECT 1079.230 21.800 1079.550 21.860 ;
        RECT 1435.730 21.800 1436.050 21.860 ;
      LAYER via ;
        RECT 1435.760 1677.940 1436.020 1678.200 ;
        RECT 1439.900 1677.940 1440.160 1678.200 ;
        RECT 1079.260 21.800 1079.520 22.060 ;
        RECT 1435.760 21.800 1436.020 22.060 ;
      LAYER met2 ;
        RECT 1441.270 1700.410 1441.550 1704.000 ;
        RECT 1439.960 1700.270 1441.550 1700.410 ;
        RECT 1439.960 1678.230 1440.100 1700.270 ;
        RECT 1441.270 1700.000 1441.550 1700.270 ;
        RECT 1435.760 1677.910 1436.020 1678.230 ;
        RECT 1439.900 1677.910 1440.160 1678.230 ;
        RECT 1435.820 22.090 1435.960 1677.910 ;
        RECT 1079.260 21.770 1079.520 22.090 ;
        RECT 1435.760 21.770 1436.020 22.090 ;
        RECT 1079.320 2.400 1079.460 21.770 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 0.300 ;
=======
      LAYER met1 ;
        RECT 1442.170 1678.140 1442.490 1678.200 ;
        RECT 1444.930 1678.140 1445.250 1678.200 ;
        RECT 1442.170 1678.000 1445.250 1678.140 ;
        RECT 1442.170 1677.940 1442.490 1678.000 ;
        RECT 1444.930 1677.940 1445.250 1678.000 ;
        RECT 1096.710 21.660 1097.030 21.720 ;
        RECT 1442.170 21.660 1442.490 21.720 ;
        RECT 1096.710 21.520 1442.490 21.660 ;
        RECT 1096.710 21.460 1097.030 21.520 ;
        RECT 1442.170 21.460 1442.490 21.520 ;
      LAYER via ;
        RECT 1442.200 1677.940 1442.460 1678.200 ;
        RECT 1444.960 1677.940 1445.220 1678.200 ;
        RECT 1096.740 21.460 1097.000 21.720 ;
        RECT 1442.200 21.460 1442.460 21.720 ;
      LAYER met2 ;
        RECT 1445.870 1700.410 1446.150 1704.000 ;
        RECT 1445.020 1700.270 1446.150 1700.410 ;
        RECT 1445.020 1678.230 1445.160 1700.270 ;
        RECT 1445.870 1700.000 1446.150 1700.270 ;
        RECT 1442.200 1677.910 1442.460 1678.230 ;
        RECT 1444.960 1677.910 1445.220 1678.230 ;
        RECT 1442.260 21.750 1442.400 1677.910 ;
        RECT 1096.740 21.430 1097.000 21.750 ;
        RECT 1442.200 21.430 1442.460 21.750 ;
        RECT 1096.800 2.400 1096.940 21.430 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1449.530 1658.420 1449.850 1658.480 ;
        RECT 1450.450 1658.420 1450.770 1658.480 ;
        RECT 1449.530 1658.280 1450.770 1658.420 ;
        RECT 1449.530 1658.220 1449.850 1658.280 ;
        RECT 1450.450 1658.220 1450.770 1658.280 ;
        RECT 1449.530 290.060 1449.850 290.320 ;
        RECT 1449.620 289.640 1449.760 290.060 ;
        RECT 1449.530 289.380 1449.850 289.640 ;
        RECT 1114.650 21.320 1114.970 21.380 ;
        RECT 1449.530 21.320 1449.850 21.380 ;
        RECT 1114.650 21.180 1449.850 21.320 ;
        RECT 1114.650 21.120 1114.970 21.180 ;
        RECT 1449.530 21.120 1449.850 21.180 ;
      LAYER via ;
        RECT 1449.560 1658.220 1449.820 1658.480 ;
        RECT 1450.480 1658.220 1450.740 1658.480 ;
        RECT 1449.560 290.060 1449.820 290.320 ;
        RECT 1449.560 289.380 1449.820 289.640 ;
        RECT 1114.680 21.120 1114.940 21.380 ;
        RECT 1449.560 21.120 1449.820 21.380 ;
      LAYER met2 ;
        RECT 1450.470 1700.000 1450.750 1704.000 ;
        RECT 1450.540 1658.510 1450.680 1700.000 ;
        RECT 1449.560 1658.190 1449.820 1658.510 ;
        RECT 1450.480 1658.190 1450.740 1658.510 ;
        RECT 1449.620 290.350 1449.760 1658.190 ;
        RECT 1449.560 290.030 1449.820 290.350 ;
        RECT 1449.560 289.350 1449.820 289.670 ;
        RECT 1449.620 21.410 1449.760 289.350 ;
        RECT 1114.680 21.090 1114.940 21.410 ;
        RECT 1449.560 21.090 1449.820 21.410 ;
        RECT 1114.740 2.400 1114.880 21.090 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 0.300 ;
=======
      LAYER li1 ;
        RECT 1451.445 964.665 1451.615 966.535 ;
      LAYER mcon ;
        RECT 1451.445 966.365 1451.615 966.535 ;
      LAYER met1 ;
        RECT 1451.370 1678.140 1451.690 1678.200 ;
        RECT 1454.130 1678.140 1454.450 1678.200 ;
        RECT 1451.370 1678.000 1454.450 1678.140 ;
        RECT 1451.370 1677.940 1451.690 1678.000 ;
        RECT 1454.130 1677.940 1454.450 1678.000 ;
        RECT 1451.370 1153.320 1451.690 1153.580 ;
        RECT 1451.460 1152.560 1451.600 1153.320 ;
        RECT 1451.370 1152.300 1451.690 1152.560 ;
        RECT 1451.370 966.520 1451.690 966.580 ;
        RECT 1451.175 966.380 1451.690 966.520 ;
        RECT 1451.370 966.320 1451.690 966.380 ;
        RECT 1451.370 964.820 1451.690 964.880 ;
        RECT 1451.175 964.680 1451.690 964.820 ;
        RECT 1451.370 964.620 1451.690 964.680 ;
        RECT 1132.590 20.980 1132.910 21.040 ;
        RECT 1451.370 20.980 1451.690 21.040 ;
        RECT 1132.590 20.840 1451.690 20.980 ;
        RECT 1132.590 20.780 1132.910 20.840 ;
        RECT 1451.370 20.780 1451.690 20.840 ;
      LAYER via ;
        RECT 1451.400 1677.940 1451.660 1678.200 ;
        RECT 1454.160 1677.940 1454.420 1678.200 ;
        RECT 1451.400 1153.320 1451.660 1153.580 ;
        RECT 1451.400 1152.300 1451.660 1152.560 ;
        RECT 1451.400 966.320 1451.660 966.580 ;
        RECT 1451.400 964.620 1451.660 964.880 ;
        RECT 1132.620 20.780 1132.880 21.040 ;
        RECT 1451.400 20.780 1451.660 21.040 ;
      LAYER met2 ;
        RECT 1455.530 1700.410 1455.810 1704.000 ;
        RECT 1454.220 1700.270 1455.810 1700.410 ;
        RECT 1454.220 1678.230 1454.360 1700.270 ;
        RECT 1455.530 1700.000 1455.810 1700.270 ;
        RECT 1451.400 1677.910 1451.660 1678.230 ;
        RECT 1454.160 1677.910 1454.420 1678.230 ;
        RECT 1451.460 1153.610 1451.600 1677.910 ;
        RECT 1451.400 1153.290 1451.660 1153.610 ;
        RECT 1451.400 1152.270 1451.660 1152.590 ;
        RECT 1451.460 966.610 1451.600 1152.270 ;
        RECT 1451.400 966.290 1451.660 966.610 ;
        RECT 1451.400 964.590 1451.660 964.910 ;
        RECT 1451.460 21.070 1451.600 964.590 ;
        RECT 1132.620 20.750 1132.880 21.070 ;
        RECT 1451.400 20.750 1451.660 21.070 ;
        RECT 1132.680 2.400 1132.820 20.750 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 0.300 ;
=======
      LAYER met1 ;
        RECT 1456.430 1678.140 1456.750 1678.200 ;
        RECT 1459.190 1678.140 1459.510 1678.200 ;
        RECT 1456.430 1678.000 1459.510 1678.140 ;
        RECT 1456.430 1677.940 1456.750 1678.000 ;
        RECT 1459.190 1677.940 1459.510 1678.000 ;
        RECT 1150.530 24.040 1150.850 24.100 ;
        RECT 1456.430 24.040 1456.750 24.100 ;
        RECT 1150.530 23.900 1456.750 24.040 ;
        RECT 1150.530 23.840 1150.850 23.900 ;
        RECT 1456.430 23.840 1456.750 23.900 ;
      LAYER via ;
        RECT 1456.460 1677.940 1456.720 1678.200 ;
        RECT 1459.220 1677.940 1459.480 1678.200 ;
        RECT 1150.560 23.840 1150.820 24.100 ;
        RECT 1456.460 23.840 1456.720 24.100 ;
      LAYER met2 ;
        RECT 1460.130 1700.410 1460.410 1704.000 ;
        RECT 1459.280 1700.270 1460.410 1700.410 ;
        RECT 1459.280 1678.230 1459.420 1700.270 ;
        RECT 1460.130 1700.000 1460.410 1700.270 ;
        RECT 1456.460 1677.910 1456.720 1678.230 ;
        RECT 1459.220 1677.910 1459.480 1678.230 ;
        RECT 1456.520 24.130 1456.660 1677.910 ;
        RECT 1150.560 23.810 1150.820 24.130 ;
        RECT 1456.460 23.810 1456.720 24.130 ;
        RECT 1150.620 2.400 1150.760 23.810 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 0.300 ;
=======
      LAYER li1 ;
        RECT 1326.785 1345.125 1326.955 1368.075 ;
        RECT 1326.785 642.345 1326.955 710.515 ;
        RECT 1327.245 559.045 1327.415 607.155 ;
        RECT 1327.705 475.745 1327.875 537.115 ;
      LAYER mcon ;
        RECT 1326.785 1367.905 1326.955 1368.075 ;
        RECT 1326.785 710.345 1326.955 710.515 ;
        RECT 1327.245 606.985 1327.415 607.155 ;
        RECT 1327.705 536.945 1327.875 537.115 ;
      LAYER met1 ;
        RECT 1326.710 1642.440 1327.030 1642.500 ;
        RECT 1329.470 1642.440 1329.790 1642.500 ;
        RECT 1326.710 1642.300 1329.790 1642.440 ;
        RECT 1326.710 1642.240 1327.030 1642.300 ;
        RECT 1329.470 1642.240 1329.790 1642.300 ;
        RECT 1326.710 1545.880 1327.030 1545.940 ;
        RECT 1327.170 1545.880 1327.490 1545.940 ;
        RECT 1326.710 1545.740 1327.490 1545.880 ;
        RECT 1326.710 1545.680 1327.030 1545.740 ;
        RECT 1327.170 1545.680 1327.490 1545.740 ;
        RECT 1327.630 1401.380 1327.950 1401.440 ;
        RECT 1326.800 1401.240 1327.950 1401.380 ;
        RECT 1326.800 1401.100 1326.940 1401.240 ;
        RECT 1327.630 1401.180 1327.950 1401.240 ;
        RECT 1326.710 1400.840 1327.030 1401.100 ;
        RECT 1326.710 1368.060 1327.030 1368.120 ;
        RECT 1326.515 1367.920 1327.030 1368.060 ;
        RECT 1326.710 1367.860 1327.030 1367.920 ;
        RECT 1326.725 1345.280 1327.015 1345.325 ;
        RECT 1327.630 1345.280 1327.950 1345.340 ;
        RECT 1326.725 1345.140 1327.950 1345.280 ;
        RECT 1326.725 1345.095 1327.015 1345.140 ;
        RECT 1327.630 1345.080 1327.950 1345.140 ;
        RECT 1327.170 1297.340 1327.490 1297.400 ;
        RECT 1327.630 1297.340 1327.950 1297.400 ;
        RECT 1327.170 1297.200 1327.950 1297.340 ;
        RECT 1327.170 1297.140 1327.490 1297.200 ;
        RECT 1327.630 1297.140 1327.950 1297.200 ;
        RECT 1326.710 1249.060 1327.030 1249.120 ;
        RECT 1327.170 1249.060 1327.490 1249.120 ;
        RECT 1326.710 1248.920 1327.490 1249.060 ;
        RECT 1326.710 1248.860 1327.030 1248.920 ;
        RECT 1327.170 1248.860 1327.490 1248.920 ;
        RECT 1327.170 814.540 1327.490 814.600 ;
        RECT 1326.800 814.400 1327.490 814.540 ;
        RECT 1326.800 814.260 1326.940 814.400 ;
        RECT 1327.170 814.340 1327.490 814.400 ;
        RECT 1326.710 814.000 1327.030 814.260 ;
        RECT 1326.710 710.500 1327.030 710.560 ;
        RECT 1326.515 710.360 1327.030 710.500 ;
        RECT 1326.710 710.300 1327.030 710.360 ;
        RECT 1326.725 642.500 1327.015 642.545 ;
        RECT 1327.170 642.500 1327.490 642.560 ;
        RECT 1326.725 642.360 1327.490 642.500 ;
        RECT 1326.725 642.315 1327.015 642.360 ;
        RECT 1327.170 642.300 1327.490 642.360 ;
        RECT 1327.170 607.140 1327.490 607.200 ;
        RECT 1326.975 607.000 1327.490 607.140 ;
        RECT 1327.170 606.940 1327.490 607.000 ;
        RECT 1326.710 559.200 1327.030 559.260 ;
        RECT 1327.185 559.200 1327.475 559.245 ;
        RECT 1326.710 559.060 1327.475 559.200 ;
        RECT 1326.710 559.000 1327.030 559.060 ;
        RECT 1327.185 559.015 1327.475 559.060 ;
        RECT 1326.710 537.100 1327.030 537.160 ;
        RECT 1327.645 537.100 1327.935 537.145 ;
        RECT 1326.710 536.960 1327.935 537.100 ;
        RECT 1326.710 536.900 1327.030 536.960 ;
        RECT 1327.645 536.915 1327.935 536.960 ;
        RECT 1327.630 475.900 1327.950 475.960 ;
        RECT 1327.435 475.760 1327.950 475.900 ;
        RECT 1327.630 475.700 1327.950 475.760 ;
        RECT 1327.170 427.960 1327.490 428.020 ;
        RECT 1327.630 427.960 1327.950 428.020 ;
        RECT 1327.170 427.820 1327.950 427.960 ;
        RECT 1327.170 427.760 1327.490 427.820 ;
        RECT 1327.630 427.760 1327.950 427.820 ;
        RECT 1326.710 379.680 1327.030 379.740 ;
        RECT 1327.170 379.680 1327.490 379.740 ;
        RECT 1326.710 379.540 1327.490 379.680 ;
        RECT 1326.710 379.480 1327.030 379.540 ;
        RECT 1327.170 379.480 1327.490 379.540 ;
        RECT 1326.710 331.060 1327.030 331.120 ;
        RECT 1327.170 331.060 1327.490 331.120 ;
        RECT 1326.710 330.920 1327.490 331.060 ;
        RECT 1326.710 330.860 1327.030 330.920 ;
        RECT 1327.170 330.860 1327.490 330.920 ;
        RECT 1327.170 186.900 1327.490 186.960 ;
        RECT 1326.800 186.760 1327.490 186.900 ;
        RECT 1326.800 186.620 1326.940 186.760 ;
        RECT 1327.170 186.700 1327.490 186.760 ;
        RECT 1326.710 186.360 1327.030 186.620 ;
        RECT 1326.710 110.540 1327.030 110.800 ;
        RECT 1326.800 110.060 1326.940 110.540 ;
        RECT 1327.170 110.060 1327.490 110.120 ;
        RECT 1326.800 109.920 1327.490 110.060 ;
        RECT 1327.170 109.860 1327.490 109.920 ;
        RECT 668.910 25.740 669.230 25.800 ;
        RECT 1326.710 25.740 1327.030 25.800 ;
        RECT 668.910 25.600 1327.030 25.740 ;
        RECT 668.910 25.540 669.230 25.600 ;
        RECT 1326.710 25.540 1327.030 25.600 ;
      LAYER via ;
        RECT 1326.740 1642.240 1327.000 1642.500 ;
        RECT 1329.500 1642.240 1329.760 1642.500 ;
        RECT 1326.740 1545.680 1327.000 1545.940 ;
        RECT 1327.200 1545.680 1327.460 1545.940 ;
        RECT 1327.660 1401.180 1327.920 1401.440 ;
        RECT 1326.740 1400.840 1327.000 1401.100 ;
        RECT 1326.740 1367.860 1327.000 1368.120 ;
        RECT 1327.660 1345.080 1327.920 1345.340 ;
        RECT 1327.200 1297.140 1327.460 1297.400 ;
        RECT 1327.660 1297.140 1327.920 1297.400 ;
        RECT 1326.740 1248.860 1327.000 1249.120 ;
        RECT 1327.200 1248.860 1327.460 1249.120 ;
        RECT 1327.200 814.340 1327.460 814.600 ;
        RECT 1326.740 814.000 1327.000 814.260 ;
        RECT 1326.740 710.300 1327.000 710.560 ;
        RECT 1327.200 642.300 1327.460 642.560 ;
        RECT 1327.200 606.940 1327.460 607.200 ;
        RECT 1326.740 559.000 1327.000 559.260 ;
        RECT 1326.740 536.900 1327.000 537.160 ;
        RECT 1327.660 475.700 1327.920 475.960 ;
        RECT 1327.200 427.760 1327.460 428.020 ;
        RECT 1327.660 427.760 1327.920 428.020 ;
        RECT 1326.740 379.480 1327.000 379.740 ;
        RECT 1327.200 379.480 1327.460 379.740 ;
        RECT 1326.740 330.860 1327.000 331.120 ;
        RECT 1327.200 330.860 1327.460 331.120 ;
        RECT 1327.200 186.700 1327.460 186.960 ;
        RECT 1326.740 186.360 1327.000 186.620 ;
        RECT 1326.740 110.540 1327.000 110.800 ;
        RECT 1327.200 109.860 1327.460 110.120 ;
        RECT 668.940 25.540 669.200 25.800 ;
        RECT 1326.740 25.540 1327.000 25.800 ;
      LAYER met2 ;
        RECT 1330.410 1700.410 1330.690 1704.000 ;
        RECT 1329.560 1700.270 1330.690 1700.410 ;
        RECT 1329.560 1642.530 1329.700 1700.270 ;
        RECT 1330.410 1700.000 1330.690 1700.270 ;
        RECT 1326.740 1642.210 1327.000 1642.530 ;
        RECT 1329.500 1642.210 1329.760 1642.530 ;
        RECT 1326.800 1545.970 1326.940 1642.210 ;
        RECT 1326.740 1545.650 1327.000 1545.970 ;
        RECT 1327.200 1545.650 1327.460 1545.970 ;
        RECT 1327.260 1425.010 1327.400 1545.650 ;
        RECT 1327.260 1424.870 1327.860 1425.010 ;
        RECT 1327.720 1401.470 1327.860 1424.870 ;
        RECT 1327.660 1401.150 1327.920 1401.470 ;
        RECT 1326.740 1400.810 1327.000 1401.130 ;
        RECT 1326.800 1368.150 1326.940 1400.810 ;
        RECT 1326.740 1367.830 1327.000 1368.150 ;
        RECT 1327.660 1345.050 1327.920 1345.370 ;
        RECT 1327.720 1297.430 1327.860 1345.050 ;
        RECT 1327.200 1297.110 1327.460 1297.430 ;
        RECT 1327.660 1297.110 1327.920 1297.430 ;
        RECT 1327.260 1249.150 1327.400 1297.110 ;
        RECT 1326.740 1248.830 1327.000 1249.150 ;
        RECT 1327.200 1248.830 1327.460 1249.150 ;
        RECT 1326.800 1110.965 1326.940 1248.830 ;
        RECT 1326.730 1110.595 1327.010 1110.965 ;
        RECT 1327.190 1109.915 1327.470 1110.285 ;
        RECT 1327.260 814.630 1327.400 1109.915 ;
        RECT 1327.200 814.310 1327.460 814.630 ;
        RECT 1326.740 813.970 1327.000 814.290 ;
        RECT 1326.800 710.590 1326.940 813.970 ;
        RECT 1326.740 710.270 1327.000 710.590 ;
        RECT 1327.200 642.270 1327.460 642.590 ;
        RECT 1327.260 607.230 1327.400 642.270 ;
        RECT 1327.200 606.910 1327.460 607.230 ;
        RECT 1326.740 558.970 1327.000 559.290 ;
        RECT 1326.800 537.190 1326.940 558.970 ;
        RECT 1326.740 536.870 1327.000 537.190 ;
        RECT 1327.660 475.670 1327.920 475.990 ;
        RECT 1327.720 428.050 1327.860 475.670 ;
        RECT 1327.200 427.730 1327.460 428.050 ;
        RECT 1327.660 427.730 1327.920 428.050 ;
        RECT 1327.260 379.770 1327.400 427.730 ;
        RECT 1326.740 379.450 1327.000 379.770 ;
        RECT 1327.200 379.450 1327.460 379.770 ;
        RECT 1326.800 331.150 1326.940 379.450 ;
        RECT 1326.740 330.830 1327.000 331.150 ;
        RECT 1327.200 330.830 1327.460 331.150 ;
        RECT 1327.260 186.990 1327.400 330.830 ;
        RECT 1327.200 186.670 1327.460 186.990 ;
        RECT 1326.740 186.330 1327.000 186.650 ;
        RECT 1326.800 110.830 1326.940 186.330 ;
        RECT 1326.740 110.510 1327.000 110.830 ;
        RECT 1327.200 109.830 1327.460 110.150 ;
        RECT 1327.260 41.210 1327.400 109.830 ;
        RECT 1326.800 41.070 1327.400 41.210 ;
        RECT 1326.800 25.830 1326.940 41.070 ;
        RECT 668.940 25.510 669.200 25.830 ;
        RECT 1326.740 25.510 1327.000 25.830 ;
        RECT 669.000 2.400 669.140 25.510 ;
        RECT 668.790 -4.800 669.350 2.400 ;
      LAYER via2 ;
        RECT 1326.730 1110.640 1327.010 1110.920 ;
        RECT 1327.190 1109.960 1327.470 1110.240 ;
      LAYER met3 ;
        RECT 1326.705 1110.930 1327.035 1110.945 ;
        RECT 1326.705 1110.615 1327.250 1110.930 ;
        RECT 1326.950 1110.265 1327.250 1110.615 ;
        RECT 1326.950 1109.950 1327.495 1110.265 ;
        RECT 1327.165 1109.935 1327.495 1109.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1168.470 25.060 1168.790 25.120 ;
        RECT 1464.250 25.060 1464.570 25.120 ;
        RECT 1168.470 24.920 1464.570 25.060 ;
        RECT 1168.470 24.860 1168.790 24.920 ;
        RECT 1464.250 24.860 1464.570 24.920 ;
      LAYER via ;
        RECT 1168.500 24.860 1168.760 25.120 ;
        RECT 1464.280 24.860 1464.540 25.120 ;
      LAYER met2 ;
        RECT 1465.190 1700.410 1465.470 1704.000 ;
        RECT 1464.340 1700.270 1465.470 1700.410 ;
        RECT 1464.340 25.150 1464.480 1700.270 ;
        RECT 1465.190 1700.000 1465.470 1700.270 ;
        RECT 1168.500 24.830 1168.760 25.150 ;
        RECT 1464.280 24.830 1464.540 25.150 ;
        RECT 1168.560 2.400 1168.700 24.830 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1185.830 -4.800 1186.390 0.300 ;
=======
        RECT 1469.790 1700.000 1470.070 1704.000 ;
        RECT 1469.860 16.845 1470.000 1700.000 ;
        RECT 1185.970 16.475 1186.250 16.845 ;
        RECT 1469.790 16.475 1470.070 16.845 ;
        RECT 1186.040 2.400 1186.180 16.475 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
      LAYER via2 ;
        RECT 1185.970 16.520 1186.250 16.800 ;
        RECT 1469.790 16.520 1470.070 16.800 ;
      LAYER met3 ;
        RECT 1185.945 16.810 1186.275 16.825 ;
        RECT 1469.765 16.810 1470.095 16.825 ;
        RECT 1185.945 16.510 1470.095 16.810 ;
        RECT 1185.945 16.495 1186.275 16.510 ;
        RECT 1469.765 16.495 1470.095 16.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1470.690 1678.140 1471.010 1678.200 ;
        RECT 1473.450 1678.140 1473.770 1678.200 ;
        RECT 1470.690 1678.000 1473.770 1678.140 ;
        RECT 1470.690 1677.940 1471.010 1678.000 ;
        RECT 1473.450 1677.940 1473.770 1678.000 ;
      LAYER via ;
        RECT 1470.720 1677.940 1470.980 1678.200 ;
        RECT 1473.480 1677.940 1473.740 1678.200 ;
      LAYER met2 ;
        RECT 1474.850 1700.410 1475.130 1704.000 ;
        RECT 1473.540 1700.270 1475.130 1700.410 ;
        RECT 1473.540 1678.230 1473.680 1700.270 ;
        RECT 1474.850 1700.000 1475.130 1700.270 ;
        RECT 1470.720 1677.910 1470.980 1678.230 ;
        RECT 1473.480 1677.910 1473.740 1678.230 ;
        RECT 1470.780 19.565 1470.920 1677.910 ;
        RECT 1203.910 19.195 1204.190 19.565 ;
        RECT 1470.710 19.195 1470.990 19.565 ;
        RECT 1203.980 2.400 1204.120 19.195 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
      LAYER via2 ;
        RECT 1203.910 19.240 1204.190 19.520 ;
        RECT 1470.710 19.240 1470.990 19.520 ;
      LAYER met3 ;
        RECT 1203.885 19.530 1204.215 19.545 ;
        RECT 1470.685 19.530 1471.015 19.545 ;
        RECT 1203.885 19.230 1471.015 19.530 ;
        RECT 1203.885 19.215 1204.215 19.230 ;
        RECT 1470.685 19.215 1471.015 19.230 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 0.300 ;
=======
      LAYER li1 ;
        RECT 1422.925 14.025 1423.095 17.935 ;
      LAYER mcon ;
        RECT 1422.925 17.765 1423.095 17.935 ;
      LAYER met1 ;
        RECT 1477.590 1666.240 1477.910 1666.300 ;
        RECT 1478.510 1666.240 1478.830 1666.300 ;
        RECT 1477.590 1666.100 1478.830 1666.240 ;
        RECT 1477.590 1666.040 1477.910 1666.100 ;
        RECT 1478.510 1666.040 1478.830 1666.100 ;
        RECT 1221.830 17.920 1222.150 17.980 ;
        RECT 1422.865 17.920 1423.155 17.965 ;
        RECT 1221.830 17.780 1423.155 17.920 ;
        RECT 1221.830 17.720 1222.150 17.780 ;
        RECT 1422.865 17.735 1423.155 17.780 ;
        RECT 1422.865 14.180 1423.155 14.225 ;
        RECT 1422.865 14.040 1471.380 14.180 ;
        RECT 1422.865 13.995 1423.155 14.040 ;
        RECT 1471.240 13.840 1471.380 14.040 ;
        RECT 1478.050 13.840 1478.370 13.900 ;
        RECT 1471.240 13.700 1478.370 13.840 ;
        RECT 1478.050 13.640 1478.370 13.700 ;
      LAYER via ;
        RECT 1477.620 1666.040 1477.880 1666.300 ;
        RECT 1478.540 1666.040 1478.800 1666.300 ;
        RECT 1221.860 17.720 1222.120 17.980 ;
        RECT 1478.080 13.640 1478.340 13.900 ;
      LAYER met2 ;
        RECT 1479.450 1700.410 1479.730 1704.000 ;
        RECT 1478.600 1700.270 1479.730 1700.410 ;
        RECT 1478.600 1666.330 1478.740 1700.270 ;
        RECT 1479.450 1700.000 1479.730 1700.270 ;
        RECT 1477.620 1666.010 1477.880 1666.330 ;
        RECT 1478.540 1666.010 1478.800 1666.330 ;
        RECT 1477.680 37.810 1477.820 1666.010 ;
        RECT 1477.680 37.670 1478.280 37.810 ;
        RECT 1221.860 17.690 1222.120 18.010 ;
        RECT 1221.920 2.400 1222.060 17.690 ;
        RECT 1478.140 13.930 1478.280 37.670 ;
        RECT 1478.080 13.610 1478.340 13.930 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 0.300 ;
=======
      LAYER li1 ;
        RECT 1463.865 18.445 1464.955 18.615 ;
      LAYER mcon ;
        RECT 1464.785 18.445 1464.955 18.615 ;
      LAYER met1 ;
        RECT 1239.770 18.600 1240.090 18.660 ;
        RECT 1463.805 18.600 1464.095 18.645 ;
        RECT 1239.770 18.460 1464.095 18.600 ;
        RECT 1239.770 18.400 1240.090 18.460 ;
        RECT 1463.805 18.415 1464.095 18.460 ;
        RECT 1464.725 18.600 1465.015 18.645 ;
        RECT 1484.950 18.600 1485.270 18.660 ;
        RECT 1464.725 18.460 1485.270 18.600 ;
        RECT 1464.725 18.415 1465.015 18.460 ;
        RECT 1484.950 18.400 1485.270 18.460 ;
      LAYER via ;
        RECT 1239.800 18.400 1240.060 18.660 ;
        RECT 1484.980 18.400 1485.240 18.660 ;
      LAYER met2 ;
        RECT 1484.510 1700.410 1484.790 1704.000 ;
        RECT 1484.510 1700.270 1485.180 1700.410 ;
        RECT 1484.510 1700.000 1484.790 1700.270 ;
        RECT 1485.040 18.690 1485.180 1700.270 ;
        RECT 1239.800 18.370 1240.060 18.690 ;
        RECT 1484.980 18.370 1485.240 18.690 ;
        RECT 1239.860 2.400 1240.000 18.370 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1484.030 1678.140 1484.350 1678.200 ;
        RECT 1488.170 1678.140 1488.490 1678.200 ;
        RECT 1484.030 1678.000 1488.490 1678.140 ;
        RECT 1484.030 1677.940 1484.350 1678.000 ;
        RECT 1488.170 1677.940 1488.490 1678.000 ;
        RECT 1257.250 25.400 1257.570 25.460 ;
        RECT 1484.030 25.400 1484.350 25.460 ;
        RECT 1257.250 25.260 1484.350 25.400 ;
        RECT 1257.250 25.200 1257.570 25.260 ;
        RECT 1484.030 25.200 1484.350 25.260 ;
      LAYER via ;
        RECT 1484.060 1677.940 1484.320 1678.200 ;
        RECT 1488.200 1677.940 1488.460 1678.200 ;
        RECT 1257.280 25.200 1257.540 25.460 ;
        RECT 1484.060 25.200 1484.320 25.460 ;
      LAYER met2 ;
        RECT 1489.110 1700.410 1489.390 1704.000 ;
        RECT 1488.260 1700.270 1489.390 1700.410 ;
        RECT 1488.260 1678.230 1488.400 1700.270 ;
        RECT 1489.110 1700.000 1489.390 1700.270 ;
        RECT 1484.060 1677.910 1484.320 1678.230 ;
        RECT 1488.200 1677.910 1488.460 1678.230 ;
        RECT 1484.120 25.490 1484.260 1677.910 ;
        RECT 1257.280 25.170 1257.540 25.490 ;
        RECT 1484.060 25.170 1484.320 25.490 ;
        RECT 1257.340 2.400 1257.480 25.170 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 0.300 ;
=======
      LAYER li1 ;
        RECT 1492.845 1393.745 1493.015 1401.055 ;
        RECT 1492.385 1290.385 1492.555 1304.495 ;
        RECT 1492.385 1152.345 1492.555 1183.795 ;
        RECT 1492.385 582.845 1492.555 620.755 ;
        RECT 1492.385 434.605 1492.555 475.915 ;
        RECT 1492.845 372.725 1493.015 420.835 ;
        RECT 1492.845 276.165 1493.015 324.275 ;
        RECT 1491.925 234.685 1492.095 255.935 ;
        RECT 1491.925 179.605 1492.095 227.715 ;
        RECT 1470.765 19.125 1471.395 19.295 ;
        RECT 1471.225 14.195 1471.395 19.125 ;
        RECT 1471.225 14.025 1471.855 14.195 ;
      LAYER mcon ;
        RECT 1492.845 1400.885 1493.015 1401.055 ;
        RECT 1492.385 1304.325 1492.555 1304.495 ;
        RECT 1492.385 1183.625 1492.555 1183.795 ;
        RECT 1492.385 620.585 1492.555 620.755 ;
        RECT 1492.385 475.745 1492.555 475.915 ;
        RECT 1492.845 420.665 1493.015 420.835 ;
        RECT 1492.845 324.105 1493.015 324.275 ;
        RECT 1491.925 255.765 1492.095 255.935 ;
        RECT 1491.925 227.545 1492.095 227.715 ;
        RECT 1471.685 14.025 1471.855 14.195 ;
      LAYER met1 ;
        RECT 1492.770 1607.900 1493.090 1608.160 ;
        RECT 1492.860 1607.480 1493.000 1607.900 ;
        RECT 1492.770 1607.220 1493.090 1607.480 ;
        RECT 1492.310 1442.520 1492.630 1442.580 ;
        RECT 1493.230 1442.520 1493.550 1442.580 ;
        RECT 1492.310 1442.380 1493.550 1442.520 ;
        RECT 1492.310 1442.320 1492.630 1442.380 ;
        RECT 1493.230 1442.320 1493.550 1442.380 ;
        RECT 1492.770 1401.040 1493.090 1401.100 ;
        RECT 1492.575 1400.900 1493.090 1401.040 ;
        RECT 1492.770 1400.840 1493.090 1400.900 ;
        RECT 1492.770 1393.900 1493.090 1393.960 ;
        RECT 1492.575 1393.760 1493.090 1393.900 ;
        RECT 1492.770 1393.700 1493.090 1393.760 ;
        RECT 1492.310 1304.480 1492.630 1304.540 ;
        RECT 1492.115 1304.340 1492.630 1304.480 ;
        RECT 1492.310 1304.280 1492.630 1304.340 ;
        RECT 1492.310 1290.540 1492.630 1290.600 ;
        RECT 1492.115 1290.400 1492.630 1290.540 ;
        RECT 1492.310 1290.340 1492.630 1290.400 ;
        RECT 1491.850 1242.260 1492.170 1242.320 ;
        RECT 1492.310 1242.260 1492.630 1242.320 ;
        RECT 1491.850 1242.120 1492.630 1242.260 ;
        RECT 1491.850 1242.060 1492.170 1242.120 ;
        RECT 1492.310 1242.060 1492.630 1242.120 ;
        RECT 1491.850 1241.580 1492.170 1241.640 ;
        RECT 1492.310 1241.580 1492.630 1241.640 ;
        RECT 1491.850 1241.440 1492.630 1241.580 ;
        RECT 1491.850 1241.380 1492.170 1241.440 ;
        RECT 1492.310 1241.380 1492.630 1241.440 ;
        RECT 1492.325 1183.780 1492.615 1183.825 ;
        RECT 1492.770 1183.780 1493.090 1183.840 ;
        RECT 1492.325 1183.640 1493.090 1183.780 ;
        RECT 1492.325 1183.595 1492.615 1183.640 ;
        RECT 1492.770 1183.580 1493.090 1183.640 ;
        RECT 1492.310 1152.500 1492.630 1152.560 ;
        RECT 1492.115 1152.360 1492.630 1152.500 ;
        RECT 1492.310 1152.300 1492.630 1152.360 ;
        RECT 1491.850 724.440 1492.170 724.500 ;
        RECT 1492.770 724.440 1493.090 724.500 ;
        RECT 1491.850 724.300 1493.090 724.440 ;
        RECT 1491.850 724.240 1492.170 724.300 ;
        RECT 1492.770 724.240 1493.090 724.300 ;
        RECT 1491.850 676.640 1492.170 676.900 ;
        RECT 1491.940 676.220 1492.080 676.640 ;
        RECT 1491.850 675.960 1492.170 676.220 ;
        RECT 1492.310 620.740 1492.630 620.800 ;
        RECT 1492.115 620.600 1492.630 620.740 ;
        RECT 1492.310 620.540 1492.630 620.600 ;
        RECT 1492.310 583.000 1492.630 583.060 ;
        RECT 1492.115 582.860 1492.630 583.000 ;
        RECT 1492.310 582.800 1492.630 582.860 ;
        RECT 1493.230 483.380 1493.550 483.440 ;
        RECT 1492.400 483.240 1493.550 483.380 ;
        RECT 1492.400 483.100 1492.540 483.240 ;
        RECT 1493.230 483.180 1493.550 483.240 ;
        RECT 1492.310 482.840 1492.630 483.100 ;
        RECT 1492.310 475.900 1492.630 475.960 ;
        RECT 1492.115 475.760 1492.630 475.900 ;
        RECT 1492.310 475.700 1492.630 475.760 ;
        RECT 1492.325 434.760 1492.615 434.805 ;
        RECT 1492.770 434.760 1493.090 434.820 ;
        RECT 1492.325 434.620 1493.090 434.760 ;
        RECT 1492.325 434.575 1492.615 434.620 ;
        RECT 1492.770 434.560 1493.090 434.620 ;
        RECT 1492.770 420.820 1493.090 420.880 ;
        RECT 1492.575 420.680 1493.090 420.820 ;
        RECT 1492.770 420.620 1493.090 420.680 ;
        RECT 1492.770 372.880 1493.090 372.940 ;
        RECT 1492.575 372.740 1493.090 372.880 ;
        RECT 1492.770 372.680 1493.090 372.740 ;
        RECT 1492.770 324.260 1493.090 324.320 ;
        RECT 1492.575 324.120 1493.090 324.260 ;
        RECT 1492.770 324.060 1493.090 324.120 ;
        RECT 1492.770 276.320 1493.090 276.380 ;
        RECT 1492.575 276.180 1493.090 276.320 ;
        RECT 1492.770 276.120 1493.090 276.180 ;
        RECT 1491.865 255.920 1492.155 255.965 ;
        RECT 1492.770 255.920 1493.090 255.980 ;
        RECT 1491.865 255.780 1493.090 255.920 ;
        RECT 1491.865 255.735 1492.155 255.780 ;
        RECT 1492.770 255.720 1493.090 255.780 ;
        RECT 1491.850 234.840 1492.170 234.900 ;
        RECT 1491.655 234.700 1492.170 234.840 ;
        RECT 1491.850 234.640 1492.170 234.700 ;
        RECT 1491.850 227.700 1492.170 227.760 ;
        RECT 1491.655 227.560 1492.170 227.700 ;
        RECT 1491.850 227.500 1492.170 227.560 ;
        RECT 1491.865 179.760 1492.155 179.805 ;
        RECT 1492.310 179.760 1492.630 179.820 ;
        RECT 1491.865 179.620 1492.630 179.760 ;
        RECT 1491.865 179.575 1492.155 179.620 ;
        RECT 1492.310 179.560 1492.630 179.620 ;
        RECT 1492.310 96.600 1492.630 96.860 ;
        RECT 1492.400 96.120 1492.540 96.600 ;
        RECT 1492.770 96.120 1493.090 96.180 ;
        RECT 1492.400 95.980 1493.090 96.120 ;
        RECT 1492.770 95.920 1493.090 95.980 ;
        RECT 1492.310 48.520 1492.630 48.580 ;
        RECT 1492.770 48.520 1493.090 48.580 ;
        RECT 1492.310 48.380 1493.090 48.520 ;
        RECT 1492.310 48.320 1492.630 48.380 ;
        RECT 1492.770 48.320 1493.090 48.380 ;
        RECT 1470.705 19.280 1470.995 19.325 ;
        RECT 1463.880 19.140 1470.995 19.280 ;
        RECT 1275.190 18.940 1275.510 19.000 ;
        RECT 1463.880 18.940 1464.020 19.140 ;
        RECT 1470.705 19.095 1470.995 19.140 ;
        RECT 1275.190 18.800 1464.020 18.940 ;
        RECT 1275.190 18.740 1275.510 18.800 ;
        RECT 1471.625 14.180 1471.915 14.225 ;
        RECT 1492.310 14.180 1492.630 14.240 ;
        RECT 1471.625 14.040 1492.630 14.180 ;
        RECT 1471.625 13.995 1471.915 14.040 ;
        RECT 1492.310 13.980 1492.630 14.040 ;
      LAYER via ;
        RECT 1492.800 1607.900 1493.060 1608.160 ;
        RECT 1492.800 1607.220 1493.060 1607.480 ;
        RECT 1492.340 1442.320 1492.600 1442.580 ;
        RECT 1493.260 1442.320 1493.520 1442.580 ;
        RECT 1492.800 1400.840 1493.060 1401.100 ;
        RECT 1492.800 1393.700 1493.060 1393.960 ;
        RECT 1492.340 1304.280 1492.600 1304.540 ;
        RECT 1492.340 1290.340 1492.600 1290.600 ;
        RECT 1491.880 1242.060 1492.140 1242.320 ;
        RECT 1492.340 1242.060 1492.600 1242.320 ;
        RECT 1491.880 1241.380 1492.140 1241.640 ;
        RECT 1492.340 1241.380 1492.600 1241.640 ;
        RECT 1492.800 1183.580 1493.060 1183.840 ;
        RECT 1492.340 1152.300 1492.600 1152.560 ;
        RECT 1491.880 724.240 1492.140 724.500 ;
        RECT 1492.800 724.240 1493.060 724.500 ;
        RECT 1491.880 676.640 1492.140 676.900 ;
        RECT 1491.880 675.960 1492.140 676.220 ;
        RECT 1492.340 620.540 1492.600 620.800 ;
        RECT 1492.340 582.800 1492.600 583.060 ;
        RECT 1493.260 483.180 1493.520 483.440 ;
        RECT 1492.340 482.840 1492.600 483.100 ;
        RECT 1492.340 475.700 1492.600 475.960 ;
        RECT 1492.800 434.560 1493.060 434.820 ;
        RECT 1492.800 420.620 1493.060 420.880 ;
        RECT 1492.800 372.680 1493.060 372.940 ;
        RECT 1492.800 324.060 1493.060 324.320 ;
        RECT 1492.800 276.120 1493.060 276.380 ;
        RECT 1492.800 255.720 1493.060 255.980 ;
        RECT 1491.880 234.640 1492.140 234.900 ;
        RECT 1491.880 227.500 1492.140 227.760 ;
        RECT 1492.340 179.560 1492.600 179.820 ;
        RECT 1492.340 96.600 1492.600 96.860 ;
        RECT 1492.800 95.920 1493.060 96.180 ;
        RECT 1492.340 48.320 1492.600 48.580 ;
        RECT 1492.800 48.320 1493.060 48.580 ;
        RECT 1275.220 18.740 1275.480 19.000 ;
        RECT 1492.340 13.980 1492.600 14.240 ;
      LAYER met2 ;
        RECT 1494.170 1700.410 1494.450 1704.000 ;
        RECT 1493.320 1700.270 1494.450 1700.410 ;
        RECT 1493.320 1678.480 1493.460 1700.270 ;
        RECT 1494.170 1700.000 1494.450 1700.270 ;
        RECT 1492.400 1678.340 1493.460 1678.480 ;
        RECT 1492.400 1655.530 1492.540 1678.340 ;
        RECT 1492.400 1655.390 1493.000 1655.530 ;
        RECT 1492.860 1608.190 1493.000 1655.390 ;
        RECT 1492.800 1607.870 1493.060 1608.190 ;
        RECT 1492.800 1607.190 1493.060 1607.510 ;
        RECT 1492.860 1497.770 1493.000 1607.190 ;
        RECT 1492.400 1497.630 1493.000 1497.770 ;
        RECT 1492.400 1442.610 1492.540 1497.630 ;
        RECT 1492.340 1442.290 1492.600 1442.610 ;
        RECT 1493.260 1442.290 1493.520 1442.610 ;
        RECT 1493.320 1442.010 1493.460 1442.290 ;
        RECT 1492.860 1441.870 1493.460 1442.010 ;
        RECT 1492.860 1401.130 1493.000 1441.870 ;
        RECT 1492.800 1400.810 1493.060 1401.130 ;
        RECT 1492.800 1393.670 1493.060 1393.990 ;
        RECT 1492.860 1366.530 1493.000 1393.670 ;
        RECT 1492.860 1366.390 1493.460 1366.530 ;
        RECT 1493.320 1343.410 1493.460 1366.390 ;
        RECT 1492.860 1343.270 1493.460 1343.410 ;
        RECT 1492.860 1338.650 1493.000 1343.270 ;
        RECT 1492.400 1338.510 1493.000 1338.650 ;
        RECT 1492.400 1304.570 1492.540 1338.510 ;
        RECT 1492.340 1304.250 1492.600 1304.570 ;
        RECT 1492.340 1290.310 1492.600 1290.630 ;
        RECT 1492.400 1242.350 1492.540 1290.310 ;
        RECT 1491.880 1242.030 1492.140 1242.350 ;
        RECT 1492.340 1242.030 1492.600 1242.350 ;
        RECT 1491.940 1241.670 1492.080 1242.030 ;
        RECT 1491.880 1241.350 1492.140 1241.670 ;
        RECT 1492.340 1241.350 1492.600 1241.670 ;
        RECT 1492.400 1193.810 1492.540 1241.350 ;
        RECT 1492.400 1193.670 1493.000 1193.810 ;
        RECT 1492.860 1183.870 1493.000 1193.670 ;
        RECT 1492.800 1183.550 1493.060 1183.870 ;
        RECT 1492.340 1152.270 1492.600 1152.590 ;
        RECT 1492.400 1124.450 1492.540 1152.270 ;
        RECT 1492.400 1124.310 1493.000 1124.450 ;
        RECT 1492.860 883.050 1493.000 1124.310 ;
        RECT 1492.400 882.910 1493.000 883.050 ;
        RECT 1492.400 881.690 1492.540 882.910 ;
        RECT 1492.400 881.550 1493.000 881.690 ;
        RECT 1492.860 786.490 1493.000 881.550 ;
        RECT 1492.400 786.350 1493.000 786.490 ;
        RECT 1492.400 785.130 1492.540 786.350 ;
        RECT 1492.400 784.990 1493.000 785.130 ;
        RECT 1492.860 724.530 1493.000 784.990 ;
        RECT 1491.880 724.210 1492.140 724.530 ;
        RECT 1492.800 724.210 1493.060 724.530 ;
        RECT 1491.940 676.930 1492.080 724.210 ;
        RECT 1491.880 676.610 1492.140 676.930 ;
        RECT 1491.880 675.930 1492.140 676.250 ;
        RECT 1491.940 651.170 1492.080 675.930 ;
        RECT 1491.940 651.030 1492.540 651.170 ;
        RECT 1492.400 620.830 1492.540 651.030 ;
        RECT 1492.340 620.510 1492.600 620.830 ;
        RECT 1492.340 582.770 1492.600 583.090 ;
        RECT 1492.400 531.605 1492.540 582.770 ;
        RECT 1492.330 531.235 1492.610 531.605 ;
        RECT 1493.250 530.555 1493.530 530.925 ;
        RECT 1493.320 483.470 1493.460 530.555 ;
        RECT 1493.260 483.150 1493.520 483.470 ;
        RECT 1492.340 482.810 1492.600 483.130 ;
        RECT 1492.400 475.990 1492.540 482.810 ;
        RECT 1492.340 475.670 1492.600 475.990 ;
        RECT 1492.800 434.530 1493.060 434.850 ;
        RECT 1492.860 420.910 1493.000 434.530 ;
        RECT 1492.800 420.590 1493.060 420.910 ;
        RECT 1492.800 372.650 1493.060 372.970 ;
        RECT 1492.860 324.350 1493.000 372.650 ;
        RECT 1492.800 324.030 1493.060 324.350 ;
        RECT 1492.800 276.090 1493.060 276.410 ;
        RECT 1492.860 256.010 1493.000 276.090 ;
        RECT 1492.800 255.690 1493.060 256.010 ;
        RECT 1491.880 234.610 1492.140 234.930 ;
        RECT 1491.940 227.790 1492.080 234.610 ;
        RECT 1491.880 227.470 1492.140 227.790 ;
        RECT 1492.340 179.530 1492.600 179.850 ;
        RECT 1492.400 96.890 1492.540 179.530 ;
        RECT 1492.340 96.570 1492.600 96.890 ;
        RECT 1492.800 95.890 1493.060 96.210 ;
        RECT 1492.860 48.610 1493.000 95.890 ;
        RECT 1492.340 48.290 1492.600 48.610 ;
        RECT 1492.800 48.290 1493.060 48.610 ;
        RECT 1275.220 18.710 1275.480 19.030 ;
        RECT 1275.280 2.400 1275.420 18.710 ;
        RECT 1492.400 14.270 1492.540 48.290 ;
        RECT 1492.340 13.950 1492.600 14.270 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
      LAYER via2 ;
        RECT 1492.330 531.280 1492.610 531.560 ;
        RECT 1493.250 530.600 1493.530 530.880 ;
      LAYER met3 ;
        RECT 1492.305 531.570 1492.635 531.585 ;
        RECT 1492.305 531.255 1492.850 531.570 ;
        RECT 1492.550 530.890 1492.850 531.255 ;
        RECT 1493.225 530.890 1493.555 530.905 ;
        RECT 1492.550 530.590 1493.555 530.890 ;
        RECT 1493.225 530.575 1493.555 530.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 0.300 ;
=======
      LAYER li1 ;
        RECT 1463.405 18.275 1463.575 19.295 ;
        RECT 1463.405 18.105 1465.875 18.275 ;
        RECT 1465.705 17.085 1465.875 18.105 ;
      LAYER mcon ;
        RECT 1463.405 19.125 1463.575 19.295 ;
      LAYER met1 ;
        RECT 1293.130 19.280 1293.450 19.340 ;
        RECT 1463.345 19.280 1463.635 19.325 ;
        RECT 1293.130 19.140 1463.635 19.280 ;
        RECT 1293.130 19.080 1293.450 19.140 ;
        RECT 1463.345 19.095 1463.635 19.140 ;
        RECT 1487.250 18.260 1487.570 18.320 ;
        RECT 1498.750 18.260 1499.070 18.320 ;
        RECT 1487.250 18.120 1499.070 18.260 ;
        RECT 1487.250 18.060 1487.570 18.120 ;
        RECT 1498.750 18.060 1499.070 18.120 ;
        RECT 1465.645 17.240 1465.935 17.285 ;
        RECT 1484.030 17.240 1484.350 17.300 ;
        RECT 1465.645 17.100 1484.350 17.240 ;
        RECT 1465.645 17.055 1465.935 17.100 ;
        RECT 1484.030 17.040 1484.350 17.100 ;
      LAYER via ;
        RECT 1293.160 19.080 1293.420 19.340 ;
        RECT 1487.280 18.060 1487.540 18.320 ;
        RECT 1498.780 18.060 1499.040 18.320 ;
        RECT 1484.060 17.040 1484.320 17.300 ;
      LAYER met2 ;
        RECT 1498.770 1700.000 1499.050 1704.000 ;
        RECT 1293.160 19.050 1293.420 19.370 ;
        RECT 1293.220 2.400 1293.360 19.050 ;
        RECT 1498.840 18.350 1498.980 1700.000 ;
        RECT 1484.120 17.950 1485.180 18.090 ;
        RECT 1487.280 18.030 1487.540 18.350 ;
        RECT 1498.780 18.030 1499.040 18.350 ;
        RECT 1484.120 17.330 1484.260 17.950 ;
        RECT 1485.040 17.410 1485.180 17.950 ;
        RECT 1487.340 17.410 1487.480 18.030 ;
        RECT 1484.060 17.010 1484.320 17.330 ;
        RECT 1485.040 17.270 1487.480 17.410 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 0.300 ;
=======
      LAYER met1 ;
        RECT 1498.290 1678.140 1498.610 1678.200 ;
        RECT 1502.430 1678.140 1502.750 1678.200 ;
        RECT 1498.290 1678.000 1502.750 1678.140 ;
        RECT 1498.290 1677.940 1498.610 1678.000 ;
        RECT 1502.430 1677.940 1502.750 1678.000 ;
        RECT 1311.070 19.620 1311.390 19.680 ;
        RECT 1311.070 19.480 1471.380 19.620 ;
        RECT 1311.070 19.420 1311.390 19.480 ;
        RECT 1471.240 19.280 1471.380 19.480 ;
        RECT 1471.240 19.140 1485.640 19.280 ;
        RECT 1485.500 18.600 1485.640 19.140 ;
        RECT 1498.290 18.600 1498.610 18.660 ;
        RECT 1485.500 18.460 1498.610 18.600 ;
        RECT 1498.290 18.400 1498.610 18.460 ;
      LAYER via ;
        RECT 1498.320 1677.940 1498.580 1678.200 ;
        RECT 1502.460 1677.940 1502.720 1678.200 ;
        RECT 1311.100 19.420 1311.360 19.680 ;
        RECT 1498.320 18.400 1498.580 18.660 ;
      LAYER met2 ;
        RECT 1503.830 1700.410 1504.110 1704.000 ;
        RECT 1502.520 1700.270 1504.110 1700.410 ;
        RECT 1502.520 1678.230 1502.660 1700.270 ;
        RECT 1503.830 1700.000 1504.110 1700.270 ;
        RECT 1498.320 1677.910 1498.580 1678.230 ;
        RECT 1502.460 1677.910 1502.720 1678.230 ;
        RECT 1311.100 19.390 1311.360 19.710 ;
        RECT 1311.160 2.400 1311.300 19.390 ;
        RECT 1498.380 18.690 1498.520 1677.910 ;
        RECT 1498.320 18.370 1498.580 18.690 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 0.300 ;
=======
      LAYER li1 ;
        RECT 1505.725 1338.665 1505.895 1366.035 ;
        RECT 1505.725 766.105 1505.895 814.215 ;
      LAYER mcon ;
        RECT 1505.725 1365.865 1505.895 1366.035 ;
        RECT 1505.725 814.045 1505.895 814.215 ;
      LAYER met1 ;
        RECT 1505.650 1642.440 1505.970 1642.500 ;
        RECT 1507.030 1642.440 1507.350 1642.500 ;
        RECT 1505.650 1642.300 1507.350 1642.440 ;
        RECT 1505.650 1642.240 1505.970 1642.300 ;
        RECT 1507.030 1642.240 1507.350 1642.300 ;
        RECT 1505.650 1366.020 1505.970 1366.080 ;
        RECT 1505.455 1365.880 1505.970 1366.020 ;
        RECT 1505.650 1365.820 1505.970 1365.880 ;
        RECT 1505.650 1338.820 1505.970 1338.880 ;
        RECT 1505.455 1338.680 1505.970 1338.820 ;
        RECT 1505.650 1338.620 1505.970 1338.680 ;
        RECT 1505.650 1257.700 1505.970 1257.960 ;
        RECT 1505.740 1257.280 1505.880 1257.700 ;
        RECT 1505.650 1257.020 1505.970 1257.280 ;
        RECT 1504.730 886.620 1505.050 886.680 ;
        RECT 1505.650 886.620 1505.970 886.680 ;
        RECT 1504.730 886.480 1505.970 886.620 ;
        RECT 1504.730 886.420 1505.050 886.480 ;
        RECT 1505.650 886.420 1505.970 886.480 ;
        RECT 1505.650 814.200 1505.970 814.260 ;
        RECT 1505.455 814.060 1505.970 814.200 ;
        RECT 1505.650 814.000 1505.970 814.060 ;
        RECT 1505.650 766.260 1505.970 766.320 ;
        RECT 1505.455 766.120 1505.970 766.260 ;
        RECT 1505.650 766.060 1505.970 766.120 ;
        RECT 1506.110 676.300 1506.430 676.560 ;
        RECT 1506.200 675.820 1506.340 676.300 ;
        RECT 1506.570 675.820 1506.890 675.880 ;
        RECT 1506.200 675.680 1506.890 675.820 ;
        RECT 1506.570 675.620 1506.890 675.680 ;
        RECT 1505.650 593.340 1505.970 593.600 ;
        RECT 1505.740 592.920 1505.880 593.340 ;
        RECT 1505.650 592.660 1505.970 592.920 ;
        RECT 1505.190 62.460 1505.510 62.520 ;
        RECT 1504.820 62.320 1505.510 62.460 ;
        RECT 1504.820 62.180 1504.960 62.320 ;
        RECT 1505.190 62.260 1505.510 62.320 ;
        RECT 1504.730 61.920 1505.050 62.180 ;
        RECT 1329.010 25.740 1329.330 25.800 ;
        RECT 1504.730 25.740 1505.050 25.800 ;
        RECT 1329.010 25.600 1505.050 25.740 ;
        RECT 1329.010 25.540 1329.330 25.600 ;
        RECT 1504.730 25.540 1505.050 25.600 ;
      LAYER via ;
        RECT 1505.680 1642.240 1505.940 1642.500 ;
        RECT 1507.060 1642.240 1507.320 1642.500 ;
        RECT 1505.680 1365.820 1505.940 1366.080 ;
        RECT 1505.680 1338.620 1505.940 1338.880 ;
        RECT 1505.680 1257.700 1505.940 1257.960 ;
        RECT 1505.680 1257.020 1505.940 1257.280 ;
        RECT 1504.760 886.420 1505.020 886.680 ;
        RECT 1505.680 886.420 1505.940 886.680 ;
        RECT 1505.680 814.000 1505.940 814.260 ;
        RECT 1505.680 766.060 1505.940 766.320 ;
        RECT 1506.140 676.300 1506.400 676.560 ;
        RECT 1506.600 675.620 1506.860 675.880 ;
        RECT 1505.680 593.340 1505.940 593.600 ;
        RECT 1505.680 592.660 1505.940 592.920 ;
        RECT 1505.220 62.260 1505.480 62.520 ;
        RECT 1504.760 61.920 1505.020 62.180 ;
        RECT 1329.040 25.540 1329.300 25.800 ;
        RECT 1504.760 25.540 1505.020 25.800 ;
      LAYER met2 ;
        RECT 1508.430 1700.410 1508.710 1704.000 ;
        RECT 1507.580 1700.270 1508.710 1700.410 ;
        RECT 1507.580 1672.530 1507.720 1700.270 ;
        RECT 1508.430 1700.000 1508.710 1700.270 ;
        RECT 1507.120 1672.390 1507.720 1672.530 ;
        RECT 1507.120 1642.530 1507.260 1672.390 ;
        RECT 1505.680 1642.210 1505.940 1642.530 ;
        RECT 1507.060 1642.210 1507.320 1642.530 ;
        RECT 1505.740 1366.110 1505.880 1642.210 ;
        RECT 1505.680 1365.790 1505.940 1366.110 ;
        RECT 1505.680 1338.590 1505.940 1338.910 ;
        RECT 1505.740 1257.990 1505.880 1338.590 ;
        RECT 1505.680 1257.670 1505.940 1257.990 ;
        RECT 1505.680 1256.990 1505.940 1257.310 ;
        RECT 1505.740 1076.850 1505.880 1256.990 ;
        RECT 1505.280 1076.710 1505.880 1076.850 ;
        RECT 1505.280 1076.170 1505.420 1076.710 ;
        RECT 1505.280 1076.030 1505.880 1076.170 ;
        RECT 1505.740 886.710 1505.880 1076.030 ;
        RECT 1504.760 886.390 1505.020 886.710 ;
        RECT 1505.680 886.390 1505.940 886.710 ;
        RECT 1504.820 862.765 1504.960 886.390 ;
        RECT 1504.750 862.395 1505.030 862.765 ;
        RECT 1505.670 862.395 1505.950 862.765 ;
        RECT 1505.740 814.290 1505.880 862.395 ;
        RECT 1505.680 813.970 1505.940 814.290 ;
        RECT 1505.680 766.030 1505.940 766.350 ;
        RECT 1505.740 749.090 1505.880 766.030 ;
        RECT 1505.740 748.950 1506.800 749.090 ;
        RECT 1506.660 724.610 1506.800 748.950 ;
        RECT 1506.200 724.470 1506.800 724.610 ;
        RECT 1506.200 676.590 1506.340 724.470 ;
        RECT 1506.140 676.270 1506.400 676.590 ;
        RECT 1506.600 675.590 1506.860 675.910 ;
        RECT 1506.660 628.165 1506.800 675.590 ;
        RECT 1505.670 627.795 1505.950 628.165 ;
        RECT 1506.590 627.795 1506.870 628.165 ;
        RECT 1505.740 593.630 1505.880 627.795 ;
        RECT 1505.680 593.310 1505.940 593.630 ;
        RECT 1505.680 592.630 1505.940 592.950 ;
        RECT 1505.740 303.690 1505.880 592.630 ;
        RECT 1505.280 303.550 1505.880 303.690 ;
        RECT 1505.280 303.010 1505.420 303.550 ;
        RECT 1505.280 302.870 1505.880 303.010 ;
        RECT 1505.740 207.130 1505.880 302.870 ;
        RECT 1505.280 206.990 1505.880 207.130 ;
        RECT 1505.280 206.450 1505.420 206.990 ;
        RECT 1505.280 206.310 1505.880 206.450 ;
        RECT 1505.740 110.570 1505.880 206.310 ;
        RECT 1505.280 110.430 1505.880 110.570 ;
        RECT 1505.280 62.550 1505.420 110.430 ;
        RECT 1505.220 62.230 1505.480 62.550 ;
        RECT 1504.760 61.890 1505.020 62.210 ;
        RECT 1504.820 25.830 1504.960 61.890 ;
        RECT 1329.040 25.510 1329.300 25.830 ;
        RECT 1504.760 25.510 1505.020 25.830 ;
        RECT 1329.100 2.400 1329.240 25.510 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
      LAYER via2 ;
        RECT 1504.750 862.440 1505.030 862.720 ;
        RECT 1505.670 862.440 1505.950 862.720 ;
        RECT 1505.670 627.840 1505.950 628.120 ;
        RECT 1506.590 627.840 1506.870 628.120 ;
      LAYER met3 ;
        RECT 1504.725 862.730 1505.055 862.745 ;
        RECT 1505.645 862.730 1505.975 862.745 ;
        RECT 1504.725 862.430 1505.975 862.730 ;
        RECT 1504.725 862.415 1505.055 862.430 ;
        RECT 1505.645 862.415 1505.975 862.430 ;
        RECT 1505.645 628.130 1505.975 628.145 ;
        RECT 1506.565 628.130 1506.895 628.145 ;
        RECT 1505.645 627.830 1506.895 628.130 ;
        RECT 1505.645 627.815 1505.975 627.830 ;
        RECT 1506.565 627.815 1506.895 627.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 0.300 ;
=======
      LAYER met1 ;
        RECT 686.390 26.080 686.710 26.140 ;
        RECT 1334.070 26.080 1334.390 26.140 ;
        RECT 686.390 25.940 1334.390 26.080 ;
        RECT 686.390 25.880 686.710 25.940 ;
        RECT 1334.070 25.880 1334.390 25.940 ;
      LAYER via ;
        RECT 686.420 25.880 686.680 26.140 ;
        RECT 1334.100 25.880 1334.360 26.140 ;
      LAYER met2 ;
        RECT 1335.010 1700.410 1335.290 1704.000 ;
        RECT 1334.160 1700.270 1335.290 1700.410 ;
        RECT 1334.160 26.170 1334.300 1700.270 ;
        RECT 1335.010 1700.000 1335.290 1700.270 ;
        RECT 686.420 25.850 686.680 26.170 ;
        RECT 1334.100 25.850 1334.360 26.170 ;
        RECT 686.480 2.400 686.620 25.850 ;
        RECT 686.270 -4.800 686.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1346.490 26.080 1346.810 26.140 ;
        RECT 1512.090 26.080 1512.410 26.140 ;
        RECT 1346.490 25.940 1512.410 26.080 ;
        RECT 1346.490 25.880 1346.810 25.940 ;
        RECT 1512.090 25.880 1512.410 25.940 ;
      LAYER via ;
        RECT 1346.520 25.880 1346.780 26.140 ;
        RECT 1512.120 25.880 1512.380 26.140 ;
      LAYER met2 ;
        RECT 1513.490 1700.410 1513.770 1704.000 ;
        RECT 1512.180 1700.270 1513.770 1700.410 ;
        RECT 1512.180 26.170 1512.320 1700.270 ;
        RECT 1513.490 1700.000 1513.770 1700.270 ;
        RECT 1346.520 25.850 1346.780 26.170 ;
        RECT 1512.120 25.850 1512.380 26.170 ;
        RECT 1346.580 2.400 1346.720 25.850 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 0.300 ;
=======
      LAYER li1 ;
        RECT 1486.865 1686.825 1487.035 1690.395 ;
      LAYER mcon ;
        RECT 1486.865 1690.225 1487.035 1690.395 ;
      LAYER met1 ;
        RECT 1369.490 1690.380 1369.810 1690.440 ;
        RECT 1486.805 1690.380 1487.095 1690.425 ;
        RECT 1369.490 1690.240 1487.095 1690.380 ;
        RECT 1369.490 1690.180 1369.810 1690.240 ;
        RECT 1486.805 1690.195 1487.095 1690.240 ;
        RECT 1486.805 1686.980 1487.095 1687.025 ;
        RECT 1518.070 1686.980 1518.390 1687.040 ;
        RECT 1486.805 1686.840 1518.390 1686.980 ;
        RECT 1486.805 1686.795 1487.095 1686.840 ;
        RECT 1518.070 1686.780 1518.390 1686.840 ;
        RECT 1364.430 16.900 1364.750 16.960 ;
        RECT 1369.490 16.900 1369.810 16.960 ;
        RECT 1364.430 16.760 1369.810 16.900 ;
        RECT 1364.430 16.700 1364.750 16.760 ;
        RECT 1369.490 16.700 1369.810 16.760 ;
      LAYER via ;
        RECT 1369.520 1690.180 1369.780 1690.440 ;
        RECT 1518.100 1686.780 1518.360 1687.040 ;
        RECT 1364.460 16.700 1364.720 16.960 ;
        RECT 1369.520 16.700 1369.780 16.960 ;
      LAYER met2 ;
        RECT 1518.090 1700.000 1518.370 1704.000 ;
        RECT 1369.520 1690.150 1369.780 1690.470 ;
        RECT 1369.580 16.990 1369.720 1690.150 ;
        RECT 1518.160 1687.070 1518.300 1700.000 ;
        RECT 1518.100 1686.750 1518.360 1687.070 ;
        RECT 1364.460 16.670 1364.720 16.990 ;
        RECT 1369.520 16.670 1369.780 16.990 ;
        RECT 1364.520 2.400 1364.660 16.670 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 0.300 ;
=======
      LAYER li1 ;
        RECT 1438.565 1684.785 1438.735 1686.655 ;
      LAYER mcon ;
        RECT 1438.565 1686.485 1438.735 1686.655 ;
      LAYER met1 ;
        RECT 1438.505 1686.640 1438.795 1686.685 ;
        RECT 1438.505 1686.500 1487.020 1686.640 ;
        RECT 1438.505 1686.455 1438.795 1686.500 ;
        RECT 1486.880 1686.300 1487.020 1686.500 ;
        RECT 1523.130 1686.300 1523.450 1686.360 ;
        RECT 1486.880 1686.160 1523.450 1686.300 ;
        RECT 1523.130 1686.100 1523.450 1686.160 ;
        RECT 1390.650 1684.940 1390.970 1685.000 ;
        RECT 1438.505 1684.940 1438.795 1684.985 ;
        RECT 1390.650 1684.800 1438.795 1684.940 ;
        RECT 1390.650 1684.740 1390.970 1684.800 ;
        RECT 1438.505 1684.755 1438.795 1684.800 ;
        RECT 1382.370 20.640 1382.690 20.700 ;
        RECT 1390.190 20.640 1390.510 20.700 ;
        RECT 1382.370 20.500 1390.510 20.640 ;
        RECT 1382.370 20.440 1382.690 20.500 ;
        RECT 1390.190 20.440 1390.510 20.500 ;
      LAYER via ;
        RECT 1523.160 1686.100 1523.420 1686.360 ;
        RECT 1390.680 1684.740 1390.940 1685.000 ;
        RECT 1382.400 20.440 1382.660 20.700 ;
        RECT 1390.220 20.440 1390.480 20.700 ;
      LAYER met2 ;
        RECT 1523.150 1700.000 1523.430 1704.000 ;
        RECT 1523.220 1686.390 1523.360 1700.000 ;
        RECT 1523.160 1686.070 1523.420 1686.390 ;
        RECT 1390.680 1684.710 1390.940 1685.030 ;
        RECT 1390.740 1670.490 1390.880 1684.710 ;
        RECT 1390.280 1670.350 1390.880 1670.490 ;
        RECT 1390.280 20.730 1390.420 1670.350 ;
        RECT 1382.400 20.410 1382.660 20.730 ;
        RECT 1390.220 20.410 1390.480 20.730 ;
        RECT 1382.460 2.400 1382.600 20.410 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 0.300 ;
=======
      LAYER li1 ;
        RECT 1459.265 16.065 1462.655 16.235 ;
        RECT 1465.245 16.065 1465.415 17.935 ;
        RECT 1508.025 17.765 1508.195 19.635 ;
        RECT 1437.645 14.535 1437.815 15.555 ;
        RECT 1437.645 14.365 1439.655 14.535 ;
        RECT 1459.265 14.365 1459.435 16.065 ;
      LAYER mcon ;
        RECT 1508.025 19.465 1508.195 19.635 ;
        RECT 1465.245 17.765 1465.415 17.935 ;
        RECT 1462.485 16.065 1462.655 16.235 ;
        RECT 1437.645 15.385 1437.815 15.555 ;
        RECT 1439.485 14.365 1439.655 14.535 ;
      LAYER met1 ;
        RECT 1526.810 19.960 1527.130 20.020 ;
        RECT 1518.620 19.820 1527.130 19.960 ;
        RECT 1507.965 19.620 1508.255 19.665 ;
        RECT 1518.620 19.620 1518.760 19.820 ;
        RECT 1526.810 19.760 1527.130 19.820 ;
        RECT 1507.965 19.480 1518.760 19.620 ;
        RECT 1507.965 19.435 1508.255 19.480 ;
        RECT 1465.185 17.920 1465.475 17.965 ;
        RECT 1507.965 17.920 1508.255 17.965 ;
        RECT 1465.185 17.780 1508.255 17.920 ;
        RECT 1465.185 17.735 1465.475 17.780 ;
        RECT 1507.965 17.735 1508.255 17.780 ;
        RECT 1462.425 16.220 1462.715 16.265 ;
        RECT 1465.185 16.220 1465.475 16.265 ;
        RECT 1462.425 16.080 1465.475 16.220 ;
        RECT 1462.425 16.035 1462.715 16.080 ;
        RECT 1465.185 16.035 1465.475 16.080 ;
        RECT 1400.310 15.540 1400.630 15.600 ;
        RECT 1437.585 15.540 1437.875 15.585 ;
        RECT 1400.310 15.400 1437.875 15.540 ;
        RECT 1400.310 15.340 1400.630 15.400 ;
        RECT 1437.585 15.355 1437.875 15.400 ;
        RECT 1439.425 14.520 1439.715 14.565 ;
        RECT 1459.205 14.520 1459.495 14.565 ;
        RECT 1439.425 14.380 1459.495 14.520 ;
        RECT 1439.425 14.335 1439.715 14.380 ;
        RECT 1459.205 14.335 1459.495 14.380 ;
      LAYER via ;
        RECT 1526.840 19.760 1527.100 20.020 ;
        RECT 1400.340 15.340 1400.600 15.600 ;
      LAYER met2 ;
        RECT 1527.750 1700.410 1528.030 1704.000 ;
        RECT 1526.900 1700.270 1528.030 1700.410 ;
        RECT 1526.900 20.050 1527.040 1700.270 ;
        RECT 1527.750 1700.000 1528.030 1700.270 ;
        RECT 1526.840 19.730 1527.100 20.050 ;
        RECT 1400.340 15.310 1400.600 15.630 ;
        RECT 1400.400 2.400 1400.540 15.310 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1424.690 1685.960 1425.010 1686.020 ;
        RECT 1532.790 1685.960 1533.110 1686.020 ;
        RECT 1424.690 1685.820 1533.110 1685.960 ;
        RECT 1424.690 1685.760 1425.010 1685.820 ;
        RECT 1532.790 1685.760 1533.110 1685.820 ;
        RECT 1418.250 16.560 1418.570 16.620 ;
        RECT 1424.690 16.560 1425.010 16.620 ;
        RECT 1418.250 16.420 1425.010 16.560 ;
        RECT 1418.250 16.360 1418.570 16.420 ;
        RECT 1424.690 16.360 1425.010 16.420 ;
      LAYER via ;
        RECT 1424.720 1685.760 1424.980 1686.020 ;
        RECT 1532.820 1685.760 1533.080 1686.020 ;
        RECT 1418.280 16.360 1418.540 16.620 ;
        RECT 1424.720 16.360 1424.980 16.620 ;
      LAYER met2 ;
        RECT 1532.810 1700.000 1533.090 1704.000 ;
        RECT 1532.880 1686.050 1533.020 1700.000 ;
        RECT 1424.720 1685.730 1424.980 1686.050 ;
        RECT 1532.820 1685.730 1533.080 1686.050 ;
        RECT 1424.780 16.650 1424.920 1685.730 ;
        RECT 1418.280 16.330 1418.540 16.650 ;
        RECT 1424.720 16.330 1424.980 16.650 ;
        RECT 1418.340 2.400 1418.480 16.330 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1487.250 1686.640 1487.570 1686.700 ;
        RECT 1537.390 1686.640 1537.710 1686.700 ;
        RECT 1487.250 1686.500 1537.710 1686.640 ;
        RECT 1487.250 1686.440 1487.570 1686.500 ;
        RECT 1537.390 1686.440 1537.710 1686.500 ;
        RECT 1483.570 18.940 1483.890 19.000 ;
        RECT 1464.340 18.800 1483.890 18.940 ;
        RECT 1436.650 18.260 1436.970 18.320 ;
        RECT 1464.340 18.260 1464.480 18.800 ;
        RECT 1483.570 18.740 1483.890 18.800 ;
        RECT 1436.650 18.120 1464.480 18.260 ;
        RECT 1483.570 18.260 1483.890 18.320 ;
        RECT 1486.790 18.260 1487.110 18.320 ;
        RECT 1483.570 18.120 1487.110 18.260 ;
        RECT 1436.650 18.060 1436.970 18.120 ;
        RECT 1483.570 18.060 1483.890 18.120 ;
        RECT 1486.790 18.060 1487.110 18.120 ;
      LAYER via ;
        RECT 1487.280 1686.440 1487.540 1686.700 ;
        RECT 1537.420 1686.440 1537.680 1686.700 ;
        RECT 1436.680 18.060 1436.940 18.320 ;
        RECT 1483.600 18.740 1483.860 19.000 ;
        RECT 1483.600 18.060 1483.860 18.320 ;
        RECT 1486.820 18.060 1487.080 18.320 ;
      LAYER met2 ;
        RECT 1537.410 1700.000 1537.690 1704.000 ;
        RECT 1537.480 1686.730 1537.620 1700.000 ;
        RECT 1487.280 1686.410 1487.540 1686.730 ;
        RECT 1537.420 1686.410 1537.680 1686.730 ;
        RECT 1487.340 1671.170 1487.480 1686.410 ;
        RECT 1486.880 1671.030 1487.480 1671.170 ;
        RECT 1483.600 18.710 1483.860 19.030 ;
        RECT 1483.660 18.350 1483.800 18.710 ;
        RECT 1486.880 18.350 1487.020 1671.030 ;
        RECT 1436.680 18.030 1436.940 18.350 ;
        RECT 1483.600 18.030 1483.860 18.350 ;
        RECT 1486.820 18.030 1487.080 18.350 ;
        RECT 1436.740 9.250 1436.880 18.030 ;
        RECT 1435.820 9.110 1436.880 9.250 ;
        RECT 1435.820 2.400 1435.960 9.110 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1453.670 14.860 1453.990 14.920 ;
        RECT 1541.070 14.860 1541.390 14.920 ;
        RECT 1453.670 14.720 1541.390 14.860 ;
        RECT 1453.670 14.660 1453.990 14.720 ;
        RECT 1541.070 14.660 1541.390 14.720 ;
      LAYER via ;
        RECT 1453.700 14.660 1453.960 14.920 ;
        RECT 1541.100 14.660 1541.360 14.920 ;
      LAYER met2 ;
        RECT 1542.470 1700.410 1542.750 1704.000 ;
        RECT 1541.160 1700.270 1542.750 1700.410 ;
        RECT 1541.160 14.950 1541.300 1700.270 ;
        RECT 1542.470 1700.000 1542.750 1700.270 ;
        RECT 1453.700 14.630 1453.960 14.950 ;
        RECT 1541.100 14.630 1541.360 14.950 ;
        RECT 1453.760 2.400 1453.900 14.630 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1507.950 1687.320 1508.270 1687.380 ;
        RECT 1547.050 1687.320 1547.370 1687.380 ;
        RECT 1507.950 1687.180 1547.370 1687.320 ;
        RECT 1507.950 1687.120 1508.270 1687.180 ;
        RECT 1547.050 1687.120 1547.370 1687.180 ;
        RECT 1471.610 19.620 1471.930 19.680 ;
        RECT 1507.490 19.620 1507.810 19.680 ;
        RECT 1471.610 19.480 1507.810 19.620 ;
        RECT 1471.610 19.420 1471.930 19.480 ;
        RECT 1507.490 19.420 1507.810 19.480 ;
      LAYER via ;
        RECT 1507.980 1687.120 1508.240 1687.380 ;
        RECT 1547.080 1687.120 1547.340 1687.380 ;
        RECT 1471.640 19.420 1471.900 19.680 ;
        RECT 1507.520 19.420 1507.780 19.680 ;
      LAYER met2 ;
        RECT 1547.070 1700.000 1547.350 1704.000 ;
        RECT 1547.140 1687.410 1547.280 1700.000 ;
        RECT 1507.980 1687.090 1508.240 1687.410 ;
        RECT 1547.080 1687.090 1547.340 1687.410 ;
        RECT 1508.040 1671.850 1508.180 1687.090 ;
        RECT 1507.580 1671.710 1508.180 1671.850 ;
        RECT 1507.580 19.710 1507.720 1671.710 ;
        RECT 1471.640 19.390 1471.900 19.710 ;
        RECT 1507.520 19.390 1507.780 19.710 ;
        RECT 1471.700 2.400 1471.840 19.390 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1521.750 1684.260 1522.070 1684.320 ;
        RECT 1551.650 1684.260 1551.970 1684.320 ;
        RECT 1521.750 1684.120 1551.970 1684.260 ;
        RECT 1521.750 1684.060 1522.070 1684.120 ;
        RECT 1551.650 1684.060 1551.970 1684.120 ;
        RECT 1489.550 15.880 1489.870 15.940 ;
        RECT 1521.750 15.880 1522.070 15.940 ;
        RECT 1489.550 15.740 1522.070 15.880 ;
        RECT 1489.550 15.680 1489.870 15.740 ;
        RECT 1521.750 15.680 1522.070 15.740 ;
      LAYER via ;
        RECT 1521.780 1684.060 1522.040 1684.320 ;
        RECT 1551.680 1684.060 1551.940 1684.320 ;
        RECT 1489.580 15.680 1489.840 15.940 ;
        RECT 1521.780 15.680 1522.040 15.940 ;
      LAYER met2 ;
        RECT 1551.670 1700.000 1551.950 1704.000 ;
        RECT 1551.740 1684.350 1551.880 1700.000 ;
        RECT 1521.780 1684.030 1522.040 1684.350 ;
        RECT 1551.680 1684.030 1551.940 1684.350 ;
        RECT 1521.840 15.970 1521.980 1684.030 ;
        RECT 1489.580 15.650 1489.840 15.970 ;
        RECT 1521.780 15.650 1522.040 15.970 ;
        RECT 1489.640 2.400 1489.780 15.650 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 0.300 ;
=======
      LAYER met1 ;
        RECT 1528.190 1683.920 1528.510 1683.980 ;
        RECT 1556.710 1683.920 1557.030 1683.980 ;
        RECT 1528.190 1683.780 1557.030 1683.920 ;
        RECT 1528.190 1683.720 1528.510 1683.780 ;
        RECT 1556.710 1683.720 1557.030 1683.780 ;
        RECT 1507.030 18.600 1507.350 18.660 ;
        RECT 1528.190 18.600 1528.510 18.660 ;
        RECT 1507.030 18.460 1528.510 18.600 ;
        RECT 1507.030 18.400 1507.350 18.460 ;
        RECT 1528.190 18.400 1528.510 18.460 ;
      LAYER via ;
        RECT 1528.220 1683.720 1528.480 1683.980 ;
        RECT 1556.740 1683.720 1557.000 1683.980 ;
        RECT 1507.060 18.400 1507.320 18.660 ;
        RECT 1528.220 18.400 1528.480 18.660 ;
      LAYER met2 ;
        RECT 1556.730 1700.000 1557.010 1704.000 ;
        RECT 1556.800 1684.010 1556.940 1700.000 ;
        RECT 1528.220 1683.690 1528.480 1684.010 ;
        RECT 1556.740 1683.690 1557.000 1684.010 ;
        RECT 1528.280 18.690 1528.420 1683.690 ;
        RECT 1507.060 18.370 1507.320 18.690 ;
        RECT 1528.220 18.370 1528.480 18.690 ;
        RECT 1507.120 2.400 1507.260 18.370 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1340.050 1656.380 1340.370 1656.440 ;
        RECT 1339.680 1656.240 1340.370 1656.380 ;
        RECT 1339.680 1656.100 1339.820 1656.240 ;
        RECT 1340.050 1656.180 1340.370 1656.240 ;
        RECT 1339.590 1655.840 1339.910 1656.100 ;
        RECT 710.310 54.980 710.630 55.040 ;
        RECT 1339.590 54.980 1339.910 55.040 ;
        RECT 710.310 54.840 1339.910 54.980 ;
        RECT 710.310 54.780 710.630 54.840 ;
        RECT 1339.590 54.780 1339.910 54.840 ;
        RECT 704.330 20.980 704.650 21.040 ;
        RECT 710.310 20.980 710.630 21.040 ;
        RECT 704.330 20.840 710.630 20.980 ;
        RECT 704.330 20.780 704.650 20.840 ;
        RECT 710.310 20.780 710.630 20.840 ;
      LAYER via ;
        RECT 1340.080 1656.180 1340.340 1656.440 ;
        RECT 1339.620 1655.840 1339.880 1656.100 ;
        RECT 710.340 54.780 710.600 55.040 ;
        RECT 1339.620 54.780 1339.880 55.040 ;
        RECT 704.360 20.780 704.620 21.040 ;
        RECT 710.340 20.780 710.600 21.040 ;
      LAYER met2 ;
        RECT 1340.070 1700.000 1340.350 1704.000 ;
        RECT 1340.140 1656.470 1340.280 1700.000 ;
        RECT 1340.080 1656.150 1340.340 1656.470 ;
        RECT 1339.620 1655.810 1339.880 1656.130 ;
        RECT 1339.680 55.070 1339.820 1655.810 ;
        RECT 710.340 54.750 710.600 55.070 ;
        RECT 1339.620 54.750 1339.880 55.070 ;
        RECT 710.400 21.070 710.540 54.750 ;
        RECT 704.360 20.750 704.620 21.070 ;
        RECT 710.340 20.750 710.600 21.070 ;
        RECT 704.420 2.400 704.560 20.750 ;
        RECT 704.210 -4.800 704.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1541.990 1689.360 1542.310 1689.420 ;
        RECT 1561.310 1689.360 1561.630 1689.420 ;
        RECT 1541.990 1689.220 1561.630 1689.360 ;
        RECT 1541.990 1689.160 1542.310 1689.220 ;
        RECT 1561.310 1689.160 1561.630 1689.220 ;
        RECT 1524.970 15.880 1525.290 15.940 ;
        RECT 1541.990 15.880 1542.310 15.940 ;
        RECT 1524.970 15.740 1542.310 15.880 ;
        RECT 1524.970 15.680 1525.290 15.740 ;
        RECT 1541.990 15.680 1542.310 15.740 ;
      LAYER via ;
        RECT 1542.020 1689.160 1542.280 1689.420 ;
        RECT 1561.340 1689.160 1561.600 1689.420 ;
        RECT 1525.000 15.680 1525.260 15.940 ;
        RECT 1542.020 15.680 1542.280 15.940 ;
      LAYER met2 ;
        RECT 1561.330 1700.000 1561.610 1704.000 ;
        RECT 1561.400 1689.450 1561.540 1700.000 ;
        RECT 1542.020 1689.130 1542.280 1689.450 ;
        RECT 1561.340 1689.130 1561.600 1689.450 ;
        RECT 1542.080 15.970 1542.220 1689.130 ;
        RECT 1525.000 15.650 1525.260 15.970 ;
        RECT 1542.020 15.650 1542.280 15.970 ;
        RECT 1525.060 2.400 1525.200 15.650 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1545.210 1686.640 1545.530 1686.700 ;
        RECT 1566.370 1686.640 1566.690 1686.700 ;
        RECT 1545.210 1686.500 1566.690 1686.640 ;
        RECT 1545.210 1686.440 1545.530 1686.500 ;
        RECT 1566.370 1686.440 1566.690 1686.500 ;
        RECT 1542.910 20.640 1543.230 20.700 ;
        RECT 1545.210 20.640 1545.530 20.700 ;
        RECT 1542.910 20.500 1545.530 20.640 ;
        RECT 1542.910 20.440 1543.230 20.500 ;
        RECT 1545.210 20.440 1545.530 20.500 ;
      LAYER via ;
        RECT 1545.240 1686.440 1545.500 1686.700 ;
        RECT 1566.400 1686.440 1566.660 1686.700 ;
        RECT 1542.940 20.440 1543.200 20.700 ;
        RECT 1545.240 20.440 1545.500 20.700 ;
      LAYER met2 ;
        RECT 1566.390 1700.000 1566.670 1704.000 ;
        RECT 1566.460 1686.730 1566.600 1700.000 ;
        RECT 1545.240 1686.410 1545.500 1686.730 ;
        RECT 1566.400 1686.410 1566.660 1686.730 ;
        RECT 1545.300 20.730 1545.440 1686.410 ;
        RECT 1542.940 20.410 1543.200 20.730 ;
        RECT 1545.240 20.410 1545.500 20.730 ;
        RECT 1543.000 2.400 1543.140 20.410 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1565.910 1683.920 1566.230 1683.980 ;
        RECT 1570.970 1683.920 1571.290 1683.980 ;
        RECT 1565.910 1683.780 1571.290 1683.920 ;
        RECT 1565.910 1683.720 1566.230 1683.780 ;
        RECT 1570.970 1683.720 1571.290 1683.780 ;
        RECT 1560.850 20.640 1561.170 20.700 ;
        RECT 1565.910 20.640 1566.230 20.700 ;
        RECT 1560.850 20.500 1566.230 20.640 ;
        RECT 1560.850 20.440 1561.170 20.500 ;
        RECT 1565.910 20.440 1566.230 20.500 ;
      LAYER via ;
        RECT 1565.940 1683.720 1566.200 1683.980 ;
        RECT 1571.000 1683.720 1571.260 1683.980 ;
        RECT 1560.880 20.440 1561.140 20.700 ;
        RECT 1565.940 20.440 1566.200 20.700 ;
      LAYER met2 ;
        RECT 1570.990 1700.000 1571.270 1704.000 ;
        RECT 1571.060 1684.010 1571.200 1700.000 ;
        RECT 1565.940 1683.690 1566.200 1684.010 ;
        RECT 1571.000 1683.690 1571.260 1684.010 ;
        RECT 1566.000 20.730 1566.140 1683.690 ;
        RECT 1560.880 20.410 1561.140 20.730 ;
        RECT 1565.940 20.410 1566.200 20.730 ;
        RECT 1560.940 2.400 1561.080 20.410 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 0.300 ;
=======
      LAYER met1 ;
        RECT 1575.110 20.640 1575.430 20.700 ;
        RECT 1578.790 20.640 1579.110 20.700 ;
        RECT 1575.110 20.500 1579.110 20.640 ;
        RECT 1575.110 20.440 1575.430 20.500 ;
        RECT 1578.790 20.440 1579.110 20.500 ;
      LAYER via ;
        RECT 1575.140 20.440 1575.400 20.700 ;
        RECT 1578.820 20.440 1579.080 20.700 ;
      LAYER met2 ;
        RECT 1576.050 1700.410 1576.330 1704.000 ;
        RECT 1575.200 1700.270 1576.330 1700.410 ;
        RECT 1575.200 20.730 1575.340 1700.270 ;
        RECT 1576.050 1700.000 1576.330 1700.270 ;
        RECT 1575.140 20.410 1575.400 20.730 ;
        RECT 1578.820 20.410 1579.080 20.730 ;
        RECT 1578.880 2.400 1579.020 20.410 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 0.300 ;
=======
      LAYER met1 ;
        RECT 1580.630 1684.600 1580.950 1684.660 ;
        RECT 1594.430 1684.600 1594.750 1684.660 ;
        RECT 1580.630 1684.460 1594.750 1684.600 ;
        RECT 1580.630 1684.400 1580.950 1684.460 ;
        RECT 1594.430 1684.400 1594.750 1684.460 ;
        RECT 1594.430 2.960 1594.750 3.020 ;
        RECT 1596.270 2.960 1596.590 3.020 ;
        RECT 1594.430 2.820 1596.590 2.960 ;
        RECT 1594.430 2.760 1594.750 2.820 ;
        RECT 1596.270 2.760 1596.590 2.820 ;
      LAYER via ;
        RECT 1580.660 1684.400 1580.920 1684.660 ;
        RECT 1594.460 1684.400 1594.720 1684.660 ;
        RECT 1594.460 2.760 1594.720 3.020 ;
        RECT 1596.300 2.760 1596.560 3.020 ;
      LAYER met2 ;
        RECT 1580.650 1700.000 1580.930 1704.000 ;
        RECT 1580.720 1684.690 1580.860 1700.000 ;
        RECT 1580.660 1684.370 1580.920 1684.690 ;
        RECT 1594.460 1684.370 1594.720 1684.690 ;
        RECT 1594.520 3.050 1594.660 1684.370 ;
        RECT 1594.460 2.730 1594.720 3.050 ;
        RECT 1596.300 2.730 1596.560 3.050 ;
        RECT 1596.360 2.400 1596.500 2.730 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1586.150 16.220 1586.470 16.280 ;
        RECT 1614.210 16.220 1614.530 16.280 ;
        RECT 1586.150 16.080 1614.530 16.220 ;
        RECT 1586.150 16.020 1586.470 16.080 ;
        RECT 1614.210 16.020 1614.530 16.080 ;
      LAYER via ;
        RECT 1586.180 16.020 1586.440 16.280 ;
        RECT 1614.240 16.020 1614.500 16.280 ;
      LAYER met2 ;
        RECT 1585.710 1700.410 1585.990 1704.000 ;
        RECT 1585.710 1700.270 1586.380 1700.410 ;
        RECT 1585.710 1700.000 1585.990 1700.270 ;
        RECT 1586.240 16.310 1586.380 1700.270 ;
        RECT 1586.180 15.990 1586.440 16.310 ;
        RECT 1614.240 15.990 1614.500 16.310 ;
        RECT 1614.300 2.400 1614.440 15.990 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1590.290 1684.260 1590.610 1684.320 ;
        RECT 1597.190 1684.260 1597.510 1684.320 ;
        RECT 1590.290 1684.120 1597.510 1684.260 ;
        RECT 1590.290 1684.060 1590.610 1684.120 ;
        RECT 1597.190 1684.060 1597.510 1684.120 ;
        RECT 1632.150 16.220 1632.470 16.280 ;
        RECT 1614.760 16.080 1632.470 16.220 ;
        RECT 1597.190 15.880 1597.510 15.940 ;
        RECT 1614.760 15.880 1614.900 16.080 ;
        RECT 1632.150 16.020 1632.470 16.080 ;
        RECT 1597.190 15.740 1614.900 15.880 ;
        RECT 1597.190 15.680 1597.510 15.740 ;
      LAYER via ;
        RECT 1590.320 1684.060 1590.580 1684.320 ;
        RECT 1597.220 1684.060 1597.480 1684.320 ;
        RECT 1597.220 15.680 1597.480 15.940 ;
        RECT 1632.180 16.020 1632.440 16.280 ;
      LAYER met2 ;
        RECT 1590.310 1700.000 1590.590 1704.000 ;
        RECT 1590.380 1684.350 1590.520 1700.000 ;
        RECT 1590.320 1684.030 1590.580 1684.350 ;
        RECT 1597.220 1684.030 1597.480 1684.350 ;
        RECT 1597.280 15.970 1597.420 1684.030 ;
        RECT 1632.180 15.990 1632.440 16.310 ;
        RECT 1597.220 15.650 1597.480 15.970 ;
        RECT 1632.240 2.400 1632.380 15.990 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1595.350 1684.600 1595.670 1684.660 ;
        RECT 1604.550 1684.600 1604.870 1684.660 ;
        RECT 1595.350 1684.460 1604.870 1684.600 ;
        RECT 1595.350 1684.400 1595.670 1684.460 ;
        RECT 1604.550 1684.400 1604.870 1684.460 ;
        RECT 1604.550 17.580 1604.870 17.640 ;
        RECT 1604.550 17.440 1608.920 17.580 ;
        RECT 1604.550 17.380 1604.870 17.440 ;
        RECT 1608.780 17.240 1608.920 17.440 ;
        RECT 1650.090 17.240 1650.410 17.300 ;
        RECT 1608.780 17.100 1650.410 17.240 ;
        RECT 1650.090 17.040 1650.410 17.100 ;
      LAYER via ;
        RECT 1595.380 1684.400 1595.640 1684.660 ;
        RECT 1604.580 1684.400 1604.840 1684.660 ;
        RECT 1604.580 17.380 1604.840 17.640 ;
        RECT 1650.120 17.040 1650.380 17.300 ;
      LAYER met2 ;
        RECT 1595.370 1700.000 1595.650 1704.000 ;
        RECT 1595.440 1684.690 1595.580 1700.000 ;
        RECT 1595.380 1684.370 1595.640 1684.690 ;
        RECT 1604.580 1684.370 1604.840 1684.690 ;
        RECT 1604.640 17.670 1604.780 1684.370 ;
        RECT 1604.580 17.350 1604.840 17.670 ;
        RECT 1650.120 17.010 1650.380 17.330 ;
        RECT 1650.180 2.400 1650.320 17.010 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 0.300 ;
=======
      LAYER met1 ;
        RECT 1599.950 20.640 1600.270 20.700 ;
        RECT 1668.030 20.640 1668.350 20.700 ;
        RECT 1599.950 20.500 1668.350 20.640 ;
        RECT 1599.950 20.440 1600.270 20.500 ;
        RECT 1668.030 20.440 1668.350 20.500 ;
      LAYER via ;
        RECT 1599.980 20.440 1600.240 20.700 ;
        RECT 1668.060 20.440 1668.320 20.700 ;
      LAYER met2 ;
        RECT 1599.970 1700.000 1600.250 1704.000 ;
        RECT 1600.040 20.730 1600.180 1700.000 ;
        RECT 1599.980 20.410 1600.240 20.730 ;
        RECT 1668.060 20.410 1668.320 20.730 ;
        RECT 1668.120 2.400 1668.260 20.410 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 0.300 ;
=======
      LAYER li1 ;
        RECT 1674.085 17.425 1674.255 20.315 ;
      LAYER mcon ;
        RECT 1674.085 20.145 1674.255 20.315 ;
      LAYER met1 ;
        RECT 1605.010 1683.920 1605.330 1683.980 ;
        RECT 1606.850 1683.920 1607.170 1683.980 ;
        RECT 1605.010 1683.780 1607.170 1683.920 ;
        RECT 1605.010 1683.720 1605.330 1683.780 ;
        RECT 1606.850 1683.720 1607.170 1683.780 ;
        RECT 1606.850 20.300 1607.170 20.360 ;
        RECT 1674.025 20.300 1674.315 20.345 ;
        RECT 1606.850 20.160 1674.315 20.300 ;
        RECT 1606.850 20.100 1607.170 20.160 ;
        RECT 1674.025 20.115 1674.315 20.160 ;
        RECT 1674.025 17.580 1674.315 17.625 ;
        RECT 1685.510 17.580 1685.830 17.640 ;
        RECT 1674.025 17.440 1685.830 17.580 ;
        RECT 1674.025 17.395 1674.315 17.440 ;
        RECT 1685.510 17.380 1685.830 17.440 ;
      LAYER via ;
        RECT 1605.040 1683.720 1605.300 1683.980 ;
        RECT 1606.880 1683.720 1607.140 1683.980 ;
        RECT 1606.880 20.100 1607.140 20.360 ;
        RECT 1685.540 17.380 1685.800 17.640 ;
      LAYER met2 ;
        RECT 1605.030 1700.000 1605.310 1704.000 ;
        RECT 1605.100 1684.010 1605.240 1700.000 ;
        RECT 1605.040 1683.690 1605.300 1684.010 ;
        RECT 1606.880 1683.690 1607.140 1684.010 ;
        RECT 1606.940 20.390 1607.080 1683.690 ;
        RECT 1606.880 20.070 1607.140 20.390 ;
        RECT 1685.540 17.350 1685.800 17.670 ;
        RECT 1685.600 2.400 1685.740 17.350 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 0.300 ;
=======
      LAYER li1 ;
        RECT 1340.585 1580.065 1340.755 1594.515 ;
        RECT 1340.585 1435.225 1340.755 1442.195 ;
        RECT 1340.585 565.845 1340.755 613.275 ;
        RECT 1341.045 421.345 1341.215 475.915 ;
        RECT 1341.045 324.785 1341.215 372.555 ;
        RECT 1341.045 276.165 1341.215 324.275 ;
      LAYER mcon ;
        RECT 1340.585 1594.345 1340.755 1594.515 ;
        RECT 1340.585 1442.025 1340.755 1442.195 ;
        RECT 1340.585 613.105 1340.755 613.275 ;
        RECT 1341.045 475.745 1341.215 475.915 ;
        RECT 1341.045 372.385 1341.215 372.555 ;
        RECT 1341.045 324.105 1341.215 324.275 ;
      LAYER met1 ;
        RECT 1341.430 1666.580 1341.750 1666.640 ;
        RECT 1344.190 1666.580 1344.510 1666.640 ;
        RECT 1341.430 1666.440 1344.510 1666.580 ;
        RECT 1341.430 1666.380 1341.750 1666.440 ;
        RECT 1344.190 1666.380 1344.510 1666.440 ;
        RECT 1340.525 1594.500 1340.815 1594.545 ;
        RECT 1341.430 1594.500 1341.750 1594.560 ;
        RECT 1340.525 1594.360 1341.750 1594.500 ;
        RECT 1340.525 1594.315 1340.815 1594.360 ;
        RECT 1341.430 1594.300 1341.750 1594.360 ;
        RECT 1340.510 1580.220 1340.830 1580.280 ;
        RECT 1340.315 1580.080 1340.830 1580.220 ;
        RECT 1340.510 1580.020 1340.830 1580.080 ;
        RECT 1340.525 1442.180 1340.815 1442.225 ;
        RECT 1340.970 1442.180 1341.290 1442.240 ;
        RECT 1340.525 1442.040 1341.290 1442.180 ;
        RECT 1340.525 1441.995 1340.815 1442.040 ;
        RECT 1340.970 1441.980 1341.290 1442.040 ;
        RECT 1340.510 1435.380 1340.830 1435.440 ;
        RECT 1340.315 1435.240 1340.830 1435.380 ;
        RECT 1340.510 1435.180 1340.830 1435.240 ;
        RECT 1340.510 1076.480 1340.830 1076.740 ;
        RECT 1340.600 1076.340 1340.740 1076.480 ;
        RECT 1340.970 1076.340 1341.290 1076.400 ;
        RECT 1340.600 1076.200 1341.290 1076.340 ;
        RECT 1340.970 1076.140 1341.290 1076.200 ;
        RECT 1340.510 917.900 1340.830 917.960 ;
        RECT 1341.430 917.900 1341.750 917.960 ;
        RECT 1340.510 917.760 1341.750 917.900 ;
        RECT 1340.510 917.700 1340.830 917.760 ;
        RECT 1341.430 917.700 1341.750 917.760 ;
        RECT 1340.510 613.740 1340.830 614.000 ;
        RECT 1340.600 613.305 1340.740 613.740 ;
        RECT 1340.525 613.075 1340.815 613.305 ;
        RECT 1340.510 566.000 1340.830 566.060 ;
        RECT 1340.315 565.860 1340.830 566.000 ;
        RECT 1340.510 565.800 1340.830 565.860 ;
        RECT 1340.970 475.900 1341.290 475.960 ;
        RECT 1340.775 475.760 1341.290 475.900 ;
        RECT 1340.970 475.700 1341.290 475.760 ;
        RECT 1340.510 421.500 1340.830 421.560 ;
        RECT 1340.985 421.500 1341.275 421.545 ;
        RECT 1340.510 421.360 1341.275 421.500 ;
        RECT 1340.510 421.300 1340.830 421.360 ;
        RECT 1340.985 421.315 1341.275 421.360 ;
        RECT 1340.510 420.820 1340.830 420.880 ;
        RECT 1341.430 420.820 1341.750 420.880 ;
        RECT 1340.510 420.680 1341.750 420.820 ;
        RECT 1340.510 420.620 1340.830 420.680 ;
        RECT 1341.430 420.620 1341.750 420.680 ;
        RECT 1340.970 372.540 1341.290 372.600 ;
        RECT 1340.775 372.400 1341.290 372.540 ;
        RECT 1340.970 372.340 1341.290 372.400 ;
        RECT 1340.970 324.940 1341.290 325.000 ;
        RECT 1340.775 324.800 1341.290 324.940 ;
        RECT 1340.970 324.740 1341.290 324.800 ;
        RECT 1340.970 324.260 1341.290 324.320 ;
        RECT 1340.775 324.120 1341.290 324.260 ;
        RECT 1340.970 324.060 1341.290 324.120 ;
        RECT 1340.985 276.320 1341.275 276.365 ;
        RECT 1341.430 276.320 1341.750 276.380 ;
        RECT 1340.985 276.180 1341.750 276.320 ;
        RECT 1340.985 276.135 1341.275 276.180 ;
        RECT 1341.430 276.120 1341.750 276.180 ;
        RECT 1340.970 234.840 1341.290 234.900 ;
        RECT 1340.600 234.700 1341.290 234.840 ;
        RECT 1340.600 234.220 1340.740 234.700 ;
        RECT 1340.970 234.640 1341.290 234.700 ;
        RECT 1340.510 233.960 1340.830 234.220 ;
        RECT 724.110 51.240 724.430 51.300 ;
        RECT 1340.510 51.240 1340.830 51.300 ;
        RECT 724.110 51.100 1340.830 51.240 ;
        RECT 724.110 51.040 724.430 51.100 ;
        RECT 1340.510 51.040 1340.830 51.100 ;
      LAYER via ;
        RECT 1341.460 1666.380 1341.720 1666.640 ;
        RECT 1344.220 1666.380 1344.480 1666.640 ;
        RECT 1341.460 1594.300 1341.720 1594.560 ;
        RECT 1340.540 1580.020 1340.800 1580.280 ;
        RECT 1341.000 1441.980 1341.260 1442.240 ;
        RECT 1340.540 1435.180 1340.800 1435.440 ;
        RECT 1340.540 1076.480 1340.800 1076.740 ;
        RECT 1341.000 1076.140 1341.260 1076.400 ;
        RECT 1340.540 917.700 1340.800 917.960 ;
        RECT 1341.460 917.700 1341.720 917.960 ;
        RECT 1340.540 613.740 1340.800 614.000 ;
        RECT 1340.540 565.800 1340.800 566.060 ;
        RECT 1341.000 475.700 1341.260 475.960 ;
        RECT 1340.540 421.300 1340.800 421.560 ;
        RECT 1340.540 420.620 1340.800 420.880 ;
        RECT 1341.460 420.620 1341.720 420.880 ;
        RECT 1341.000 372.340 1341.260 372.600 ;
        RECT 1341.000 324.740 1341.260 325.000 ;
        RECT 1341.000 324.060 1341.260 324.320 ;
        RECT 1341.460 276.120 1341.720 276.380 ;
        RECT 1341.000 234.640 1341.260 234.900 ;
        RECT 1340.540 233.960 1340.800 234.220 ;
        RECT 724.140 51.040 724.400 51.300 ;
        RECT 1340.540 51.040 1340.800 51.300 ;
      LAYER met2 ;
        RECT 1344.670 1700.410 1344.950 1704.000 ;
        RECT 1344.280 1700.270 1344.950 1700.410 ;
        RECT 1344.280 1666.670 1344.420 1700.270 ;
        RECT 1344.670 1700.000 1344.950 1700.270 ;
        RECT 1341.460 1666.350 1341.720 1666.670 ;
        RECT 1344.220 1666.350 1344.480 1666.670 ;
        RECT 1341.520 1594.590 1341.660 1666.350 ;
        RECT 1341.460 1594.270 1341.720 1594.590 ;
        RECT 1340.540 1580.165 1340.800 1580.310 ;
        RECT 1340.530 1579.795 1340.810 1580.165 ;
        RECT 1340.990 1537.635 1341.270 1538.005 ;
        RECT 1341.060 1442.270 1341.200 1537.635 ;
        RECT 1341.000 1441.950 1341.260 1442.270 ;
        RECT 1340.540 1435.150 1340.800 1435.470 ;
        RECT 1340.600 1076.770 1340.740 1435.150 ;
        RECT 1340.540 1076.450 1340.800 1076.770 ;
        RECT 1341.000 1076.110 1341.260 1076.430 ;
        RECT 1341.060 983.010 1341.200 1076.110 ;
        RECT 1341.060 982.870 1341.660 983.010 ;
        RECT 1341.520 917.990 1341.660 982.870 ;
        RECT 1340.540 917.670 1340.800 917.990 ;
        RECT 1341.460 917.670 1341.720 917.990 ;
        RECT 1340.600 821.965 1340.740 917.670 ;
        RECT 1340.530 821.595 1340.810 821.965 ;
        RECT 1340.530 820.915 1340.810 821.285 ;
        RECT 1340.600 719.285 1340.740 820.915 ;
        RECT 1340.530 718.915 1340.810 719.285 ;
        RECT 1340.530 717.555 1340.810 717.925 ;
        RECT 1340.600 614.030 1340.740 717.555 ;
        RECT 1340.540 613.710 1340.800 614.030 ;
        RECT 1340.540 565.770 1340.800 566.090 ;
        RECT 1340.600 549.170 1340.740 565.770 ;
        RECT 1340.600 549.030 1341.200 549.170 ;
        RECT 1341.060 475.990 1341.200 549.030 ;
        RECT 1341.000 475.670 1341.260 475.990 ;
        RECT 1340.540 421.270 1340.800 421.590 ;
        RECT 1340.600 420.910 1340.740 421.270 ;
        RECT 1340.540 420.590 1340.800 420.910 ;
        RECT 1341.460 420.590 1341.720 420.910 ;
        RECT 1341.520 373.050 1341.660 420.590 ;
        RECT 1341.060 372.910 1341.660 373.050 ;
        RECT 1341.060 372.630 1341.200 372.910 ;
        RECT 1341.000 372.310 1341.260 372.630 ;
        RECT 1341.000 324.710 1341.260 325.030 ;
        RECT 1341.060 324.350 1341.200 324.710 ;
        RECT 1341.000 324.030 1341.260 324.350 ;
        RECT 1341.460 276.090 1341.720 276.410 ;
        RECT 1341.520 275.810 1341.660 276.090 ;
        RECT 1341.060 275.670 1341.660 275.810 ;
        RECT 1341.060 234.930 1341.200 275.670 ;
        RECT 1341.000 234.610 1341.260 234.930 ;
        RECT 1340.540 233.930 1340.800 234.250 ;
        RECT 1340.600 51.330 1340.740 233.930 ;
        RECT 724.140 51.010 724.400 51.330 ;
        RECT 1340.540 51.010 1340.800 51.330 ;
        RECT 724.200 3.130 724.340 51.010 ;
        RECT 722.360 2.990 724.340 3.130 ;
        RECT 722.360 2.400 722.500 2.990 ;
        RECT 722.150 -4.800 722.710 2.400 ;
      LAYER via2 ;
        RECT 1340.530 1579.840 1340.810 1580.120 ;
        RECT 1340.990 1537.680 1341.270 1537.960 ;
        RECT 1340.530 821.640 1340.810 821.920 ;
        RECT 1340.530 820.960 1340.810 821.240 ;
        RECT 1340.530 718.960 1340.810 719.240 ;
        RECT 1340.530 717.600 1340.810 717.880 ;
      LAYER met3 ;
        RECT 1340.505 1580.140 1340.835 1580.145 ;
        RECT 1340.505 1580.130 1341.090 1580.140 ;
        RECT 1340.505 1579.830 1341.290 1580.130 ;
        RECT 1340.505 1579.820 1341.090 1579.830 ;
        RECT 1340.505 1579.815 1340.835 1579.820 ;
        RECT 1340.965 1537.980 1341.295 1537.985 ;
        RECT 1340.710 1537.970 1341.295 1537.980 ;
        RECT 1340.510 1537.670 1341.295 1537.970 ;
        RECT 1340.710 1537.660 1341.295 1537.670 ;
        RECT 1340.965 1537.655 1341.295 1537.660 ;
        RECT 1340.505 821.930 1340.835 821.945 ;
        RECT 1340.505 821.615 1341.050 821.930 ;
        RECT 1340.750 821.265 1341.050 821.615 ;
        RECT 1340.505 820.950 1341.050 821.265 ;
        RECT 1340.505 820.935 1340.835 820.950 ;
        RECT 1340.505 719.250 1340.835 719.265 ;
        RECT 1340.505 718.935 1341.050 719.250 ;
        RECT 1340.750 717.905 1341.050 718.935 ;
        RECT 1340.505 717.590 1341.050 717.905 ;
        RECT 1340.505 717.575 1340.835 717.590 ;
      LAYER via3 ;
        RECT 1340.740 1579.820 1341.060 1580.140 ;
        RECT 1340.740 1537.660 1341.060 1537.980 ;
      LAYER met4 ;
        RECT 1340.735 1579.815 1341.065 1580.145 ;
        RECT 1340.750 1537.985 1341.050 1579.815 ;
        RECT 1340.735 1537.655 1341.065 1537.985 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 0.300 ;
=======
      LAYER met1 ;
        RECT 1609.610 1686.300 1609.930 1686.360 ;
        RECT 1613.750 1686.300 1614.070 1686.360 ;
        RECT 1609.610 1686.160 1614.070 1686.300 ;
        RECT 1609.610 1686.100 1609.930 1686.160 ;
        RECT 1613.750 1686.100 1614.070 1686.160 ;
        RECT 1613.750 18.940 1614.070 19.000 ;
        RECT 1703.450 18.940 1703.770 19.000 ;
        RECT 1613.750 18.800 1703.770 18.940 ;
        RECT 1613.750 18.740 1614.070 18.800 ;
        RECT 1703.450 18.740 1703.770 18.800 ;
      LAYER via ;
        RECT 1609.640 1686.100 1609.900 1686.360 ;
        RECT 1613.780 1686.100 1614.040 1686.360 ;
        RECT 1613.780 18.740 1614.040 19.000 ;
        RECT 1703.480 18.740 1703.740 19.000 ;
      LAYER met2 ;
        RECT 1609.630 1700.000 1609.910 1704.000 ;
        RECT 1609.700 1686.390 1609.840 1700.000 ;
        RECT 1609.640 1686.070 1609.900 1686.390 ;
        RECT 1613.780 1686.070 1614.040 1686.390 ;
        RECT 1613.840 19.030 1613.980 1686.070 ;
        RECT 1613.780 18.710 1614.040 19.030 ;
        RECT 1703.480 18.710 1703.740 19.030 ;
        RECT 1703.540 2.400 1703.680 18.710 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 0.300 ;
=======
      LAYER met1 ;
        RECT 1614.670 1688.340 1614.990 1688.400 ;
        RECT 1620.650 1688.340 1620.970 1688.400 ;
        RECT 1614.670 1688.200 1620.970 1688.340 ;
        RECT 1614.670 1688.140 1614.990 1688.200 ;
        RECT 1620.650 1688.140 1620.970 1688.200 ;
        RECT 1620.650 14.180 1620.970 14.240 ;
        RECT 1721.390 14.180 1721.710 14.240 ;
        RECT 1620.650 14.040 1721.710 14.180 ;
        RECT 1620.650 13.980 1620.970 14.040 ;
        RECT 1721.390 13.980 1721.710 14.040 ;
      LAYER via ;
        RECT 1614.700 1688.140 1614.960 1688.400 ;
        RECT 1620.680 1688.140 1620.940 1688.400 ;
        RECT 1620.680 13.980 1620.940 14.240 ;
        RECT 1721.420 13.980 1721.680 14.240 ;
      LAYER met2 ;
        RECT 1614.690 1700.000 1614.970 1704.000 ;
        RECT 1614.760 1688.430 1614.900 1700.000 ;
        RECT 1614.700 1688.110 1614.960 1688.430 ;
        RECT 1620.680 1688.110 1620.940 1688.430 ;
        RECT 1620.740 14.270 1620.880 1688.110 ;
        RECT 1620.680 13.950 1620.940 14.270 ;
        RECT 1721.420 13.950 1721.680 14.270 ;
        RECT 1721.480 2.400 1721.620 13.950 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1619.730 20.980 1620.050 21.040 ;
        RECT 1739.330 20.980 1739.650 21.040 ;
        RECT 1619.730 20.840 1739.650 20.980 ;
        RECT 1619.730 20.780 1620.050 20.840 ;
        RECT 1739.330 20.780 1739.650 20.840 ;
      LAYER via ;
        RECT 1619.760 20.780 1620.020 21.040 ;
        RECT 1739.360 20.780 1739.620 21.040 ;
      LAYER met2 ;
        RECT 1619.290 1700.410 1619.570 1704.000 ;
        RECT 1619.290 1700.270 1619.960 1700.410 ;
        RECT 1619.290 1700.000 1619.570 1700.270 ;
        RECT 1619.820 21.070 1619.960 1700.270 ;
        RECT 1619.760 20.750 1620.020 21.070 ;
        RECT 1739.360 20.750 1739.620 21.070 ;
        RECT 1739.420 2.400 1739.560 20.750 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1624.330 1689.020 1624.650 1689.080 ;
        RECT 1626.630 1689.020 1626.950 1689.080 ;
        RECT 1624.330 1688.880 1626.950 1689.020 ;
        RECT 1624.330 1688.820 1624.650 1688.880 ;
        RECT 1626.630 1688.820 1626.950 1688.880 ;
        RECT 1626.630 21.320 1626.950 21.380 ;
        RECT 1756.810 21.320 1757.130 21.380 ;
        RECT 1626.630 21.180 1757.130 21.320 ;
        RECT 1626.630 21.120 1626.950 21.180 ;
        RECT 1756.810 21.120 1757.130 21.180 ;
      LAYER via ;
        RECT 1624.360 1688.820 1624.620 1689.080 ;
        RECT 1626.660 1688.820 1626.920 1689.080 ;
        RECT 1626.660 21.120 1626.920 21.380 ;
        RECT 1756.840 21.120 1757.100 21.380 ;
      LAYER met2 ;
        RECT 1624.350 1700.000 1624.630 1704.000 ;
        RECT 1624.420 1689.110 1624.560 1700.000 ;
        RECT 1624.360 1688.790 1624.620 1689.110 ;
        RECT 1626.660 1688.790 1626.920 1689.110 ;
        RECT 1626.720 21.410 1626.860 1688.790 ;
        RECT 1626.660 21.090 1626.920 21.410 ;
        RECT 1756.840 21.090 1757.100 21.410 ;
        RECT 1756.900 2.400 1757.040 21.090 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1628.930 1688.000 1629.250 1688.060 ;
        RECT 1633.990 1688.000 1634.310 1688.060 ;
        RECT 1628.930 1687.860 1634.310 1688.000 ;
        RECT 1628.930 1687.800 1629.250 1687.860 ;
        RECT 1633.990 1687.800 1634.310 1687.860 ;
        RECT 1633.990 21.660 1634.310 21.720 ;
        RECT 1774.750 21.660 1775.070 21.720 ;
        RECT 1633.990 21.520 1775.070 21.660 ;
        RECT 1633.990 21.460 1634.310 21.520 ;
        RECT 1774.750 21.460 1775.070 21.520 ;
      LAYER via ;
        RECT 1628.960 1687.800 1629.220 1688.060 ;
        RECT 1634.020 1687.800 1634.280 1688.060 ;
        RECT 1634.020 21.460 1634.280 21.720 ;
        RECT 1774.780 21.460 1775.040 21.720 ;
      LAYER met2 ;
        RECT 1628.950 1700.000 1629.230 1704.000 ;
        RECT 1629.020 1688.090 1629.160 1700.000 ;
        RECT 1628.960 1687.770 1629.220 1688.090 ;
        RECT 1634.020 1687.770 1634.280 1688.090 ;
        RECT 1634.080 21.750 1634.220 1687.770 ;
        RECT 1634.020 21.430 1634.280 21.750 ;
        RECT 1774.780 21.430 1775.040 21.750 ;
        RECT 1774.840 2.400 1774.980 21.430 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 0.300 ;
=======
      LAYER met1 ;
        RECT 1633.530 22.340 1633.850 22.400 ;
        RECT 1792.690 22.340 1793.010 22.400 ;
        RECT 1633.530 22.200 1793.010 22.340 ;
        RECT 1633.530 22.140 1633.850 22.200 ;
        RECT 1792.690 22.140 1793.010 22.200 ;
      LAYER via ;
        RECT 1633.560 22.140 1633.820 22.400 ;
        RECT 1792.720 22.140 1792.980 22.400 ;
      LAYER met2 ;
        RECT 1634.010 1700.410 1634.290 1704.000 ;
        RECT 1633.620 1700.270 1634.290 1700.410 ;
        RECT 1633.620 22.430 1633.760 1700.270 ;
        RECT 1634.010 1700.000 1634.290 1700.270 ;
        RECT 1633.560 22.110 1633.820 22.430 ;
        RECT 1792.720 22.110 1792.980 22.430 ;
        RECT 1792.780 2.400 1792.920 22.110 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 0.300 ;
=======
      LAYER met1 ;
        RECT 1638.590 1688.680 1638.910 1688.740 ;
        RECT 1640.430 1688.680 1640.750 1688.740 ;
        RECT 1638.590 1688.540 1640.750 1688.680 ;
        RECT 1638.590 1688.480 1638.910 1688.540 ;
        RECT 1640.430 1688.480 1640.750 1688.540 ;
        RECT 1640.430 22.680 1640.750 22.740 ;
        RECT 1810.630 22.680 1810.950 22.740 ;
        RECT 1640.430 22.540 1810.950 22.680 ;
        RECT 1640.430 22.480 1640.750 22.540 ;
        RECT 1810.630 22.480 1810.950 22.540 ;
      LAYER via ;
        RECT 1638.620 1688.480 1638.880 1688.740 ;
        RECT 1640.460 1688.480 1640.720 1688.740 ;
        RECT 1640.460 22.480 1640.720 22.740 ;
        RECT 1810.660 22.480 1810.920 22.740 ;
      LAYER met2 ;
        RECT 1638.610 1700.000 1638.890 1704.000 ;
        RECT 1638.680 1688.770 1638.820 1700.000 ;
        RECT 1638.620 1688.450 1638.880 1688.770 ;
        RECT 1640.460 1688.450 1640.720 1688.770 ;
        RECT 1640.520 22.770 1640.660 1688.450 ;
        RECT 1640.460 22.450 1640.720 22.770 ;
        RECT 1810.660 22.450 1810.920 22.770 ;
        RECT 1810.720 2.400 1810.860 22.450 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1643.650 1688.680 1643.970 1688.740 ;
        RECT 1647.330 1688.680 1647.650 1688.740 ;
        RECT 1643.650 1688.540 1647.650 1688.680 ;
        RECT 1643.650 1688.480 1643.970 1688.540 ;
        RECT 1647.330 1688.480 1647.650 1688.540 ;
        RECT 1647.330 23.700 1647.650 23.760 ;
        RECT 1828.570 23.700 1828.890 23.760 ;
        RECT 1647.330 23.560 1828.890 23.700 ;
        RECT 1647.330 23.500 1647.650 23.560 ;
        RECT 1828.570 23.500 1828.890 23.560 ;
      LAYER via ;
        RECT 1643.680 1688.480 1643.940 1688.740 ;
        RECT 1647.360 1688.480 1647.620 1688.740 ;
        RECT 1647.360 23.500 1647.620 23.760 ;
        RECT 1828.600 23.500 1828.860 23.760 ;
      LAYER met2 ;
        RECT 1643.670 1700.000 1643.950 1704.000 ;
        RECT 1643.740 1688.770 1643.880 1700.000 ;
        RECT 1643.680 1688.450 1643.940 1688.770 ;
        RECT 1647.360 1688.450 1647.620 1688.770 ;
        RECT 1647.420 23.790 1647.560 1688.450 ;
        RECT 1647.360 23.470 1647.620 23.790 ;
        RECT 1828.600 23.470 1828.860 23.790 ;
        RECT 1828.660 2.400 1828.800 23.470 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1647.790 27.440 1648.110 27.500 ;
        RECT 1846.050 27.440 1846.370 27.500 ;
        RECT 1647.790 27.300 1846.370 27.440 ;
        RECT 1647.790 27.240 1648.110 27.300 ;
        RECT 1846.050 27.240 1846.370 27.300 ;
      LAYER via ;
        RECT 1647.820 27.240 1648.080 27.500 ;
        RECT 1846.080 27.240 1846.340 27.500 ;
      LAYER met2 ;
        RECT 1648.270 1700.410 1648.550 1704.000 ;
        RECT 1647.880 1700.270 1648.550 1700.410 ;
        RECT 1647.880 27.530 1648.020 1700.270 ;
        RECT 1648.270 1700.000 1648.550 1700.270 ;
        RECT 1647.820 27.210 1648.080 27.530 ;
        RECT 1846.080 27.210 1846.340 27.530 ;
        RECT 1846.140 2.400 1846.280 27.210 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 0.300 ;
=======
      LAYER li1 ;
        RECT 1802.425 22.865 1802.595 26.775 ;
      LAYER mcon ;
        RECT 1802.425 26.605 1802.595 26.775 ;
      LAYER met1 ;
        RECT 1654.690 26.760 1655.010 26.820 ;
        RECT 1802.365 26.760 1802.655 26.805 ;
        RECT 1654.690 26.620 1802.655 26.760 ;
        RECT 1654.690 26.560 1655.010 26.620 ;
        RECT 1802.365 26.575 1802.655 26.620 ;
        RECT 1802.365 23.020 1802.655 23.065 ;
        RECT 1863.990 23.020 1864.310 23.080 ;
        RECT 1802.365 22.880 1864.310 23.020 ;
        RECT 1802.365 22.835 1802.655 22.880 ;
        RECT 1863.990 22.820 1864.310 22.880 ;
      LAYER via ;
        RECT 1654.720 26.560 1654.980 26.820 ;
        RECT 1864.020 22.820 1864.280 23.080 ;
      LAYER met2 ;
        RECT 1652.870 1700.410 1653.150 1704.000 ;
        RECT 1652.870 1700.270 1654.460 1700.410 ;
        RECT 1652.870 1700.000 1653.150 1700.270 ;
        RECT 1654.320 1688.850 1654.460 1700.270 ;
        RECT 1654.320 1688.710 1654.920 1688.850 ;
        RECT 1654.780 26.850 1654.920 1688.710 ;
        RECT 1654.720 26.530 1654.980 26.850 ;
        RECT 1864.020 22.790 1864.280 23.110 ;
        RECT 1864.080 2.400 1864.220 22.790 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1345.570 1678.140 1345.890 1678.200 ;
        RECT 1348.330 1678.140 1348.650 1678.200 ;
        RECT 1345.570 1678.000 1348.650 1678.140 ;
        RECT 1345.570 1677.940 1345.890 1678.000 ;
        RECT 1348.330 1677.940 1348.650 1678.000 ;
        RECT 740.210 30.840 740.530 30.900 ;
        RECT 1345.570 30.840 1345.890 30.900 ;
        RECT 740.210 30.700 1345.890 30.840 ;
        RECT 740.210 30.640 740.530 30.700 ;
        RECT 1345.570 30.640 1345.890 30.700 ;
      LAYER via ;
        RECT 1345.600 1677.940 1345.860 1678.200 ;
        RECT 1348.360 1677.940 1348.620 1678.200 ;
        RECT 740.240 30.640 740.500 30.900 ;
        RECT 1345.600 30.640 1345.860 30.900 ;
      LAYER met2 ;
        RECT 1349.730 1700.410 1350.010 1704.000 ;
        RECT 1348.420 1700.270 1350.010 1700.410 ;
        RECT 1348.420 1678.230 1348.560 1700.270 ;
        RECT 1349.730 1700.000 1350.010 1700.270 ;
        RECT 1345.600 1677.910 1345.860 1678.230 ;
        RECT 1348.360 1677.910 1348.620 1678.230 ;
        RECT 1345.660 30.930 1345.800 1677.910 ;
        RECT 740.240 30.610 740.500 30.930 ;
        RECT 1345.600 30.610 1345.860 30.930 ;
        RECT 740.300 2.400 740.440 30.610 ;
        RECT 740.090 -4.800 740.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 0.300 ;
=======
      LAYER met1 ;
        RECT 1657.910 1685.620 1658.230 1685.680 ;
        RECT 1662.510 1685.620 1662.830 1685.680 ;
        RECT 1657.910 1685.480 1662.830 1685.620 ;
        RECT 1657.910 1685.420 1658.230 1685.480 ;
        RECT 1662.510 1685.420 1662.830 1685.480 ;
        RECT 1662.510 26.420 1662.830 26.480 ;
        RECT 1881.930 26.420 1882.250 26.480 ;
        RECT 1662.510 26.280 1882.250 26.420 ;
        RECT 1662.510 26.220 1662.830 26.280 ;
        RECT 1881.930 26.220 1882.250 26.280 ;
      LAYER via ;
        RECT 1657.940 1685.420 1658.200 1685.680 ;
        RECT 1662.540 1685.420 1662.800 1685.680 ;
        RECT 1662.540 26.220 1662.800 26.480 ;
        RECT 1881.960 26.220 1882.220 26.480 ;
      LAYER met2 ;
        RECT 1657.930 1700.000 1658.210 1704.000 ;
        RECT 1658.000 1685.710 1658.140 1700.000 ;
        RECT 1657.940 1685.390 1658.200 1685.710 ;
        RECT 1662.540 1685.390 1662.800 1685.710 ;
        RECT 1662.600 26.510 1662.740 1685.390 ;
        RECT 1662.540 26.190 1662.800 26.510 ;
        RECT 1881.960 26.190 1882.220 26.510 ;
        RECT 1882.020 2.400 1882.160 26.190 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1662.050 25.400 1662.370 25.460 ;
        RECT 1872.270 25.400 1872.590 25.460 ;
        RECT 1662.050 25.260 1872.590 25.400 ;
        RECT 1662.050 25.200 1662.370 25.260 ;
        RECT 1872.270 25.200 1872.590 25.260 ;
        RECT 1873.650 24.720 1873.970 24.780 ;
        RECT 1899.870 24.720 1900.190 24.780 ;
        RECT 1873.650 24.580 1900.190 24.720 ;
        RECT 1873.650 24.520 1873.970 24.580 ;
        RECT 1899.870 24.520 1900.190 24.580 ;
      LAYER via ;
        RECT 1662.080 25.200 1662.340 25.460 ;
        RECT 1872.300 25.200 1872.560 25.460 ;
        RECT 1873.680 24.520 1873.940 24.780 ;
        RECT 1899.900 24.520 1900.160 24.780 ;
      LAYER met2 ;
        RECT 1662.530 1700.410 1662.810 1704.000 ;
        RECT 1662.140 1700.270 1662.810 1700.410 ;
        RECT 1662.140 25.490 1662.280 1700.270 ;
        RECT 1662.530 1700.000 1662.810 1700.270 ;
        RECT 1662.080 25.170 1662.340 25.490 ;
        RECT 1872.300 25.170 1872.560 25.490 ;
        RECT 1872.360 24.890 1872.500 25.170 ;
        RECT 1872.360 24.810 1873.880 24.890 ;
        RECT 1872.360 24.750 1873.940 24.810 ;
        RECT 1873.680 24.490 1873.940 24.750 ;
        RECT 1899.900 24.490 1900.160 24.810 ;
        RECT 1899.960 2.400 1900.100 24.490 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1667.570 1688.340 1667.890 1688.400 ;
        RECT 1668.950 1688.340 1669.270 1688.400 ;
        RECT 1667.570 1688.200 1669.270 1688.340 ;
        RECT 1667.570 1688.140 1667.890 1688.200 ;
        RECT 1668.950 1688.140 1669.270 1688.200 ;
        RECT 1873.280 25.260 1874.340 25.400 ;
        RECT 1668.950 24.720 1669.270 24.780 ;
        RECT 1873.280 24.720 1873.420 25.260 ;
        RECT 1874.200 25.060 1874.340 25.260 ;
        RECT 1874.200 24.920 1900.560 25.060 ;
        RECT 1668.950 24.580 1873.420 24.720 ;
        RECT 1900.420 24.720 1900.560 24.920 ;
        RECT 1917.810 24.720 1918.130 24.780 ;
        RECT 1900.420 24.580 1918.130 24.720 ;
        RECT 1668.950 24.520 1669.270 24.580 ;
        RECT 1917.810 24.520 1918.130 24.580 ;
      LAYER via ;
        RECT 1667.600 1688.140 1667.860 1688.400 ;
        RECT 1668.980 1688.140 1669.240 1688.400 ;
        RECT 1668.980 24.520 1669.240 24.780 ;
        RECT 1917.840 24.520 1918.100 24.780 ;
      LAYER met2 ;
        RECT 1667.590 1700.000 1667.870 1704.000 ;
        RECT 1667.660 1688.430 1667.800 1700.000 ;
        RECT 1667.600 1688.110 1667.860 1688.430 ;
        RECT 1668.980 1688.110 1669.240 1688.430 ;
        RECT 1669.040 24.810 1669.180 1688.110 ;
        RECT 1668.980 24.490 1669.240 24.810 ;
        RECT 1917.840 24.490 1918.100 24.810 ;
        RECT 1917.900 2.400 1918.040 24.490 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 0.300 ;
=======
      LAYER li1 ;
        RECT 1919.265 24.055 1919.435 24.735 ;
        RECT 1918.345 23.885 1919.435 24.055 ;
      LAYER mcon ;
        RECT 1919.265 24.565 1919.435 24.735 ;
      LAYER met1 ;
        RECT 1672.170 1688.680 1672.490 1688.740 ;
        RECT 1675.390 1688.680 1675.710 1688.740 ;
        RECT 1672.170 1688.540 1675.710 1688.680 ;
        RECT 1672.170 1688.480 1672.490 1688.540 ;
        RECT 1675.390 1688.480 1675.710 1688.540 ;
        RECT 1919.205 24.720 1919.495 24.765 ;
        RECT 1935.290 24.720 1935.610 24.780 ;
        RECT 1919.205 24.580 1935.610 24.720 ;
        RECT 1919.205 24.535 1919.495 24.580 ;
        RECT 1935.290 24.520 1935.610 24.580 ;
        RECT 1675.390 24.040 1675.710 24.100 ;
        RECT 1918.285 24.040 1918.575 24.085 ;
        RECT 1675.390 23.900 1918.575 24.040 ;
        RECT 1675.390 23.840 1675.710 23.900 ;
        RECT 1918.285 23.855 1918.575 23.900 ;
      LAYER via ;
        RECT 1672.200 1688.480 1672.460 1688.740 ;
        RECT 1675.420 1688.480 1675.680 1688.740 ;
        RECT 1935.320 24.520 1935.580 24.780 ;
        RECT 1675.420 23.840 1675.680 24.100 ;
      LAYER met2 ;
        RECT 1672.190 1700.000 1672.470 1704.000 ;
        RECT 1672.260 1688.770 1672.400 1700.000 ;
        RECT 1672.200 1688.450 1672.460 1688.770 ;
        RECT 1675.420 1688.450 1675.680 1688.770 ;
        RECT 1675.480 24.130 1675.620 1688.450 ;
        RECT 1935.320 24.490 1935.580 24.810 ;
        RECT 1675.420 23.810 1675.680 24.130 ;
        RECT 1935.380 2.400 1935.520 24.490 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1677.230 1688.340 1677.550 1688.400 ;
        RECT 1682.750 1688.340 1683.070 1688.400 ;
        RECT 1677.230 1688.200 1683.070 1688.340 ;
        RECT 1677.230 1688.140 1677.550 1688.200 ;
        RECT 1682.750 1688.140 1683.070 1688.200 ;
      LAYER via ;
        RECT 1677.260 1688.140 1677.520 1688.400 ;
        RECT 1682.780 1688.140 1683.040 1688.400 ;
      LAYER met2 ;
        RECT 1677.250 1700.000 1677.530 1704.000 ;
        RECT 1677.320 1688.430 1677.460 1700.000 ;
        RECT 1677.260 1688.110 1677.520 1688.430 ;
        RECT 1682.780 1688.110 1683.040 1688.430 ;
        RECT 1682.840 27.725 1682.980 1688.110 ;
        RECT 1682.770 27.355 1683.050 27.725 ;
        RECT 1953.250 27.355 1953.530 27.725 ;
        RECT 1953.320 2.400 1953.460 27.355 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
      LAYER via2 ;
        RECT 1682.770 27.400 1683.050 27.680 ;
        RECT 1953.250 27.400 1953.530 27.680 ;
      LAYER met3 ;
        RECT 1682.745 27.690 1683.075 27.705 ;
        RECT 1953.225 27.690 1953.555 27.705 ;
        RECT 1682.745 27.390 1953.555 27.690 ;
        RECT 1682.745 27.375 1683.075 27.390 ;
        RECT 1953.225 27.375 1953.555 27.390 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1681.830 41.720 1682.150 41.780 ;
        RECT 1971.170 41.720 1971.490 41.780 ;
        RECT 1681.830 41.580 1971.490 41.720 ;
        RECT 1681.830 41.520 1682.150 41.580 ;
        RECT 1971.170 41.520 1971.490 41.580 ;
      LAYER via ;
        RECT 1681.860 41.520 1682.120 41.780 ;
        RECT 1971.200 41.520 1971.460 41.780 ;
      LAYER met2 ;
        RECT 1681.850 1700.000 1682.130 1704.000 ;
        RECT 1681.920 41.810 1682.060 1700.000 ;
        RECT 1681.860 41.490 1682.120 41.810 ;
        RECT 1971.200 41.490 1971.460 41.810 ;
        RECT 1971.260 2.400 1971.400 41.490 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1688.270 42.060 1688.590 42.120 ;
        RECT 1989.110 42.060 1989.430 42.120 ;
        RECT 1688.270 41.920 1989.430 42.060 ;
        RECT 1688.270 41.860 1688.590 41.920 ;
        RECT 1989.110 41.860 1989.430 41.920 ;
      LAYER via ;
        RECT 1688.300 41.860 1688.560 42.120 ;
        RECT 1989.140 41.860 1989.400 42.120 ;
      LAYER met2 ;
        RECT 1686.910 1700.410 1687.190 1704.000 ;
        RECT 1686.910 1700.270 1687.580 1700.410 ;
        RECT 1686.910 1700.000 1687.190 1700.270 ;
        RECT 1687.440 1688.680 1687.580 1700.270 ;
        RECT 1687.440 1688.540 1688.500 1688.680 ;
        RECT 1688.360 42.150 1688.500 1688.540 ;
        RECT 1688.300 41.830 1688.560 42.150 ;
        RECT 1989.140 41.830 1989.400 42.150 ;
        RECT 1989.200 2.400 1989.340 41.830 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1691.490 1688.680 1691.810 1688.740 ;
        RECT 1696.090 1688.680 1696.410 1688.740 ;
        RECT 1691.490 1688.540 1696.410 1688.680 ;
        RECT 1691.490 1688.480 1691.810 1688.540 ;
        RECT 1696.090 1688.480 1696.410 1688.540 ;
        RECT 1696.090 42.400 1696.410 42.460 ;
        RECT 2006.590 42.400 2006.910 42.460 ;
        RECT 1696.090 42.260 2006.910 42.400 ;
        RECT 1696.090 42.200 1696.410 42.260 ;
        RECT 2006.590 42.200 2006.910 42.260 ;
      LAYER via ;
        RECT 1691.520 1688.480 1691.780 1688.740 ;
        RECT 1696.120 1688.480 1696.380 1688.740 ;
        RECT 1696.120 42.200 1696.380 42.460 ;
        RECT 2006.620 42.200 2006.880 42.460 ;
      LAYER met2 ;
        RECT 1691.510 1700.000 1691.790 1704.000 ;
        RECT 1691.580 1688.770 1691.720 1700.000 ;
        RECT 1691.520 1688.450 1691.780 1688.770 ;
        RECT 1696.120 1688.450 1696.380 1688.770 ;
        RECT 1696.180 42.490 1696.320 1688.450 ;
        RECT 1696.120 42.170 1696.380 42.490 ;
        RECT 2006.620 42.170 2006.880 42.490 ;
        RECT 2006.680 2.400 2006.820 42.170 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 0.300 ;
=======
      LAYER met1 ;
        RECT 1695.630 43.080 1695.950 43.140 ;
        RECT 2024.530 43.080 2024.850 43.140 ;
        RECT 1695.630 42.940 2024.850 43.080 ;
        RECT 1695.630 42.880 1695.950 42.940 ;
        RECT 2024.530 42.880 2024.850 42.940 ;
      LAYER via ;
        RECT 1695.660 42.880 1695.920 43.140 ;
        RECT 2024.560 42.880 2024.820 43.140 ;
      LAYER met2 ;
        RECT 1696.570 1700.410 1696.850 1704.000 ;
        RECT 1695.720 1700.270 1696.850 1700.410 ;
        RECT 1695.720 43.170 1695.860 1700.270 ;
        RECT 1696.570 1700.000 1696.850 1700.270 ;
        RECT 1695.660 42.850 1695.920 43.170 ;
        RECT 2024.560 42.850 2024.820 43.170 ;
        RECT 2024.620 2.400 2024.760 42.850 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1701.150 1688.680 1701.470 1688.740 ;
        RECT 1703.450 1688.680 1703.770 1688.740 ;
        RECT 1701.150 1688.540 1703.770 1688.680 ;
        RECT 1701.150 1688.480 1701.470 1688.540 ;
        RECT 1703.450 1688.480 1703.770 1688.540 ;
        RECT 1703.450 27.780 1703.770 27.840 ;
        RECT 2042.470 27.780 2042.790 27.840 ;
        RECT 1703.450 27.640 2042.790 27.780 ;
        RECT 1703.450 27.580 1703.770 27.640 ;
        RECT 2042.470 27.580 2042.790 27.640 ;
      LAYER via ;
        RECT 1701.180 1688.480 1701.440 1688.740 ;
        RECT 1703.480 1688.480 1703.740 1688.740 ;
        RECT 1703.480 27.580 1703.740 27.840 ;
        RECT 2042.500 27.580 2042.760 27.840 ;
      LAYER met2 ;
        RECT 1701.170 1700.000 1701.450 1704.000 ;
        RECT 1701.240 1688.770 1701.380 1700.000 ;
        RECT 1701.180 1688.450 1701.440 1688.770 ;
        RECT 1703.480 1688.450 1703.740 1688.770 ;
        RECT 1703.540 27.870 1703.680 1688.450 ;
        RECT 1703.480 27.550 1703.740 27.870 ;
        RECT 2042.500 27.550 2042.760 27.870 ;
        RECT 2042.560 2.400 2042.700 27.550 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 0.300 ;
=======
      LAYER met1 ;
        RECT 757.690 31.180 758.010 31.240 ;
        RECT 1352.930 31.180 1353.250 31.240 ;
        RECT 757.690 31.040 1353.250 31.180 ;
        RECT 757.690 30.980 758.010 31.040 ;
        RECT 1352.930 30.980 1353.250 31.040 ;
      LAYER via ;
        RECT 757.720 30.980 757.980 31.240 ;
        RECT 1352.960 30.980 1353.220 31.240 ;
      LAYER met2 ;
        RECT 1354.330 1700.410 1354.610 1704.000 ;
        RECT 1353.020 1700.270 1354.610 1700.410 ;
        RECT 1353.020 31.270 1353.160 1700.270 ;
        RECT 1354.330 1700.000 1354.610 1700.270 ;
        RECT 757.720 30.950 757.980 31.270 ;
        RECT 1352.960 30.950 1353.220 31.270 ;
        RECT 757.780 2.400 757.920 30.950 ;
        RECT 757.570 -4.800 758.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1706.210 1688.000 1706.530 1688.060 ;
        RECT 1709.890 1688.000 1710.210 1688.060 ;
        RECT 1706.210 1687.860 1710.210 1688.000 ;
        RECT 1706.210 1687.800 1706.530 1687.860 ;
        RECT 1709.890 1687.800 1710.210 1687.860 ;
        RECT 1709.890 28.120 1710.210 28.180 ;
        RECT 2060.410 28.120 2060.730 28.180 ;
        RECT 1709.890 27.980 2060.730 28.120 ;
        RECT 1709.890 27.920 1710.210 27.980 ;
        RECT 2060.410 27.920 2060.730 27.980 ;
      LAYER via ;
        RECT 1706.240 1687.800 1706.500 1688.060 ;
        RECT 1709.920 1687.800 1710.180 1688.060 ;
        RECT 1709.920 27.920 1710.180 28.180 ;
        RECT 2060.440 27.920 2060.700 28.180 ;
      LAYER met2 ;
        RECT 1706.230 1700.000 1706.510 1704.000 ;
        RECT 1706.300 1688.090 1706.440 1700.000 ;
        RECT 1706.240 1687.770 1706.500 1688.090 ;
        RECT 1709.920 1687.770 1710.180 1688.090 ;
        RECT 1709.980 28.210 1710.120 1687.770 ;
        RECT 1709.920 27.890 1710.180 28.210 ;
        RECT 2060.440 27.890 2060.700 28.210 ;
        RECT 2060.500 2.400 2060.640 27.890 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 0.300 ;
=======
      LAYER met1 ;
        RECT 1709.430 28.460 1709.750 28.520 ;
        RECT 2078.350 28.460 2078.670 28.520 ;
        RECT 1709.430 28.320 2078.670 28.460 ;
        RECT 1709.430 28.260 1709.750 28.320 ;
        RECT 2078.350 28.260 2078.670 28.320 ;
      LAYER via ;
        RECT 1709.460 28.260 1709.720 28.520 ;
        RECT 2078.380 28.260 2078.640 28.520 ;
      LAYER met2 ;
        RECT 1710.830 1700.410 1711.110 1704.000 ;
        RECT 1709.980 1700.270 1711.110 1700.410 ;
        RECT 1709.980 1688.680 1710.120 1700.270 ;
        RECT 1710.830 1700.000 1711.110 1700.270 ;
        RECT 1709.520 1688.540 1710.120 1688.680 ;
        RECT 1709.520 28.550 1709.660 1688.540 ;
        RECT 1709.460 28.230 1709.720 28.550 ;
        RECT 2078.380 28.230 2078.640 28.550 ;
        RECT 2078.440 2.400 2078.580 28.230 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1715.870 1688.000 1716.190 1688.060 ;
        RECT 1717.710 1688.000 1718.030 1688.060 ;
        RECT 1715.870 1687.860 1718.030 1688.000 ;
        RECT 1715.870 1687.800 1716.190 1687.860 ;
        RECT 1717.710 1687.800 1718.030 1687.860 ;
        RECT 1717.710 28.800 1718.030 28.860 ;
        RECT 2095.830 28.800 2096.150 28.860 ;
        RECT 1717.710 28.660 2096.150 28.800 ;
        RECT 1717.710 28.600 1718.030 28.660 ;
        RECT 2095.830 28.600 2096.150 28.660 ;
      LAYER via ;
        RECT 1715.900 1687.800 1716.160 1688.060 ;
        RECT 1717.740 1687.800 1718.000 1688.060 ;
        RECT 1717.740 28.600 1718.000 28.860 ;
        RECT 2095.860 28.600 2096.120 28.860 ;
      LAYER met2 ;
        RECT 1715.890 1700.000 1716.170 1704.000 ;
        RECT 1715.960 1688.090 1716.100 1700.000 ;
        RECT 1715.900 1687.770 1716.160 1688.090 ;
        RECT 1717.740 1687.770 1718.000 1688.090 ;
        RECT 1717.800 28.890 1717.940 1687.770 ;
        RECT 1717.740 28.570 1718.000 28.890 ;
        RECT 2095.860 28.570 2096.120 28.890 ;
        RECT 2095.920 2.400 2096.060 28.570 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 0.300 ;
=======
      LAYER met1 ;
        RECT 1720.470 1688.680 1720.790 1688.740 ;
        RECT 1724.610 1688.680 1724.930 1688.740 ;
        RECT 1720.470 1688.540 1724.930 1688.680 ;
        RECT 1720.470 1688.480 1720.790 1688.540 ;
        RECT 1724.610 1688.480 1724.930 1688.540 ;
        RECT 1724.610 29.140 1724.930 29.200 ;
        RECT 2113.770 29.140 2114.090 29.200 ;
        RECT 1724.610 29.000 2114.090 29.140 ;
        RECT 1724.610 28.940 1724.930 29.000 ;
        RECT 2113.770 28.940 2114.090 29.000 ;
      LAYER via ;
        RECT 1720.500 1688.480 1720.760 1688.740 ;
        RECT 1724.640 1688.480 1724.900 1688.740 ;
        RECT 1724.640 28.940 1724.900 29.200 ;
        RECT 2113.800 28.940 2114.060 29.200 ;
      LAYER met2 ;
        RECT 1720.490 1700.000 1720.770 1704.000 ;
        RECT 1720.560 1688.770 1720.700 1700.000 ;
        RECT 1720.500 1688.450 1720.760 1688.770 ;
        RECT 1724.640 1688.450 1724.900 1688.770 ;
        RECT 1724.700 29.230 1724.840 1688.450 ;
        RECT 1724.640 28.910 1724.900 29.230 ;
        RECT 2113.800 28.910 2114.060 29.230 ;
        RECT 2113.860 2.400 2114.000 28.910 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 0.300 ;
=======
      LAYER met1 ;
        RECT 1725.530 1688.000 1725.850 1688.060 ;
        RECT 1731.050 1688.000 1731.370 1688.060 ;
        RECT 1725.530 1687.860 1731.370 1688.000 ;
        RECT 1725.530 1687.800 1725.850 1687.860 ;
        RECT 1731.050 1687.800 1731.370 1687.860 ;
        RECT 1731.050 29.480 1731.370 29.540 ;
        RECT 2131.710 29.480 2132.030 29.540 ;
        RECT 1731.050 29.340 2132.030 29.480 ;
        RECT 1731.050 29.280 1731.370 29.340 ;
        RECT 2131.710 29.280 2132.030 29.340 ;
      LAYER via ;
        RECT 1725.560 1687.800 1725.820 1688.060 ;
        RECT 1731.080 1687.800 1731.340 1688.060 ;
        RECT 1731.080 29.280 1731.340 29.540 ;
        RECT 2131.740 29.280 2132.000 29.540 ;
      LAYER met2 ;
        RECT 1725.550 1700.000 1725.830 1704.000 ;
        RECT 1725.620 1688.090 1725.760 1700.000 ;
        RECT 1725.560 1687.770 1725.820 1688.090 ;
        RECT 1731.080 1687.770 1731.340 1688.090 ;
        RECT 1731.140 29.570 1731.280 1687.770 ;
        RECT 1731.080 29.250 1731.340 29.570 ;
        RECT 2131.740 29.250 2132.000 29.570 ;
        RECT 2131.800 2.400 2131.940 29.250 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1730.590 29.820 1730.910 29.880 ;
        RECT 2149.650 29.820 2149.970 29.880 ;
        RECT 1730.590 29.680 2149.970 29.820 ;
        RECT 1730.590 29.620 1730.910 29.680 ;
        RECT 2149.650 29.620 2149.970 29.680 ;
      LAYER via ;
        RECT 1730.620 29.620 1730.880 29.880 ;
        RECT 2149.680 29.620 2149.940 29.880 ;
      LAYER met2 ;
        RECT 1730.150 1700.410 1730.430 1704.000 ;
        RECT 1730.150 1700.270 1730.820 1700.410 ;
        RECT 1730.150 1700.000 1730.430 1700.270 ;
        RECT 1730.680 29.910 1730.820 1700.270 ;
        RECT 1730.620 29.590 1730.880 29.910 ;
        RECT 2149.680 29.590 2149.940 29.910 ;
        RECT 2149.740 2.400 2149.880 29.590 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1735.190 1688.680 1735.510 1688.740 ;
        RECT 1738.410 1688.680 1738.730 1688.740 ;
        RECT 1735.190 1688.540 1738.730 1688.680 ;
        RECT 1735.190 1688.480 1735.510 1688.540 ;
        RECT 1738.410 1688.480 1738.730 1688.540 ;
        RECT 1738.410 30.160 1738.730 30.220 ;
        RECT 2167.590 30.160 2167.910 30.220 ;
        RECT 1738.410 30.020 2167.910 30.160 ;
        RECT 1738.410 29.960 1738.730 30.020 ;
        RECT 2167.590 29.960 2167.910 30.020 ;
      LAYER via ;
        RECT 1735.220 1688.480 1735.480 1688.740 ;
        RECT 1738.440 1688.480 1738.700 1688.740 ;
        RECT 1738.440 29.960 1738.700 30.220 ;
        RECT 2167.620 29.960 2167.880 30.220 ;
      LAYER met2 ;
        RECT 1735.210 1700.000 1735.490 1704.000 ;
        RECT 1735.280 1688.770 1735.420 1700.000 ;
        RECT 1735.220 1688.450 1735.480 1688.770 ;
        RECT 1738.440 1688.450 1738.700 1688.770 ;
        RECT 1738.500 30.250 1738.640 1688.450 ;
        RECT 1738.440 29.930 1738.700 30.250 ;
        RECT 2167.620 29.930 2167.880 30.250 ;
        RECT 2167.680 2.400 2167.820 29.930 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 0.300 ;
=======
      LAYER met1 ;
        RECT 1739.790 1688.680 1740.110 1688.740 ;
        RECT 1744.850 1688.680 1745.170 1688.740 ;
        RECT 1739.790 1688.540 1745.170 1688.680 ;
        RECT 1739.790 1688.480 1740.110 1688.540 ;
        RECT 1744.850 1688.480 1745.170 1688.540 ;
        RECT 1744.850 30.500 1745.170 30.560 ;
        RECT 2185.070 30.500 2185.390 30.560 ;
        RECT 1744.850 30.360 2185.390 30.500 ;
        RECT 1744.850 30.300 1745.170 30.360 ;
        RECT 2185.070 30.300 2185.390 30.360 ;
      LAYER via ;
        RECT 1739.820 1688.480 1740.080 1688.740 ;
        RECT 1744.880 1688.480 1745.140 1688.740 ;
        RECT 1744.880 30.300 1745.140 30.560 ;
        RECT 2185.100 30.300 2185.360 30.560 ;
      LAYER met2 ;
        RECT 1739.810 1700.000 1740.090 1704.000 ;
        RECT 1739.880 1688.770 1740.020 1700.000 ;
        RECT 1739.820 1688.450 1740.080 1688.770 ;
        RECT 1744.880 1688.450 1745.140 1688.770 ;
        RECT 1744.940 30.590 1745.080 1688.450 ;
        RECT 1744.880 30.270 1745.140 30.590 ;
        RECT 2185.100 30.270 2185.360 30.590 ;
        RECT 2185.160 2.400 2185.300 30.270 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1745.310 34.240 1745.630 34.300 ;
        RECT 2203.010 34.240 2203.330 34.300 ;
        RECT 1745.310 34.100 2203.330 34.240 ;
        RECT 1745.310 34.040 1745.630 34.100 ;
        RECT 2203.010 34.040 2203.330 34.100 ;
      LAYER via ;
        RECT 1745.340 34.040 1745.600 34.300 ;
        RECT 2203.040 34.040 2203.300 34.300 ;
      LAYER met2 ;
        RECT 1744.870 1700.410 1745.150 1704.000 ;
        RECT 1744.870 1700.270 1745.540 1700.410 ;
        RECT 1744.870 1700.000 1745.150 1700.270 ;
        RECT 1745.400 34.330 1745.540 1700.270 ;
        RECT 1745.340 34.010 1745.600 34.330 ;
        RECT 2203.040 34.010 2203.300 34.330 ;
        RECT 2203.100 2.400 2203.240 34.010 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1749.450 1688.680 1749.770 1688.740 ;
        RECT 1751.750 1688.680 1752.070 1688.740 ;
        RECT 1749.450 1688.540 1752.070 1688.680 ;
        RECT 1749.450 1688.480 1749.770 1688.540 ;
        RECT 1751.750 1688.480 1752.070 1688.540 ;
        RECT 1751.750 33.900 1752.070 33.960 ;
        RECT 2220.950 33.900 2221.270 33.960 ;
        RECT 1751.750 33.760 2221.270 33.900 ;
        RECT 1751.750 33.700 1752.070 33.760 ;
        RECT 2220.950 33.700 2221.270 33.760 ;
      LAYER via ;
        RECT 1749.480 1688.480 1749.740 1688.740 ;
        RECT 1751.780 1688.480 1752.040 1688.740 ;
        RECT 1751.780 33.700 1752.040 33.960 ;
        RECT 2220.980 33.700 2221.240 33.960 ;
      LAYER met2 ;
        RECT 1749.470 1700.000 1749.750 1704.000 ;
        RECT 1749.540 1688.770 1749.680 1700.000 ;
        RECT 1749.480 1688.450 1749.740 1688.770 ;
        RECT 1751.780 1688.450 1752.040 1688.770 ;
        RECT 1751.840 33.990 1751.980 1688.450 ;
        RECT 1751.780 33.670 1752.040 33.990 ;
        RECT 2220.980 33.670 2221.240 33.990 ;
        RECT 2221.040 2.400 2221.180 33.670 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 0.300 ;
=======
      LAYER li1 ;
        RECT 1354.385 1607.605 1354.555 1642.115 ;
        RECT 1354.385 1545.725 1354.555 1593.835 ;
        RECT 1354.385 1400.885 1354.555 1414.995 ;
        RECT 1354.385 1207.425 1354.555 1255.875 ;
        RECT 1354.385 1062.585 1354.555 1110.695 ;
        RECT 1354.385 821.185 1354.555 910.775 ;
        RECT 1354.385 766.105 1354.555 814.215 ;
        RECT 1354.385 524.365 1354.555 572.475 ;
        RECT 1354.845 469.285 1355.015 517.395 ;
      LAYER mcon ;
        RECT 1354.385 1641.945 1354.555 1642.115 ;
        RECT 1354.385 1593.665 1354.555 1593.835 ;
        RECT 1354.385 1414.825 1354.555 1414.995 ;
        RECT 1354.385 1255.705 1354.555 1255.875 ;
        RECT 1354.385 1110.525 1354.555 1110.695 ;
        RECT 1354.385 910.605 1354.555 910.775 ;
        RECT 1354.385 814.045 1354.555 814.215 ;
        RECT 1354.385 572.305 1354.555 572.475 ;
        RECT 1354.845 517.225 1355.015 517.395 ;
      LAYER met1 ;
        RECT 1354.310 1642.100 1354.630 1642.160 ;
        RECT 1354.115 1641.960 1354.630 1642.100 ;
        RECT 1354.310 1641.900 1354.630 1641.960 ;
        RECT 1354.310 1607.760 1354.630 1607.820 ;
        RECT 1354.115 1607.620 1354.630 1607.760 ;
        RECT 1354.310 1607.560 1354.630 1607.620 ;
        RECT 1354.310 1593.820 1354.630 1593.880 ;
        RECT 1354.115 1593.680 1354.630 1593.820 ;
        RECT 1354.310 1593.620 1354.630 1593.680 ;
        RECT 1354.325 1545.880 1354.615 1545.925 ;
        RECT 1354.770 1545.880 1355.090 1545.940 ;
        RECT 1354.325 1545.740 1355.090 1545.880 ;
        RECT 1354.325 1545.695 1354.615 1545.740 ;
        RECT 1354.770 1545.680 1355.090 1545.740 ;
        RECT 1354.325 1414.980 1354.615 1415.025 ;
        RECT 1354.770 1414.980 1355.090 1415.040 ;
        RECT 1354.325 1414.840 1355.090 1414.980 ;
        RECT 1354.325 1414.795 1354.615 1414.840 ;
        RECT 1354.770 1414.780 1355.090 1414.840 ;
        RECT 1354.310 1401.040 1354.630 1401.100 ;
        RECT 1354.115 1400.900 1354.630 1401.040 ;
        RECT 1354.310 1400.840 1354.630 1400.900 ;
        RECT 1354.770 1304.820 1355.090 1304.880 ;
        RECT 1354.400 1304.680 1355.090 1304.820 ;
        RECT 1354.400 1304.540 1354.540 1304.680 ;
        RECT 1354.770 1304.620 1355.090 1304.680 ;
        RECT 1354.310 1304.280 1354.630 1304.540 ;
        RECT 1354.310 1255.860 1354.630 1255.920 ;
        RECT 1354.115 1255.720 1354.630 1255.860 ;
        RECT 1354.310 1255.660 1354.630 1255.720 ;
        RECT 1354.310 1207.580 1354.630 1207.640 ;
        RECT 1354.115 1207.440 1354.630 1207.580 ;
        RECT 1354.310 1207.380 1354.630 1207.440 ;
        RECT 1354.310 1110.680 1354.630 1110.740 ;
        RECT 1354.115 1110.540 1354.630 1110.680 ;
        RECT 1354.310 1110.480 1354.630 1110.540 ;
        RECT 1354.325 1062.740 1354.615 1062.785 ;
        RECT 1354.770 1062.740 1355.090 1062.800 ;
        RECT 1354.325 1062.600 1355.090 1062.740 ;
        RECT 1354.325 1062.555 1354.615 1062.600 ;
        RECT 1354.770 1062.540 1355.090 1062.600 ;
        RECT 1354.310 918.240 1354.630 918.300 ;
        RECT 1354.770 918.240 1355.090 918.300 ;
        RECT 1354.310 918.100 1355.090 918.240 ;
        RECT 1354.310 918.040 1354.630 918.100 ;
        RECT 1354.770 918.040 1355.090 918.100 ;
        RECT 1354.310 910.760 1354.630 910.820 ;
        RECT 1354.115 910.620 1354.630 910.760 ;
        RECT 1354.310 910.560 1354.630 910.620 ;
        RECT 1354.310 821.340 1354.630 821.400 ;
        RECT 1354.115 821.200 1354.630 821.340 ;
        RECT 1354.310 821.140 1354.630 821.200 ;
        RECT 1354.310 814.200 1354.630 814.260 ;
        RECT 1354.115 814.060 1354.630 814.200 ;
        RECT 1354.310 814.000 1354.630 814.060 ;
        RECT 1354.310 766.260 1354.630 766.320 ;
        RECT 1354.115 766.120 1354.630 766.260 ;
        RECT 1354.310 766.060 1354.630 766.120 ;
        RECT 1354.310 765.580 1354.630 765.640 ;
        RECT 1355.230 765.580 1355.550 765.640 ;
        RECT 1354.310 765.440 1355.550 765.580 ;
        RECT 1354.310 765.380 1354.630 765.440 ;
        RECT 1355.230 765.380 1355.550 765.440 ;
        RECT 1354.310 717.640 1354.630 717.700 ;
        RECT 1354.770 717.640 1355.090 717.700 ;
        RECT 1354.310 717.500 1355.090 717.640 ;
        RECT 1354.310 717.440 1354.630 717.500 ;
        RECT 1354.770 717.440 1355.090 717.500 ;
        RECT 1354.310 572.460 1354.630 572.520 ;
        RECT 1354.115 572.320 1354.630 572.460 ;
        RECT 1354.310 572.260 1354.630 572.320 ;
        RECT 1354.325 524.520 1354.615 524.565 ;
        RECT 1354.770 524.520 1355.090 524.580 ;
        RECT 1354.325 524.380 1355.090 524.520 ;
        RECT 1354.325 524.335 1354.615 524.380 ;
        RECT 1354.770 524.320 1355.090 524.380 ;
        RECT 1354.770 517.380 1355.090 517.440 ;
        RECT 1354.575 517.240 1355.090 517.380 ;
        RECT 1354.770 517.180 1355.090 517.240 ;
        RECT 1354.770 469.440 1355.090 469.500 ;
        RECT 1354.575 469.300 1355.090 469.440 ;
        RECT 1354.770 469.240 1355.090 469.300 ;
        RECT 1354.310 427.960 1354.630 428.020 ;
        RECT 1354.770 427.960 1355.090 428.020 ;
        RECT 1354.310 427.820 1355.090 427.960 ;
        RECT 1354.310 427.760 1354.630 427.820 ;
        RECT 1354.770 427.760 1355.090 427.820 ;
        RECT 1354.310 283.120 1354.630 283.180 ;
        RECT 1354.770 283.120 1355.090 283.180 ;
        RECT 1354.310 282.980 1355.090 283.120 ;
        RECT 1354.310 282.920 1354.630 282.980 ;
        RECT 1354.770 282.920 1355.090 282.980 ;
        RECT 775.630 31.520 775.950 31.580 ;
        RECT 1354.770 31.520 1355.090 31.580 ;
        RECT 775.630 31.380 1355.090 31.520 ;
        RECT 775.630 31.320 775.950 31.380 ;
        RECT 1354.770 31.320 1355.090 31.380 ;
      LAYER via ;
        RECT 1354.340 1641.900 1354.600 1642.160 ;
        RECT 1354.340 1607.560 1354.600 1607.820 ;
        RECT 1354.340 1593.620 1354.600 1593.880 ;
        RECT 1354.800 1545.680 1355.060 1545.940 ;
        RECT 1354.800 1414.780 1355.060 1415.040 ;
        RECT 1354.340 1400.840 1354.600 1401.100 ;
        RECT 1354.800 1304.620 1355.060 1304.880 ;
        RECT 1354.340 1304.280 1354.600 1304.540 ;
        RECT 1354.340 1255.660 1354.600 1255.920 ;
        RECT 1354.340 1207.380 1354.600 1207.640 ;
        RECT 1354.340 1110.480 1354.600 1110.740 ;
        RECT 1354.800 1062.540 1355.060 1062.800 ;
        RECT 1354.340 918.040 1354.600 918.300 ;
        RECT 1354.800 918.040 1355.060 918.300 ;
        RECT 1354.340 910.560 1354.600 910.820 ;
        RECT 1354.340 821.140 1354.600 821.400 ;
        RECT 1354.340 814.000 1354.600 814.260 ;
        RECT 1354.340 766.060 1354.600 766.320 ;
        RECT 1354.340 765.380 1354.600 765.640 ;
        RECT 1355.260 765.380 1355.520 765.640 ;
        RECT 1354.340 717.440 1354.600 717.700 ;
        RECT 1354.800 717.440 1355.060 717.700 ;
        RECT 1354.340 572.260 1354.600 572.520 ;
        RECT 1354.800 524.320 1355.060 524.580 ;
        RECT 1354.800 517.180 1355.060 517.440 ;
        RECT 1354.800 469.240 1355.060 469.500 ;
        RECT 1354.340 427.760 1354.600 428.020 ;
        RECT 1354.800 427.760 1355.060 428.020 ;
        RECT 1354.340 282.920 1354.600 283.180 ;
        RECT 1354.800 282.920 1355.060 283.180 ;
        RECT 775.660 31.320 775.920 31.580 ;
        RECT 1354.800 31.320 1355.060 31.580 ;
      LAYER met2 ;
        RECT 1358.930 1700.410 1359.210 1704.000 ;
        RECT 1358.540 1700.270 1359.210 1700.410 ;
        RECT 1358.540 1676.610 1358.680 1700.270 ;
        RECT 1358.930 1700.000 1359.210 1700.270 ;
        RECT 1354.400 1676.470 1358.680 1676.610 ;
        RECT 1354.400 1642.190 1354.540 1676.470 ;
        RECT 1354.340 1641.870 1354.600 1642.190 ;
        RECT 1354.340 1607.530 1354.600 1607.850 ;
        RECT 1354.400 1593.910 1354.540 1607.530 ;
        RECT 1354.340 1593.590 1354.600 1593.910 ;
        RECT 1354.800 1545.650 1355.060 1545.970 ;
        RECT 1354.860 1415.070 1355.000 1545.650 ;
        RECT 1354.800 1414.750 1355.060 1415.070 ;
        RECT 1354.340 1400.810 1354.600 1401.130 ;
        RECT 1354.400 1352.250 1354.540 1400.810 ;
        RECT 1354.400 1352.110 1355.000 1352.250 ;
        RECT 1354.860 1304.910 1355.000 1352.110 ;
        RECT 1354.800 1304.590 1355.060 1304.910 ;
        RECT 1354.340 1304.250 1354.600 1304.570 ;
        RECT 1354.400 1255.950 1354.540 1304.250 ;
        RECT 1354.340 1255.630 1354.600 1255.950 ;
        RECT 1354.340 1207.350 1354.600 1207.670 ;
        RECT 1354.400 1110.770 1354.540 1207.350 ;
        RECT 1354.340 1110.450 1354.600 1110.770 ;
        RECT 1354.800 1062.510 1355.060 1062.830 ;
        RECT 1354.860 918.330 1355.000 1062.510 ;
        RECT 1354.340 918.010 1354.600 918.330 ;
        RECT 1354.800 918.010 1355.060 918.330 ;
        RECT 1354.400 910.850 1354.540 918.010 ;
        RECT 1354.340 910.530 1354.600 910.850 ;
        RECT 1354.340 821.110 1354.600 821.430 ;
        RECT 1354.400 814.290 1354.540 821.110 ;
        RECT 1354.340 813.970 1354.600 814.290 ;
        RECT 1354.340 766.030 1354.600 766.350 ;
        RECT 1354.400 765.670 1354.540 766.030 ;
        RECT 1354.340 765.350 1354.600 765.670 ;
        RECT 1355.260 765.350 1355.520 765.670 ;
        RECT 1355.320 717.925 1355.460 765.350 ;
        RECT 1354.330 717.555 1354.610 717.925 ;
        RECT 1354.340 717.410 1354.600 717.555 ;
        RECT 1354.800 717.410 1355.060 717.730 ;
        RECT 1355.250 717.555 1355.530 717.925 ;
        RECT 1354.860 671.005 1355.000 717.410 ;
        RECT 1354.790 670.635 1355.070 671.005 ;
        RECT 1354.330 669.275 1354.610 669.645 ;
        RECT 1354.400 572.550 1354.540 669.275 ;
        RECT 1354.340 572.230 1354.600 572.550 ;
        RECT 1354.800 524.290 1355.060 524.610 ;
        RECT 1354.860 517.470 1355.000 524.290 ;
        RECT 1354.800 517.150 1355.060 517.470 ;
        RECT 1354.800 469.210 1355.060 469.530 ;
        RECT 1354.860 428.050 1355.000 469.210 ;
        RECT 1354.340 427.730 1354.600 428.050 ;
        RECT 1354.800 427.730 1355.060 428.050 ;
        RECT 1354.400 283.210 1354.540 427.730 ;
        RECT 1354.340 282.890 1354.600 283.210 ;
        RECT 1354.800 282.890 1355.060 283.210 ;
        RECT 1354.860 207.130 1355.000 282.890 ;
        RECT 1354.400 206.990 1355.000 207.130 ;
        RECT 1354.400 144.685 1354.540 206.990 ;
        RECT 1354.330 144.315 1354.610 144.685 ;
        RECT 1354.790 143.635 1355.070 144.005 ;
        RECT 1354.860 31.610 1355.000 143.635 ;
        RECT 775.660 31.290 775.920 31.610 ;
        RECT 1354.800 31.290 1355.060 31.610 ;
        RECT 775.720 2.400 775.860 31.290 ;
        RECT 775.510 -4.800 776.070 2.400 ;
      LAYER via2 ;
        RECT 1354.330 717.600 1354.610 717.880 ;
        RECT 1355.250 717.600 1355.530 717.880 ;
        RECT 1354.790 670.680 1355.070 670.960 ;
        RECT 1354.330 669.320 1354.610 669.600 ;
        RECT 1354.330 144.360 1354.610 144.640 ;
        RECT 1354.790 143.680 1355.070 143.960 ;
      LAYER met3 ;
        RECT 1354.305 717.890 1354.635 717.905 ;
        RECT 1355.225 717.890 1355.555 717.905 ;
        RECT 1354.305 717.590 1355.555 717.890 ;
        RECT 1354.305 717.575 1354.635 717.590 ;
        RECT 1355.225 717.575 1355.555 717.590 ;
        RECT 1354.765 670.970 1355.095 670.985 ;
        RECT 1353.630 670.670 1355.095 670.970 ;
        RECT 1353.630 669.610 1353.930 670.670 ;
        RECT 1354.765 670.655 1355.095 670.670 ;
        RECT 1354.305 669.610 1354.635 669.625 ;
        RECT 1353.630 669.310 1354.635 669.610 ;
        RECT 1354.305 669.295 1354.635 669.310 ;
        RECT 1354.305 144.650 1354.635 144.665 ;
        RECT 1353.630 144.350 1354.635 144.650 ;
        RECT 1353.630 143.970 1353.930 144.350 ;
        RECT 1354.305 144.335 1354.635 144.350 ;
        RECT 1354.765 143.970 1355.095 143.985 ;
        RECT 1353.630 143.670 1355.095 143.970 ;
        RECT 1354.765 143.655 1355.095 143.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1754.050 1685.280 1754.370 1685.340 ;
        RECT 1758.190 1685.280 1758.510 1685.340 ;
        RECT 1754.050 1685.140 1758.510 1685.280 ;
        RECT 1754.050 1685.080 1754.370 1685.140 ;
        RECT 1758.190 1685.080 1758.510 1685.140 ;
        RECT 1758.190 33.560 1758.510 33.620 ;
        RECT 2238.890 33.560 2239.210 33.620 ;
        RECT 1758.190 33.420 2239.210 33.560 ;
        RECT 1758.190 33.360 1758.510 33.420 ;
        RECT 2238.890 33.360 2239.210 33.420 ;
      LAYER via ;
        RECT 1754.080 1685.080 1754.340 1685.340 ;
        RECT 1758.220 1685.080 1758.480 1685.340 ;
        RECT 1758.220 33.360 1758.480 33.620 ;
        RECT 2238.920 33.360 2239.180 33.620 ;
      LAYER met2 ;
        RECT 1754.070 1700.000 1754.350 1704.000 ;
        RECT 1754.140 1685.370 1754.280 1700.000 ;
        RECT 1754.080 1685.050 1754.340 1685.370 ;
        RECT 1758.220 1685.050 1758.480 1685.370 ;
        RECT 1758.280 33.650 1758.420 1685.050 ;
        RECT 1758.220 33.330 1758.480 33.650 ;
        RECT 2238.920 33.330 2239.180 33.650 ;
        RECT 2238.980 2.400 2239.120 33.330 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1758.650 33.220 1758.970 33.280 ;
        RECT 2256.370 33.220 2256.690 33.280 ;
        RECT 1758.650 33.080 2256.690 33.220 ;
        RECT 1758.650 33.020 1758.970 33.080 ;
        RECT 2256.370 33.020 2256.690 33.080 ;
      LAYER via ;
        RECT 1758.680 33.020 1758.940 33.280 ;
        RECT 2256.400 33.020 2256.660 33.280 ;
      LAYER met2 ;
        RECT 1759.130 1700.410 1759.410 1704.000 ;
        RECT 1758.740 1700.270 1759.410 1700.410 ;
        RECT 1758.740 33.310 1758.880 1700.270 ;
        RECT 1759.130 1700.000 1759.410 1700.270 ;
        RECT 1758.680 32.990 1758.940 33.310 ;
        RECT 2256.400 32.990 2256.660 33.310 ;
        RECT 2256.460 2.400 2256.600 32.990 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1763.710 1685.960 1764.030 1686.020 ;
        RECT 1766.010 1685.960 1766.330 1686.020 ;
        RECT 1763.710 1685.820 1766.330 1685.960 ;
        RECT 1763.710 1685.760 1764.030 1685.820 ;
        RECT 1766.010 1685.760 1766.330 1685.820 ;
        RECT 1766.010 32.880 1766.330 32.940 ;
        RECT 2274.310 32.880 2274.630 32.940 ;
        RECT 1766.010 32.740 2274.630 32.880 ;
        RECT 1766.010 32.680 1766.330 32.740 ;
        RECT 2274.310 32.680 2274.630 32.740 ;
      LAYER via ;
        RECT 1763.740 1685.760 1764.000 1686.020 ;
        RECT 1766.040 1685.760 1766.300 1686.020 ;
        RECT 1766.040 32.680 1766.300 32.940 ;
        RECT 2274.340 32.680 2274.600 32.940 ;
      LAYER met2 ;
        RECT 1763.730 1700.000 1764.010 1704.000 ;
        RECT 1763.800 1686.050 1763.940 1700.000 ;
        RECT 1763.740 1685.730 1764.000 1686.050 ;
        RECT 1766.040 1685.730 1766.300 1686.050 ;
        RECT 1766.100 32.970 1766.240 1685.730 ;
        RECT 1766.040 32.650 1766.300 32.970 ;
        RECT 2274.340 32.650 2274.600 32.970 ;
        RECT 2274.400 2.400 2274.540 32.650 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1768.770 1686.640 1769.090 1686.700 ;
        RECT 1772.450 1686.640 1772.770 1686.700 ;
        RECT 1768.770 1686.500 1772.770 1686.640 ;
        RECT 1768.770 1686.440 1769.090 1686.500 ;
        RECT 1772.450 1686.440 1772.770 1686.500 ;
        RECT 1772.450 32.540 1772.770 32.600 ;
        RECT 2292.250 32.540 2292.570 32.600 ;
        RECT 1772.450 32.400 2292.570 32.540 ;
        RECT 1772.450 32.340 1772.770 32.400 ;
        RECT 2292.250 32.340 2292.570 32.400 ;
      LAYER via ;
        RECT 1768.800 1686.440 1769.060 1686.700 ;
        RECT 1772.480 1686.440 1772.740 1686.700 ;
        RECT 1772.480 32.340 1772.740 32.600 ;
        RECT 2292.280 32.340 2292.540 32.600 ;
      LAYER met2 ;
        RECT 1768.790 1700.000 1769.070 1704.000 ;
        RECT 1768.860 1686.730 1769.000 1700.000 ;
        RECT 1768.800 1686.410 1769.060 1686.730 ;
        RECT 1772.480 1686.410 1772.740 1686.730 ;
        RECT 1772.540 32.630 1772.680 1686.410 ;
        RECT 1772.480 32.310 1772.740 32.630 ;
        RECT 2292.280 32.310 2292.540 32.630 ;
        RECT 2292.340 2.400 2292.480 32.310 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 0.300 ;
=======
      LAYER met1 ;
        RECT 1773.370 1687.660 1773.690 1687.720 ;
        RECT 1778.890 1687.660 1779.210 1687.720 ;
        RECT 1773.370 1687.520 1779.210 1687.660 ;
        RECT 1773.370 1687.460 1773.690 1687.520 ;
        RECT 1778.890 1687.460 1779.210 1687.520 ;
        RECT 1778.890 32.200 1779.210 32.260 ;
        RECT 2310.190 32.200 2310.510 32.260 ;
        RECT 1778.890 32.060 2310.510 32.200 ;
        RECT 1778.890 32.000 1779.210 32.060 ;
        RECT 2310.190 32.000 2310.510 32.060 ;
      LAYER via ;
        RECT 1773.400 1687.460 1773.660 1687.720 ;
        RECT 1778.920 1687.460 1779.180 1687.720 ;
        RECT 1778.920 32.000 1779.180 32.260 ;
        RECT 2310.220 32.000 2310.480 32.260 ;
      LAYER met2 ;
        RECT 1773.390 1700.000 1773.670 1704.000 ;
        RECT 1773.460 1687.750 1773.600 1700.000 ;
        RECT 1773.400 1687.430 1773.660 1687.750 ;
        RECT 1778.920 1687.430 1779.180 1687.750 ;
        RECT 1778.980 32.290 1779.120 1687.430 ;
        RECT 1778.920 31.970 1779.180 32.290 ;
        RECT 2310.220 31.970 2310.480 32.290 ;
        RECT 2310.280 2.400 2310.420 31.970 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1779.350 31.860 1779.670 31.920 ;
        RECT 2328.130 31.860 2328.450 31.920 ;
        RECT 1779.350 31.720 2328.450 31.860 ;
        RECT 1779.350 31.660 1779.670 31.720 ;
        RECT 2328.130 31.660 2328.450 31.720 ;
      LAYER via ;
        RECT 1779.380 31.660 1779.640 31.920 ;
        RECT 2328.160 31.660 2328.420 31.920 ;
      LAYER met2 ;
        RECT 1778.450 1700.410 1778.730 1704.000 ;
        RECT 1778.450 1700.270 1779.580 1700.410 ;
        RECT 1778.450 1700.000 1778.730 1700.270 ;
        RECT 1779.440 31.950 1779.580 1700.270 ;
        RECT 1779.380 31.630 1779.640 31.950 ;
        RECT 2328.160 31.630 2328.420 31.950 ;
        RECT 2328.220 2.400 2328.360 31.630 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1783.030 1686.980 1783.350 1687.040 ;
        RECT 1786.250 1686.980 1786.570 1687.040 ;
        RECT 1783.030 1686.840 1786.570 1686.980 ;
        RECT 1783.030 1686.780 1783.350 1686.840 ;
        RECT 1786.250 1686.780 1786.570 1686.840 ;
        RECT 1786.250 31.520 1786.570 31.580 ;
        RECT 2345.610 31.520 2345.930 31.580 ;
        RECT 1786.250 31.380 2345.930 31.520 ;
        RECT 1786.250 31.320 1786.570 31.380 ;
        RECT 2345.610 31.320 2345.930 31.380 ;
      LAYER via ;
        RECT 1783.060 1686.780 1783.320 1687.040 ;
        RECT 1786.280 1686.780 1786.540 1687.040 ;
        RECT 1786.280 31.320 1786.540 31.580 ;
        RECT 2345.640 31.320 2345.900 31.580 ;
      LAYER met2 ;
        RECT 1783.050 1700.000 1783.330 1704.000 ;
        RECT 1783.120 1687.070 1783.260 1700.000 ;
        RECT 1783.060 1686.750 1783.320 1687.070 ;
        RECT 1786.280 1686.750 1786.540 1687.070 ;
        RECT 1786.340 31.610 1786.480 1686.750 ;
        RECT 1786.280 31.290 1786.540 31.610 ;
        RECT 2345.640 31.290 2345.900 31.610 ;
        RECT 2345.700 2.400 2345.840 31.290 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1788.090 1686.640 1788.410 1686.700 ;
        RECT 1793.610 1686.640 1793.930 1686.700 ;
        RECT 1788.090 1686.500 1793.930 1686.640 ;
        RECT 1788.090 1686.440 1788.410 1686.500 ;
        RECT 1793.610 1686.440 1793.930 1686.500 ;
        RECT 1793.610 31.180 1793.930 31.240 ;
        RECT 2363.550 31.180 2363.870 31.240 ;
        RECT 1793.610 31.040 2363.870 31.180 ;
        RECT 1793.610 30.980 1793.930 31.040 ;
        RECT 2363.550 30.980 2363.870 31.040 ;
      LAYER via ;
        RECT 1788.120 1686.440 1788.380 1686.700 ;
        RECT 1793.640 1686.440 1793.900 1686.700 ;
        RECT 1793.640 30.980 1793.900 31.240 ;
        RECT 2363.580 30.980 2363.840 31.240 ;
      LAYER met2 ;
        RECT 1788.110 1700.000 1788.390 1704.000 ;
        RECT 1788.180 1686.730 1788.320 1700.000 ;
        RECT 1788.120 1686.410 1788.380 1686.730 ;
        RECT 1793.640 1686.410 1793.900 1686.730 ;
        RECT 1793.700 31.270 1793.840 1686.410 ;
        RECT 1793.640 30.950 1793.900 31.270 ;
        RECT 2363.580 30.950 2363.840 31.270 ;
        RECT 2363.640 2.400 2363.780 30.950 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1793.150 30.840 1793.470 30.900 ;
        RECT 2381.490 30.840 2381.810 30.900 ;
        RECT 1793.150 30.700 2381.810 30.840 ;
        RECT 1793.150 30.640 1793.470 30.700 ;
        RECT 2381.490 30.640 2381.810 30.700 ;
      LAYER via ;
        RECT 1793.180 30.640 1793.440 30.900 ;
        RECT 2381.520 30.640 2381.780 30.900 ;
      LAYER met2 ;
        RECT 1792.710 1700.410 1792.990 1704.000 ;
        RECT 1792.710 1700.270 1793.380 1700.410 ;
        RECT 1792.710 1700.000 1792.990 1700.270 ;
        RECT 1793.240 30.930 1793.380 1700.270 ;
        RECT 1793.180 30.610 1793.440 30.930 ;
        RECT 2381.520 30.610 2381.780 30.930 ;
        RECT 2381.580 2.400 2381.720 30.610 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 0.300 ;
=======
      LAYER met1 ;
        RECT 1797.750 1689.020 1798.070 1689.080 ;
        RECT 1800.050 1689.020 1800.370 1689.080 ;
        RECT 1797.750 1688.880 1800.370 1689.020 ;
        RECT 1797.750 1688.820 1798.070 1688.880 ;
        RECT 1800.050 1688.820 1800.370 1688.880 ;
      LAYER via ;
        RECT 1797.780 1688.820 1798.040 1689.080 ;
        RECT 1800.080 1688.820 1800.340 1689.080 ;
      LAYER met2 ;
        RECT 1797.770 1700.000 1798.050 1704.000 ;
        RECT 1797.840 1689.110 1797.980 1700.000 ;
        RECT 1797.780 1688.790 1798.040 1689.110 ;
        RECT 1800.080 1688.790 1800.340 1689.110 ;
        RECT 1800.140 33.845 1800.280 1688.790 ;
        RECT 1800.070 33.475 1800.350 33.845 ;
        RECT 2399.450 33.475 2399.730 33.845 ;
        RECT 2399.520 2.400 2399.660 33.475 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
      LAYER via2 ;
        RECT 1800.070 33.520 1800.350 33.800 ;
        RECT 2399.450 33.520 2399.730 33.800 ;
      LAYER met3 ;
        RECT 1800.045 33.810 1800.375 33.825 ;
        RECT 2399.425 33.810 2399.755 33.825 ;
        RECT 1800.045 33.510 2399.755 33.810 ;
        RECT 1800.045 33.495 1800.375 33.510 ;
        RECT 2399.425 33.495 2399.755 33.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 0.300 ;
=======
      LAYER li1 ;
        RECT 1360.825 1545.725 1360.995 1593.835 ;
        RECT 1360.825 1400.885 1360.995 1448.995 ;
        RECT 1360.825 1207.425 1360.995 1255.875 ;
        RECT 1360.825 1062.585 1360.995 1110.695 ;
        RECT 1360.825 821.185 1360.995 910.775 ;
        RECT 1361.285 517.565 1361.455 565.675 ;
      LAYER mcon ;
        RECT 1360.825 1593.665 1360.995 1593.835 ;
        RECT 1360.825 1448.825 1360.995 1448.995 ;
        RECT 1360.825 1255.705 1360.995 1255.875 ;
        RECT 1360.825 1110.525 1360.995 1110.695 ;
        RECT 1360.825 910.605 1360.995 910.775 ;
        RECT 1361.285 565.505 1361.455 565.675 ;
      LAYER met1 ;
        RECT 1360.750 1593.820 1361.070 1593.880 ;
        RECT 1360.555 1593.680 1361.070 1593.820 ;
        RECT 1360.750 1593.620 1361.070 1593.680 ;
        RECT 1360.765 1545.880 1361.055 1545.925 ;
        RECT 1361.210 1545.880 1361.530 1545.940 ;
        RECT 1360.765 1545.740 1361.530 1545.880 ;
        RECT 1360.765 1545.695 1361.055 1545.740 ;
        RECT 1361.210 1545.680 1361.530 1545.740 ;
        RECT 1360.765 1448.980 1361.055 1449.025 ;
        RECT 1361.210 1448.980 1361.530 1449.040 ;
        RECT 1360.765 1448.840 1361.530 1448.980 ;
        RECT 1360.765 1448.795 1361.055 1448.840 ;
        RECT 1361.210 1448.780 1361.530 1448.840 ;
        RECT 1360.750 1401.040 1361.070 1401.100 ;
        RECT 1360.555 1400.900 1361.070 1401.040 ;
        RECT 1360.750 1400.840 1361.070 1400.900 ;
        RECT 1361.210 1304.820 1361.530 1304.880 ;
        RECT 1360.840 1304.680 1361.530 1304.820 ;
        RECT 1360.840 1304.540 1360.980 1304.680 ;
        RECT 1361.210 1304.620 1361.530 1304.680 ;
        RECT 1360.750 1304.280 1361.070 1304.540 ;
        RECT 1360.750 1255.860 1361.070 1255.920 ;
        RECT 1360.555 1255.720 1361.070 1255.860 ;
        RECT 1360.750 1255.660 1361.070 1255.720 ;
        RECT 1360.750 1207.580 1361.070 1207.640 ;
        RECT 1360.555 1207.440 1361.070 1207.580 ;
        RECT 1360.750 1207.380 1361.070 1207.440 ;
        RECT 1360.750 1110.680 1361.070 1110.740 ;
        RECT 1360.555 1110.540 1361.070 1110.680 ;
        RECT 1360.750 1110.480 1361.070 1110.540 ;
        RECT 1360.765 1062.740 1361.055 1062.785 ;
        RECT 1361.210 1062.740 1361.530 1062.800 ;
        RECT 1360.765 1062.600 1361.530 1062.740 ;
        RECT 1360.765 1062.555 1361.055 1062.600 ;
        RECT 1361.210 1062.540 1361.530 1062.600 ;
        RECT 1360.750 918.240 1361.070 918.300 ;
        RECT 1361.210 918.240 1361.530 918.300 ;
        RECT 1360.750 918.100 1361.530 918.240 ;
        RECT 1360.750 918.040 1361.070 918.100 ;
        RECT 1361.210 918.040 1361.530 918.100 ;
        RECT 1360.750 910.760 1361.070 910.820 ;
        RECT 1360.555 910.620 1361.070 910.760 ;
        RECT 1360.750 910.560 1361.070 910.620 ;
        RECT 1360.750 821.340 1361.070 821.400 ;
        RECT 1360.555 821.200 1361.070 821.340 ;
        RECT 1360.750 821.140 1361.070 821.200 ;
        RECT 1358.910 814.200 1359.230 814.260 ;
        RECT 1360.750 814.200 1361.070 814.260 ;
        RECT 1358.910 814.060 1361.070 814.200 ;
        RECT 1358.910 814.000 1359.230 814.060 ;
        RECT 1360.750 814.000 1361.070 814.060 ;
        RECT 1360.750 765.920 1361.070 765.980 ;
        RECT 1361.670 765.920 1361.990 765.980 ;
        RECT 1360.750 765.780 1361.990 765.920 ;
        RECT 1360.750 765.720 1361.070 765.780 ;
        RECT 1361.670 765.720 1361.990 765.780 ;
        RECT 1358.910 717.640 1359.230 717.700 ;
        RECT 1360.750 717.640 1361.070 717.700 ;
        RECT 1358.910 717.500 1361.070 717.640 ;
        RECT 1358.910 717.440 1359.230 717.500 ;
        RECT 1360.750 717.440 1361.070 717.500 ;
        RECT 1361.225 565.660 1361.515 565.705 ;
        RECT 1361.670 565.660 1361.990 565.720 ;
        RECT 1361.225 565.520 1361.990 565.660 ;
        RECT 1361.225 565.475 1361.515 565.520 ;
        RECT 1361.670 565.460 1361.990 565.520 ;
        RECT 1361.210 517.720 1361.530 517.780 ;
        RECT 1361.015 517.580 1361.530 517.720 ;
        RECT 1361.210 517.520 1361.530 517.580 ;
        RECT 1360.750 427.960 1361.070 428.020 ;
        RECT 1361.210 427.960 1361.530 428.020 ;
        RECT 1360.750 427.820 1361.530 427.960 ;
        RECT 1360.750 427.760 1361.070 427.820 ;
        RECT 1361.210 427.760 1361.530 427.820 ;
        RECT 1360.750 283.120 1361.070 283.180 ;
        RECT 1361.210 283.120 1361.530 283.180 ;
        RECT 1360.750 282.980 1361.530 283.120 ;
        RECT 1360.750 282.920 1361.070 282.980 ;
        RECT 1361.210 282.920 1361.530 282.980 ;
        RECT 800.010 50.900 800.330 50.960 ;
        RECT 1361.210 50.900 1361.530 50.960 ;
        RECT 800.010 50.760 1361.530 50.900 ;
        RECT 800.010 50.700 800.330 50.760 ;
        RECT 1361.210 50.700 1361.530 50.760 ;
        RECT 793.570 20.980 793.890 21.040 ;
        RECT 800.010 20.980 800.330 21.040 ;
        RECT 793.570 20.840 800.330 20.980 ;
        RECT 793.570 20.780 793.890 20.840 ;
        RECT 800.010 20.780 800.330 20.840 ;
      LAYER via ;
        RECT 1360.780 1593.620 1361.040 1593.880 ;
        RECT 1361.240 1545.680 1361.500 1545.940 ;
        RECT 1361.240 1448.780 1361.500 1449.040 ;
        RECT 1360.780 1400.840 1361.040 1401.100 ;
        RECT 1361.240 1304.620 1361.500 1304.880 ;
        RECT 1360.780 1304.280 1361.040 1304.540 ;
        RECT 1360.780 1255.660 1361.040 1255.920 ;
        RECT 1360.780 1207.380 1361.040 1207.640 ;
        RECT 1360.780 1110.480 1361.040 1110.740 ;
        RECT 1361.240 1062.540 1361.500 1062.800 ;
        RECT 1360.780 918.040 1361.040 918.300 ;
        RECT 1361.240 918.040 1361.500 918.300 ;
        RECT 1360.780 910.560 1361.040 910.820 ;
        RECT 1360.780 821.140 1361.040 821.400 ;
        RECT 1358.940 814.000 1359.200 814.260 ;
        RECT 1360.780 814.000 1361.040 814.260 ;
        RECT 1360.780 765.720 1361.040 765.980 ;
        RECT 1361.700 765.720 1361.960 765.980 ;
        RECT 1358.940 717.440 1359.200 717.700 ;
        RECT 1360.780 717.440 1361.040 717.700 ;
        RECT 1361.700 565.460 1361.960 565.720 ;
        RECT 1361.240 517.520 1361.500 517.780 ;
        RECT 1360.780 427.760 1361.040 428.020 ;
        RECT 1361.240 427.760 1361.500 428.020 ;
        RECT 1360.780 282.920 1361.040 283.180 ;
        RECT 1361.240 282.920 1361.500 283.180 ;
        RECT 800.040 50.700 800.300 50.960 ;
        RECT 1361.240 50.700 1361.500 50.960 ;
        RECT 793.600 20.780 793.860 21.040 ;
        RECT 800.040 20.780 800.300 21.040 ;
      LAYER met2 ;
        RECT 1363.990 1700.410 1364.270 1704.000 ;
        RECT 1363.140 1700.270 1364.270 1700.410 ;
        RECT 1363.140 1677.290 1363.280 1700.270 ;
        RECT 1363.990 1700.000 1364.270 1700.270 ;
        RECT 1360.840 1677.150 1363.280 1677.290 ;
        RECT 1360.840 1593.910 1360.980 1677.150 ;
        RECT 1360.780 1593.590 1361.040 1593.910 ;
        RECT 1361.240 1545.650 1361.500 1545.970 ;
        RECT 1361.300 1449.070 1361.440 1545.650 ;
        RECT 1361.240 1448.750 1361.500 1449.070 ;
        RECT 1360.780 1400.810 1361.040 1401.130 ;
        RECT 1360.840 1352.250 1360.980 1400.810 ;
        RECT 1360.840 1352.110 1361.440 1352.250 ;
        RECT 1361.300 1304.910 1361.440 1352.110 ;
        RECT 1361.240 1304.590 1361.500 1304.910 ;
        RECT 1360.780 1304.250 1361.040 1304.570 ;
        RECT 1360.840 1255.950 1360.980 1304.250 ;
        RECT 1360.780 1255.630 1361.040 1255.950 ;
        RECT 1360.780 1207.350 1361.040 1207.670 ;
        RECT 1360.840 1110.770 1360.980 1207.350 ;
        RECT 1360.780 1110.450 1361.040 1110.770 ;
        RECT 1361.240 1062.510 1361.500 1062.830 ;
        RECT 1361.300 918.330 1361.440 1062.510 ;
        RECT 1360.780 918.010 1361.040 918.330 ;
        RECT 1361.240 918.010 1361.500 918.330 ;
        RECT 1360.840 910.850 1360.980 918.010 ;
        RECT 1360.780 910.530 1361.040 910.850 ;
        RECT 1360.780 821.110 1361.040 821.430 ;
        RECT 1360.840 814.290 1360.980 821.110 ;
        RECT 1358.940 813.970 1359.200 814.290 ;
        RECT 1360.780 813.970 1361.040 814.290 ;
        RECT 1359.000 766.205 1359.140 813.970 ;
        RECT 1358.930 765.835 1359.210 766.205 ;
        RECT 1360.770 765.835 1361.050 766.205 ;
        RECT 1360.780 765.690 1361.040 765.835 ;
        RECT 1361.700 765.690 1361.960 766.010 ;
        RECT 1361.760 717.925 1361.900 765.690 ;
        RECT 1358.940 717.410 1359.200 717.730 ;
        RECT 1360.770 717.555 1361.050 717.925 ;
        RECT 1361.690 717.555 1361.970 717.925 ;
        RECT 1360.780 717.410 1361.040 717.555 ;
        RECT 1359.000 669.645 1359.140 717.410 ;
        RECT 1358.930 669.275 1359.210 669.645 ;
        RECT 1360.770 669.275 1361.050 669.645 ;
        RECT 1360.840 589.970 1360.980 669.275 ;
        RECT 1360.840 589.830 1361.440 589.970 ;
        RECT 1361.300 566.170 1361.440 589.830 ;
        RECT 1361.300 566.030 1361.900 566.170 ;
        RECT 1361.760 565.750 1361.900 566.030 ;
        RECT 1361.700 565.430 1361.960 565.750 ;
        RECT 1361.240 517.490 1361.500 517.810 ;
        RECT 1361.300 517.210 1361.440 517.490 ;
        RECT 1360.840 517.070 1361.440 517.210 ;
        RECT 1360.840 470.405 1360.980 517.070 ;
        RECT 1360.770 470.035 1361.050 470.405 ;
        RECT 1361.230 469.355 1361.510 469.725 ;
        RECT 1361.300 428.050 1361.440 469.355 ;
        RECT 1360.780 427.730 1361.040 428.050 ;
        RECT 1361.240 427.730 1361.500 428.050 ;
        RECT 1360.840 283.210 1360.980 427.730 ;
        RECT 1360.780 282.890 1361.040 283.210 ;
        RECT 1361.240 282.890 1361.500 283.210 ;
        RECT 1361.300 207.810 1361.440 282.890 ;
        RECT 1361.300 207.670 1361.900 207.810 ;
        RECT 1361.760 206.450 1361.900 207.670 ;
        RECT 1360.840 206.310 1361.900 206.450 ;
        RECT 1360.840 144.685 1360.980 206.310 ;
        RECT 1360.770 144.315 1361.050 144.685 ;
        RECT 1361.230 143.635 1361.510 144.005 ;
        RECT 1361.300 50.990 1361.440 143.635 ;
        RECT 800.040 50.670 800.300 50.990 ;
        RECT 1361.240 50.670 1361.500 50.990 ;
        RECT 800.100 21.070 800.240 50.670 ;
        RECT 793.600 20.750 793.860 21.070 ;
        RECT 800.040 20.750 800.300 21.070 ;
        RECT 793.660 2.400 793.800 20.750 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 1358.930 765.880 1359.210 766.160 ;
        RECT 1360.770 765.880 1361.050 766.160 ;
        RECT 1360.770 717.600 1361.050 717.880 ;
        RECT 1361.690 717.600 1361.970 717.880 ;
        RECT 1358.930 669.320 1359.210 669.600 ;
        RECT 1360.770 669.320 1361.050 669.600 ;
        RECT 1360.770 470.080 1361.050 470.360 ;
        RECT 1361.230 469.400 1361.510 469.680 ;
        RECT 1360.770 144.360 1361.050 144.640 ;
        RECT 1361.230 143.680 1361.510 143.960 ;
      LAYER met3 ;
        RECT 1358.905 766.170 1359.235 766.185 ;
        RECT 1360.745 766.170 1361.075 766.185 ;
        RECT 1358.905 765.870 1361.075 766.170 ;
        RECT 1358.905 765.855 1359.235 765.870 ;
        RECT 1360.745 765.855 1361.075 765.870 ;
        RECT 1360.745 717.890 1361.075 717.905 ;
        RECT 1361.665 717.890 1361.995 717.905 ;
        RECT 1360.745 717.590 1361.995 717.890 ;
        RECT 1360.745 717.575 1361.075 717.590 ;
        RECT 1361.665 717.575 1361.995 717.590 ;
        RECT 1358.905 669.610 1359.235 669.625 ;
        RECT 1360.745 669.610 1361.075 669.625 ;
        RECT 1358.905 669.310 1361.075 669.610 ;
        RECT 1358.905 669.295 1359.235 669.310 ;
        RECT 1360.745 669.295 1361.075 669.310 ;
        RECT 1360.745 470.370 1361.075 470.385 ;
        RECT 1360.745 470.070 1362.210 470.370 ;
        RECT 1360.745 470.055 1361.075 470.070 ;
        RECT 1361.205 469.690 1361.535 469.705 ;
        RECT 1361.910 469.690 1362.210 470.070 ;
        RECT 1361.205 469.390 1362.210 469.690 ;
        RECT 1361.205 469.375 1361.535 469.390 ;
        RECT 1360.745 144.650 1361.075 144.665 ;
        RECT 1360.070 144.350 1361.075 144.650 ;
        RECT 1360.070 143.970 1360.370 144.350 ;
        RECT 1360.745 144.335 1361.075 144.350 ;
        RECT 1361.205 143.970 1361.535 143.985 ;
        RECT 1360.070 143.670 1361.535 143.970 ;
        RECT 1361.205 143.655 1361.535 143.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1318.430 1678.140 1318.750 1678.200 ;
        RECT 1321.190 1678.140 1321.510 1678.200 ;
        RECT 1318.430 1678.000 1321.510 1678.140 ;
        RECT 1318.430 1677.940 1318.750 1678.000 ;
        RECT 1321.190 1677.940 1321.510 1678.000 ;
      LAYER via ;
        RECT 1318.460 1677.940 1318.720 1678.200 ;
        RECT 1321.220 1677.940 1321.480 1678.200 ;
      LAYER met2 ;
        RECT 1322.130 1700.410 1322.410 1704.000 ;
        RECT 1321.280 1700.270 1322.410 1700.410 ;
        RECT 1321.280 1678.230 1321.420 1700.270 ;
        RECT 1322.130 1700.000 1322.410 1700.270 ;
        RECT 1318.460 1677.910 1318.720 1678.230 ;
        RECT 1321.220 1677.910 1321.480 1678.230 ;
        RECT 1318.520 33.165 1318.660 1677.910 ;
        RECT 639.030 32.795 639.310 33.165 ;
        RECT 1318.450 32.795 1318.730 33.165 ;
        RECT 639.100 2.400 639.240 32.795 ;
        RECT 638.890 -4.800 639.450 2.400 ;
      LAYER via2 ;
        RECT 639.030 32.840 639.310 33.120 ;
        RECT 1318.450 32.840 1318.730 33.120 ;
      LAYER met3 ;
        RECT 639.005 33.130 639.335 33.145 ;
        RECT 1318.425 33.130 1318.755 33.145 ;
        RECT 639.005 32.830 1318.755 33.130 ;
        RECT 639.005 32.815 639.335 32.830 ;
        RECT 1318.425 32.815 1318.755 32.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1804.190 1684.260 1804.510 1684.320 ;
        RECT 1807.410 1684.260 1807.730 1684.320 ;
        RECT 1804.190 1684.120 1807.730 1684.260 ;
        RECT 1804.190 1684.060 1804.510 1684.120 ;
        RECT 1807.410 1684.060 1807.730 1684.120 ;
      LAYER via ;
        RECT 1804.220 1684.060 1804.480 1684.320 ;
        RECT 1807.440 1684.060 1807.700 1684.320 ;
      LAYER met2 ;
        RECT 1804.210 1700.000 1804.490 1704.000 ;
        RECT 1804.280 1684.350 1804.420 1700.000 ;
        RECT 1804.220 1684.030 1804.480 1684.350 ;
        RECT 1807.440 1684.030 1807.700 1684.350 ;
        RECT 1807.500 33.165 1807.640 1684.030 ;
        RECT 1807.430 32.795 1807.710 33.165 ;
        RECT 2422.910 32.795 2423.190 33.165 ;
        RECT 2422.980 2.400 2423.120 32.795 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
      LAYER via2 ;
        RECT 1807.430 32.840 1807.710 33.120 ;
        RECT 2422.910 32.840 2423.190 33.120 ;
      LAYER met3 ;
        RECT 1807.405 33.130 1807.735 33.145 ;
        RECT 2422.885 33.130 2423.215 33.145 ;
        RECT 1807.405 32.830 2423.215 33.130 ;
        RECT 1807.405 32.815 1807.735 32.830 ;
        RECT 2422.885 32.815 2423.215 32.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1808.790 1683.920 1809.110 1683.980 ;
        RECT 1814.310 1683.920 1814.630 1683.980 ;
        RECT 1808.790 1683.780 1814.630 1683.920 ;
        RECT 1808.790 1683.720 1809.110 1683.780 ;
        RECT 1814.310 1683.720 1814.630 1683.780 ;
      LAYER via ;
        RECT 1808.820 1683.720 1809.080 1683.980 ;
        RECT 1814.340 1683.720 1814.600 1683.980 ;
      LAYER met2 ;
        RECT 1808.810 1700.000 1809.090 1704.000 ;
        RECT 1808.880 1684.010 1809.020 1700.000 ;
        RECT 1808.820 1683.690 1809.080 1684.010 ;
        RECT 1814.340 1683.690 1814.600 1684.010 ;
        RECT 1814.400 32.485 1814.540 1683.690 ;
        RECT 1814.330 32.115 1814.610 32.485 ;
        RECT 2440.850 32.115 2441.130 32.485 ;
        RECT 2440.920 2.400 2441.060 32.115 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
      LAYER via2 ;
        RECT 1814.330 32.160 1814.610 32.440 ;
        RECT 2440.850 32.160 2441.130 32.440 ;
      LAYER met3 ;
        RECT 1814.305 32.450 1814.635 32.465 ;
        RECT 2440.825 32.450 2441.155 32.465 ;
        RECT 1814.305 32.150 2441.155 32.450 ;
        RECT 1814.305 32.135 1814.635 32.150 ;
        RECT 2440.825 32.135 2441.155 32.150 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2458.650 -4.800 2459.210 0.300 ;
=======
        RECT 1813.870 1700.000 1814.150 1704.000 ;
        RECT 1813.940 31.805 1814.080 1700.000 ;
        RECT 1813.870 31.435 1814.150 31.805 ;
        RECT 2458.790 31.435 2459.070 31.805 ;
        RECT 2458.860 2.400 2459.000 31.435 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
      LAYER via2 ;
        RECT 1813.870 31.480 1814.150 31.760 ;
        RECT 2458.790 31.480 2459.070 31.760 ;
      LAYER met3 ;
        RECT 1813.845 31.770 1814.175 31.785 ;
        RECT 2458.765 31.770 2459.095 31.785 ;
        RECT 1813.845 31.470 2459.095 31.770 ;
        RECT 1813.845 31.455 1814.175 31.470 ;
        RECT 2458.765 31.455 2459.095 31.470 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2476.590 -4.800 2477.150 0.300 ;
=======
        RECT 1818.470 1700.410 1818.750 1704.000 ;
        RECT 1818.470 1700.270 1820.060 1700.410 ;
        RECT 1818.470 1700.000 1818.750 1700.270 ;
        RECT 1819.920 1670.490 1820.060 1700.270 ;
        RECT 1819.920 1670.350 1820.520 1670.490 ;
        RECT 1820.380 31.125 1820.520 1670.350 ;
        RECT 1820.310 30.755 1820.590 31.125 ;
        RECT 2476.730 30.755 2477.010 31.125 ;
        RECT 2476.800 2.400 2476.940 30.755 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
      LAYER via2 ;
        RECT 1820.310 30.800 1820.590 31.080 ;
        RECT 2476.730 30.800 2477.010 31.080 ;
      LAYER met3 ;
        RECT 1820.285 31.090 1820.615 31.105 ;
        RECT 2476.705 31.090 2477.035 31.105 ;
        RECT 1820.285 30.790 2477.035 31.090 ;
        RECT 1820.285 30.775 1820.615 30.790 ;
        RECT 2476.705 30.775 2477.035 30.790 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1823.510 1683.920 1823.830 1683.980 ;
        RECT 1826.270 1683.920 1826.590 1683.980 ;
        RECT 1823.510 1683.780 1826.590 1683.920 ;
        RECT 1823.510 1683.720 1823.830 1683.780 ;
        RECT 1826.270 1683.720 1826.590 1683.780 ;
      LAYER via ;
        RECT 1823.540 1683.720 1823.800 1683.980 ;
        RECT 1826.300 1683.720 1826.560 1683.980 ;
      LAYER met2 ;
        RECT 1823.530 1700.000 1823.810 1704.000 ;
        RECT 1823.600 1684.010 1823.740 1700.000 ;
        RECT 1823.540 1683.690 1823.800 1684.010 ;
        RECT 1826.300 1683.690 1826.560 1684.010 ;
        RECT 1826.360 46.765 1826.500 1683.690 ;
        RECT 1826.290 46.395 1826.570 46.765 ;
        RECT 2494.670 46.395 2494.950 46.765 ;
        RECT 2494.740 2.400 2494.880 46.395 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
      LAYER via2 ;
        RECT 1826.290 46.440 1826.570 46.720 ;
        RECT 2494.670 46.440 2494.950 46.720 ;
      LAYER met3 ;
        RECT 1826.265 46.730 1826.595 46.745 ;
        RECT 2494.645 46.730 2494.975 46.745 ;
        RECT 1826.265 46.430 2494.975 46.730 ;
        RECT 1826.265 46.415 1826.595 46.430 ;
        RECT 2494.645 46.415 2494.975 46.430 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1826.730 1683.920 1827.050 1683.980 ;
        RECT 1828.110 1683.920 1828.430 1683.980 ;
        RECT 1826.730 1683.780 1828.430 1683.920 ;
        RECT 1826.730 1683.720 1827.050 1683.780 ;
        RECT 1828.110 1683.720 1828.430 1683.780 ;
      LAYER via ;
        RECT 1826.760 1683.720 1827.020 1683.980 ;
        RECT 1828.140 1683.720 1828.400 1683.980 ;
      LAYER met2 ;
        RECT 1828.130 1700.000 1828.410 1704.000 ;
        RECT 1828.200 1684.010 1828.340 1700.000 ;
        RECT 1826.760 1683.690 1827.020 1684.010 ;
        RECT 1828.140 1683.690 1828.400 1684.010 ;
        RECT 1826.820 46.085 1826.960 1683.690 ;
        RECT 1826.750 45.715 1827.030 46.085 ;
        RECT 2512.150 45.715 2512.430 46.085 ;
        RECT 2512.220 2.400 2512.360 45.715 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
      LAYER via2 ;
        RECT 1826.750 45.760 1827.030 46.040 ;
        RECT 2512.150 45.760 2512.430 46.040 ;
      LAYER met3 ;
        RECT 1826.725 46.050 1827.055 46.065 ;
        RECT 2512.125 46.050 2512.455 46.065 ;
        RECT 1826.725 45.750 2512.455 46.050 ;
        RECT 1826.725 45.735 1827.055 45.750 ;
        RECT 2512.125 45.735 2512.455 45.750 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 0.300 ;
=======
      LAYER met1 ;
        RECT 1832.710 110.400 1833.030 110.460 ;
        RECT 1834.090 110.400 1834.410 110.460 ;
        RECT 1832.710 110.260 1834.410 110.400 ;
        RECT 1832.710 110.200 1833.030 110.260 ;
        RECT 1834.090 110.200 1834.410 110.260 ;
      LAYER via ;
        RECT 1832.740 110.200 1833.000 110.460 ;
        RECT 1834.120 110.200 1834.380 110.460 ;
      LAYER met2 ;
        RECT 1833.190 1700.410 1833.470 1704.000 ;
        RECT 1833.190 1700.270 1834.320 1700.410 ;
        RECT 1833.190 1700.000 1833.470 1700.270 ;
        RECT 1834.180 110.490 1834.320 1700.270 ;
        RECT 1832.740 110.170 1833.000 110.490 ;
        RECT 1834.120 110.170 1834.380 110.490 ;
        RECT 1832.800 45.405 1832.940 110.170 ;
        RECT 1832.730 45.035 1833.010 45.405 ;
        RECT 2530.090 45.035 2530.370 45.405 ;
        RECT 2530.160 2.400 2530.300 45.035 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
      LAYER via2 ;
        RECT 1832.730 45.080 1833.010 45.360 ;
        RECT 2530.090 45.080 2530.370 45.360 ;
      LAYER met3 ;
        RECT 1832.705 45.370 1833.035 45.385 ;
        RECT 2530.065 45.370 2530.395 45.385 ;
        RECT 1832.705 45.070 2530.395 45.370 ;
        RECT 1832.705 45.055 1833.035 45.070 ;
        RECT 2530.065 45.055 2530.395 45.070 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1837.770 1684.600 1838.090 1684.660 ;
        RECT 1840.990 1684.600 1841.310 1684.660 ;
        RECT 1837.770 1684.460 1841.310 1684.600 ;
        RECT 1837.770 1684.400 1838.090 1684.460 ;
        RECT 1840.990 1684.400 1841.310 1684.460 ;
        RECT 1840.990 36.620 1841.310 36.680 ;
        RECT 2548.010 36.620 2548.330 36.680 ;
        RECT 1840.990 36.480 2548.330 36.620 ;
        RECT 1840.990 36.420 1841.310 36.480 ;
        RECT 2548.010 36.420 2548.330 36.480 ;
      LAYER via ;
        RECT 1837.800 1684.400 1838.060 1684.660 ;
        RECT 1841.020 1684.400 1841.280 1684.660 ;
        RECT 1841.020 36.420 1841.280 36.680 ;
        RECT 2548.040 36.420 2548.300 36.680 ;
      LAYER met2 ;
        RECT 1837.790 1700.000 1838.070 1704.000 ;
        RECT 1837.860 1684.690 1838.000 1700.000 ;
        RECT 1837.800 1684.370 1838.060 1684.690 ;
        RECT 1841.020 1684.370 1841.280 1684.690 ;
        RECT 1841.080 36.710 1841.220 1684.370 ;
        RECT 1841.020 36.390 1841.280 36.710 ;
        RECT 2548.040 36.390 2548.300 36.710 ;
        RECT 2548.100 2.400 2548.240 36.390 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1842.830 1683.920 1843.150 1683.980 ;
        RECT 1848.350 1683.920 1848.670 1683.980 ;
        RECT 1842.830 1683.780 1848.670 1683.920 ;
        RECT 1842.830 1683.720 1843.150 1683.780 ;
        RECT 1848.350 1683.720 1848.670 1683.780 ;
        RECT 1848.350 36.960 1848.670 37.020 ;
        RECT 2565.950 36.960 2566.270 37.020 ;
        RECT 1848.350 36.820 2566.270 36.960 ;
        RECT 1848.350 36.760 1848.670 36.820 ;
        RECT 2565.950 36.760 2566.270 36.820 ;
      LAYER via ;
        RECT 1842.860 1683.720 1843.120 1683.980 ;
        RECT 1848.380 1683.720 1848.640 1683.980 ;
        RECT 1848.380 36.760 1848.640 37.020 ;
        RECT 2565.980 36.760 2566.240 37.020 ;
      LAYER met2 ;
        RECT 1842.850 1700.000 1843.130 1704.000 ;
        RECT 1842.920 1684.010 1843.060 1700.000 ;
        RECT 1842.860 1683.690 1843.120 1684.010 ;
        RECT 1848.380 1683.690 1848.640 1684.010 ;
        RECT 1848.440 37.050 1848.580 1683.690 ;
        RECT 1848.380 36.730 1848.640 37.050 ;
        RECT 2565.980 36.730 2566.240 37.050 ;
        RECT 2566.040 2.400 2566.180 36.730 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1847.890 37.300 1848.210 37.360 ;
        RECT 2583.890 37.300 2584.210 37.360 ;
        RECT 1847.890 37.160 2584.210 37.300 ;
        RECT 1847.890 37.100 1848.210 37.160 ;
        RECT 2583.890 37.100 2584.210 37.160 ;
      LAYER via ;
        RECT 1847.920 37.100 1848.180 37.360 ;
        RECT 2583.920 37.100 2584.180 37.360 ;
      LAYER met2 ;
        RECT 1847.450 1700.410 1847.730 1704.000 ;
        RECT 1847.450 1700.270 1848.120 1700.410 ;
        RECT 1847.450 1700.000 1847.730 1700.270 ;
        RECT 1847.980 37.390 1848.120 1700.270 ;
        RECT 1847.920 37.070 1848.180 37.390 ;
        RECT 2583.920 37.070 2584.180 37.390 ;
        RECT 2583.980 2.400 2584.120 37.070 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1366.270 1678.140 1366.590 1678.200 ;
        RECT 1369.030 1678.140 1369.350 1678.200 ;
        RECT 1366.270 1678.000 1369.350 1678.140 ;
        RECT 1366.270 1677.940 1366.590 1678.000 ;
        RECT 1369.030 1677.940 1369.350 1678.000 ;
        RECT 817.490 31.860 817.810 31.920 ;
        RECT 1366.270 31.860 1366.590 31.920 ;
        RECT 817.490 31.720 1366.590 31.860 ;
        RECT 817.490 31.660 817.810 31.720 ;
        RECT 1366.270 31.660 1366.590 31.720 ;
      LAYER via ;
        RECT 1366.300 1677.940 1366.560 1678.200 ;
        RECT 1369.060 1677.940 1369.320 1678.200 ;
        RECT 817.520 31.660 817.780 31.920 ;
        RECT 1366.300 31.660 1366.560 31.920 ;
      LAYER met2 ;
        RECT 1370.430 1700.410 1370.710 1704.000 ;
        RECT 1369.120 1700.270 1370.710 1700.410 ;
        RECT 1369.120 1678.230 1369.260 1700.270 ;
        RECT 1370.430 1700.000 1370.710 1700.270 ;
        RECT 1366.300 1677.910 1366.560 1678.230 ;
        RECT 1369.060 1677.910 1369.320 1678.230 ;
        RECT 1366.360 31.950 1366.500 1677.910 ;
        RECT 817.520 31.630 817.780 31.950 ;
        RECT 1366.300 31.630 1366.560 31.950 ;
        RECT 817.580 2.400 817.720 31.630 ;
        RECT 817.370 -4.800 817.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1852.030 1685.960 1852.350 1686.020 ;
        RECT 1854.330 1685.960 1854.650 1686.020 ;
        RECT 1852.030 1685.820 1854.650 1685.960 ;
        RECT 1852.030 1685.760 1852.350 1685.820 ;
        RECT 1854.330 1685.760 1854.650 1685.820 ;
        RECT 1854.330 37.640 1854.650 37.700 ;
        RECT 2601.370 37.640 2601.690 37.700 ;
        RECT 1854.330 37.500 2601.690 37.640 ;
        RECT 1854.330 37.440 1854.650 37.500 ;
        RECT 2601.370 37.440 2601.690 37.500 ;
      LAYER via ;
        RECT 1852.060 1685.760 1852.320 1686.020 ;
        RECT 1854.360 1685.760 1854.620 1686.020 ;
        RECT 1854.360 37.440 1854.620 37.700 ;
        RECT 2601.400 37.440 2601.660 37.700 ;
      LAYER met2 ;
        RECT 1852.050 1700.000 1852.330 1704.000 ;
        RECT 1852.120 1686.050 1852.260 1700.000 ;
        RECT 1852.060 1685.730 1852.320 1686.050 ;
        RECT 1854.360 1685.730 1854.620 1686.050 ;
        RECT 1854.420 37.730 1854.560 1685.730 ;
        RECT 1854.360 37.410 1854.620 37.730 ;
        RECT 2601.400 37.410 2601.660 37.730 ;
        RECT 2601.460 2.400 2601.600 37.410 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1857.090 1685.620 1857.410 1685.680 ;
        RECT 1861.690 1685.620 1862.010 1685.680 ;
        RECT 1857.090 1685.480 1862.010 1685.620 ;
        RECT 1857.090 1685.420 1857.410 1685.480 ;
        RECT 1861.690 1685.420 1862.010 1685.480 ;
        RECT 1861.690 41.380 1862.010 41.440 ;
        RECT 2619.310 41.380 2619.630 41.440 ;
        RECT 1861.690 41.240 2619.630 41.380 ;
        RECT 1861.690 41.180 1862.010 41.240 ;
        RECT 2619.310 41.180 2619.630 41.240 ;
      LAYER via ;
        RECT 1857.120 1685.420 1857.380 1685.680 ;
        RECT 1861.720 1685.420 1861.980 1685.680 ;
        RECT 1861.720 41.180 1861.980 41.440 ;
        RECT 2619.340 41.180 2619.600 41.440 ;
      LAYER met2 ;
        RECT 1857.110 1700.000 1857.390 1704.000 ;
        RECT 1857.180 1685.710 1857.320 1700.000 ;
        RECT 1857.120 1685.390 1857.380 1685.710 ;
        RECT 1861.720 1685.390 1861.980 1685.710 ;
        RECT 1861.780 41.470 1861.920 1685.390 ;
        RECT 1861.720 41.150 1861.980 41.470 ;
        RECT 2619.340 41.150 2619.600 41.470 ;
        RECT 2619.400 2.400 2619.540 41.150 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1862.150 41.040 1862.470 41.100 ;
        RECT 2637.250 41.040 2637.570 41.100 ;
        RECT 1862.150 40.900 2637.570 41.040 ;
        RECT 1862.150 40.840 1862.470 40.900 ;
        RECT 2637.250 40.840 2637.570 40.900 ;
      LAYER via ;
        RECT 1862.180 40.840 1862.440 41.100 ;
        RECT 2637.280 40.840 2637.540 41.100 ;
      LAYER met2 ;
        RECT 1861.710 1700.410 1861.990 1704.000 ;
        RECT 1861.710 1700.270 1862.380 1700.410 ;
        RECT 1861.710 1700.000 1861.990 1700.270 ;
        RECT 1862.240 41.130 1862.380 1700.270 ;
        RECT 1862.180 40.810 1862.440 41.130 ;
        RECT 2637.280 40.810 2637.540 41.130 ;
        RECT 2637.340 2.400 2637.480 40.810 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 0.300 ;
=======
      LAYER met1 ;
        RECT 1866.750 1684.600 1867.070 1684.660 ;
        RECT 1869.050 1684.600 1869.370 1684.660 ;
        RECT 1866.750 1684.460 1869.370 1684.600 ;
        RECT 1866.750 1684.400 1867.070 1684.460 ;
        RECT 1869.050 1684.400 1869.370 1684.460 ;
        RECT 1869.050 40.700 1869.370 40.760 ;
        RECT 2655.190 40.700 2655.510 40.760 ;
        RECT 1869.050 40.560 2655.510 40.700 ;
        RECT 1869.050 40.500 1869.370 40.560 ;
        RECT 2655.190 40.500 2655.510 40.560 ;
      LAYER via ;
        RECT 1866.780 1684.400 1867.040 1684.660 ;
        RECT 1869.080 1684.400 1869.340 1684.660 ;
        RECT 1869.080 40.500 1869.340 40.760 ;
        RECT 2655.220 40.500 2655.480 40.760 ;
      LAYER met2 ;
        RECT 1866.770 1700.000 1867.050 1704.000 ;
        RECT 1866.840 1684.690 1866.980 1700.000 ;
        RECT 1866.780 1684.370 1867.040 1684.690 ;
        RECT 1869.080 1684.370 1869.340 1684.690 ;
        RECT 1869.140 40.790 1869.280 1684.370 ;
        RECT 1869.080 40.470 1869.340 40.790 ;
        RECT 2655.220 40.470 2655.480 40.790 ;
        RECT 2655.280 2.400 2655.420 40.470 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1871.350 1686.640 1871.670 1686.700 ;
        RECT 1875.030 1686.640 1875.350 1686.700 ;
        RECT 1871.350 1686.500 1875.350 1686.640 ;
        RECT 1871.350 1686.440 1871.670 1686.500 ;
        RECT 1875.030 1686.440 1875.350 1686.500 ;
        RECT 1875.030 40.360 1875.350 40.420 ;
        RECT 2672.670 40.360 2672.990 40.420 ;
        RECT 1875.030 40.220 2672.990 40.360 ;
        RECT 1875.030 40.160 1875.350 40.220 ;
        RECT 2672.670 40.160 2672.990 40.220 ;
      LAYER via ;
        RECT 1871.380 1686.440 1871.640 1686.700 ;
        RECT 1875.060 1686.440 1875.320 1686.700 ;
        RECT 1875.060 40.160 1875.320 40.420 ;
        RECT 2672.700 40.160 2672.960 40.420 ;
      LAYER met2 ;
        RECT 1871.370 1700.000 1871.650 1704.000 ;
        RECT 1871.440 1686.730 1871.580 1700.000 ;
        RECT 1871.380 1686.410 1871.640 1686.730 ;
        RECT 1875.060 1686.410 1875.320 1686.730 ;
        RECT 1875.120 40.450 1875.260 1686.410 ;
        RECT 1875.060 40.130 1875.320 40.450 ;
        RECT 2672.700 40.130 2672.960 40.450 ;
        RECT 2672.760 2.400 2672.900 40.130 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1874.570 1685.620 1874.890 1685.680 ;
        RECT 1876.410 1685.620 1876.730 1685.680 ;
        RECT 1874.570 1685.480 1876.730 1685.620 ;
        RECT 1874.570 1685.420 1874.890 1685.480 ;
        RECT 1876.410 1685.420 1876.730 1685.480 ;
        RECT 1874.570 40.020 1874.890 40.080 ;
        RECT 2690.610 40.020 2690.930 40.080 ;
        RECT 1874.570 39.880 2690.930 40.020 ;
        RECT 1874.570 39.820 1874.890 39.880 ;
        RECT 2690.610 39.820 2690.930 39.880 ;
      LAYER via ;
        RECT 1874.600 1685.420 1874.860 1685.680 ;
        RECT 1876.440 1685.420 1876.700 1685.680 ;
        RECT 1874.600 39.820 1874.860 40.080 ;
        RECT 2690.640 39.820 2690.900 40.080 ;
      LAYER met2 ;
        RECT 1876.430 1700.000 1876.710 1704.000 ;
        RECT 1876.500 1685.710 1876.640 1700.000 ;
        RECT 1874.600 1685.390 1874.860 1685.710 ;
        RECT 1876.440 1685.390 1876.700 1685.710 ;
        RECT 1874.660 40.110 1874.800 1685.390 ;
        RECT 1874.600 39.790 1874.860 40.110 ;
        RECT 2690.640 39.790 2690.900 40.110 ;
        RECT 2690.700 2.400 2690.840 39.790 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1882.390 1608.920 1882.710 1609.180 ;
        RECT 1882.480 1608.160 1882.620 1608.920 ;
        RECT 1882.390 1607.900 1882.710 1608.160 ;
        RECT 1882.390 39.680 1882.710 39.740 ;
        RECT 2708.550 39.680 2708.870 39.740 ;
        RECT 1882.390 39.540 2708.870 39.680 ;
        RECT 1882.390 39.480 1882.710 39.540 ;
        RECT 2708.550 39.480 2708.870 39.540 ;
      LAYER via ;
        RECT 1882.420 1608.920 1882.680 1609.180 ;
        RECT 1882.420 1607.900 1882.680 1608.160 ;
        RECT 1882.420 39.480 1882.680 39.740 ;
        RECT 2708.580 39.480 2708.840 39.740 ;
      LAYER met2 ;
        RECT 1881.030 1700.410 1881.310 1704.000 ;
        RECT 1881.030 1700.270 1882.620 1700.410 ;
        RECT 1881.030 1700.000 1881.310 1700.270 ;
        RECT 1882.480 1609.210 1882.620 1700.270 ;
        RECT 1882.420 1608.890 1882.680 1609.210 ;
        RECT 1882.420 1607.870 1882.680 1608.190 ;
        RECT 1882.480 39.770 1882.620 1607.870 ;
        RECT 1882.420 39.450 1882.680 39.770 ;
        RECT 2708.580 39.450 2708.840 39.770 ;
        RECT 2708.640 2.400 2708.780 39.450 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1886.070 1686.640 1886.390 1686.700 ;
        RECT 1889.290 1686.640 1889.610 1686.700 ;
        RECT 1886.070 1686.500 1889.610 1686.640 ;
        RECT 1886.070 1686.440 1886.390 1686.500 ;
        RECT 1889.290 1686.440 1889.610 1686.500 ;
        RECT 1889.290 39.340 1889.610 39.400 ;
        RECT 2726.490 39.340 2726.810 39.400 ;
        RECT 1889.290 39.200 2726.810 39.340 ;
        RECT 1889.290 39.140 1889.610 39.200 ;
        RECT 2726.490 39.140 2726.810 39.200 ;
      LAYER via ;
        RECT 1886.100 1686.440 1886.360 1686.700 ;
        RECT 1889.320 1686.440 1889.580 1686.700 ;
        RECT 1889.320 39.140 1889.580 39.400 ;
        RECT 2726.520 39.140 2726.780 39.400 ;
      LAYER met2 ;
        RECT 1886.090 1700.000 1886.370 1704.000 ;
        RECT 1886.160 1686.730 1886.300 1700.000 ;
        RECT 1886.100 1686.410 1886.360 1686.730 ;
        RECT 1889.320 1686.410 1889.580 1686.730 ;
        RECT 1889.380 39.430 1889.520 1686.410 ;
        RECT 1889.320 39.110 1889.580 39.430 ;
        RECT 2726.520 39.110 2726.780 39.430 ;
        RECT 2726.580 2.400 2726.720 39.110 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 0.300 ;
=======
      LAYER met1 ;
        RECT 1890.670 1685.620 1890.990 1685.680 ;
        RECT 1896.190 1685.620 1896.510 1685.680 ;
        RECT 1890.670 1685.480 1896.510 1685.620 ;
        RECT 1890.670 1685.420 1890.990 1685.480 ;
        RECT 1896.190 1685.420 1896.510 1685.480 ;
        RECT 1896.190 39.000 1896.510 39.060 ;
        RECT 2744.430 39.000 2744.750 39.060 ;
        RECT 1896.190 38.860 2744.750 39.000 ;
        RECT 1896.190 38.800 1896.510 38.860 ;
        RECT 2744.430 38.800 2744.750 38.860 ;
      LAYER via ;
        RECT 1890.700 1685.420 1890.960 1685.680 ;
        RECT 1896.220 1685.420 1896.480 1685.680 ;
        RECT 1896.220 38.800 1896.480 39.060 ;
        RECT 2744.460 38.800 2744.720 39.060 ;
      LAYER met2 ;
        RECT 1890.690 1700.000 1890.970 1704.000 ;
        RECT 1890.760 1685.710 1890.900 1700.000 ;
        RECT 1890.700 1685.390 1890.960 1685.710 ;
        RECT 1896.220 1685.390 1896.480 1685.710 ;
        RECT 1896.280 39.090 1896.420 1685.390 ;
        RECT 1896.220 38.770 1896.480 39.090 ;
        RECT 2744.460 38.770 2744.720 39.090 ;
        RECT 2744.520 2.400 2744.660 38.770 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1892.050 1686.640 1892.370 1686.700 ;
        RECT 1895.730 1686.640 1896.050 1686.700 ;
        RECT 1892.050 1686.500 1896.050 1686.640 ;
        RECT 1892.050 1686.440 1892.370 1686.500 ;
        RECT 1895.730 1686.440 1896.050 1686.500 ;
        RECT 1892.050 1631.900 1892.370 1631.960 ;
        RECT 1896.650 1631.900 1896.970 1631.960 ;
        RECT 1892.050 1631.760 1896.970 1631.900 ;
        RECT 1892.050 1631.700 1892.370 1631.760 ;
        RECT 1896.650 1631.700 1896.970 1631.760 ;
        RECT 1896.650 38.660 1896.970 38.720 ;
        RECT 2761.910 38.660 2762.230 38.720 ;
        RECT 1896.650 38.520 2762.230 38.660 ;
        RECT 1896.650 38.460 1896.970 38.520 ;
        RECT 2761.910 38.460 2762.230 38.520 ;
      LAYER via ;
        RECT 1892.080 1686.440 1892.340 1686.700 ;
        RECT 1895.760 1686.440 1896.020 1686.700 ;
        RECT 1892.080 1631.700 1892.340 1631.960 ;
        RECT 1896.680 1631.700 1896.940 1631.960 ;
        RECT 1896.680 38.460 1896.940 38.720 ;
        RECT 2761.940 38.460 2762.200 38.720 ;
      LAYER met2 ;
        RECT 1895.750 1700.000 1896.030 1704.000 ;
        RECT 1895.820 1686.730 1895.960 1700.000 ;
        RECT 1892.080 1686.410 1892.340 1686.730 ;
        RECT 1895.760 1686.410 1896.020 1686.730 ;
        RECT 1892.140 1631.990 1892.280 1686.410 ;
        RECT 1892.080 1631.670 1892.340 1631.990 ;
        RECT 1896.680 1631.670 1896.940 1631.990 ;
        RECT 1896.740 38.750 1896.880 1631.670 ;
        RECT 1896.680 38.430 1896.940 38.750 ;
        RECT 2761.940 38.430 2762.200 38.750 ;
        RECT 2762.000 2.400 2762.140 38.430 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 0.300 ;
=======
      LAYER met1 ;
        RECT 835.430 32.200 835.750 32.260 ;
        RECT 1375.010 32.200 1375.330 32.260 ;
        RECT 835.430 32.060 1375.330 32.200 ;
        RECT 835.430 32.000 835.750 32.060 ;
        RECT 1375.010 32.000 1375.330 32.060 ;
      LAYER via ;
        RECT 835.460 32.000 835.720 32.260 ;
        RECT 1375.040 32.000 1375.300 32.260 ;
      LAYER met2 ;
        RECT 1375.030 1700.000 1375.310 1704.000 ;
        RECT 1375.100 32.290 1375.240 1700.000 ;
        RECT 835.460 31.970 835.720 32.290 ;
        RECT 1375.040 31.970 1375.300 32.290 ;
        RECT 835.520 2.400 835.660 31.970 ;
        RECT 835.310 -4.800 835.870 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1900.330 1695.480 1900.650 1695.540 ;
        RECT 1902.630 1695.480 1902.950 1695.540 ;
        RECT 1900.330 1695.340 1902.950 1695.480 ;
        RECT 1900.330 1695.280 1900.650 1695.340 ;
        RECT 1902.630 1695.280 1902.950 1695.340 ;
        RECT 1902.630 38.320 1902.950 38.380 ;
        RECT 2779.850 38.320 2780.170 38.380 ;
        RECT 1902.630 38.180 2780.170 38.320 ;
        RECT 1902.630 38.120 1902.950 38.180 ;
        RECT 2779.850 38.120 2780.170 38.180 ;
      LAYER via ;
        RECT 1900.360 1695.280 1900.620 1695.540 ;
        RECT 1902.660 1695.280 1902.920 1695.540 ;
        RECT 1902.660 38.120 1902.920 38.380 ;
        RECT 2779.880 38.120 2780.140 38.380 ;
      LAYER met2 ;
        RECT 1900.350 1700.000 1900.630 1704.000 ;
        RECT 1900.420 1695.570 1900.560 1700.000 ;
        RECT 1900.360 1695.250 1900.620 1695.570 ;
        RECT 1902.660 1695.250 1902.920 1695.570 ;
        RECT 1902.720 38.410 1902.860 1695.250 ;
        RECT 1902.660 38.090 1902.920 38.410 ;
        RECT 2779.880 38.090 2780.140 38.410 ;
        RECT 2779.940 2.400 2780.080 38.090 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 0.300 ;
=======
      LAYER met1 ;
        RECT 1904.470 1631.900 1904.790 1631.960 ;
        RECT 1910.450 1631.900 1910.770 1631.960 ;
        RECT 1904.470 1631.760 1910.770 1631.900 ;
        RECT 1904.470 1631.700 1904.790 1631.760 ;
        RECT 1910.450 1631.700 1910.770 1631.760 ;
        RECT 1910.450 37.980 1910.770 38.040 ;
        RECT 2797.790 37.980 2798.110 38.040 ;
        RECT 1910.450 37.840 2798.110 37.980 ;
        RECT 1910.450 37.780 1910.770 37.840 ;
        RECT 2797.790 37.780 2798.110 37.840 ;
      LAYER via ;
        RECT 1904.500 1631.700 1904.760 1631.960 ;
        RECT 1910.480 1631.700 1910.740 1631.960 ;
        RECT 1910.480 37.780 1910.740 38.040 ;
        RECT 2797.820 37.780 2798.080 38.040 ;
      LAYER met2 ;
        RECT 1905.410 1700.410 1905.690 1704.000 ;
        RECT 1904.560 1700.270 1905.690 1700.410 ;
        RECT 1904.560 1631.990 1904.700 1700.270 ;
        RECT 1905.410 1700.000 1905.690 1700.270 ;
        RECT 1904.500 1631.670 1904.760 1631.990 ;
        RECT 1910.480 1631.670 1910.740 1631.990 ;
        RECT 1910.540 38.070 1910.680 1631.670 ;
        RECT 1910.480 37.750 1910.740 38.070 ;
        RECT 2797.820 37.750 2798.080 38.070 ;
        RECT 2797.880 2.400 2798.020 37.750 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2815.610 -4.800 2816.170 0.300 ;
=======
        RECT 1910.010 1700.000 1910.290 1704.000 ;
        RECT 1910.080 41.325 1910.220 1700.000 ;
        RECT 1910.010 40.955 1910.290 41.325 ;
        RECT 2815.750 40.955 2816.030 41.325 ;
        RECT 2815.820 2.400 2815.960 40.955 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
      LAYER via2 ;
        RECT 1910.010 41.000 1910.290 41.280 ;
        RECT 2815.750 41.000 2816.030 41.280 ;
      LAYER met3 ;
        RECT 1909.985 41.290 1910.315 41.305 ;
        RECT 2815.725 41.290 2816.055 41.305 ;
        RECT 1909.985 40.990 2816.055 41.290 ;
        RECT 1909.985 40.975 1910.315 40.990 ;
        RECT 2815.725 40.975 2816.055 40.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1911.370 1684.260 1911.690 1684.320 ;
        RECT 1915.050 1684.260 1915.370 1684.320 ;
        RECT 1911.370 1684.120 1915.370 1684.260 ;
        RECT 1911.370 1684.060 1911.690 1684.120 ;
        RECT 1915.050 1684.060 1915.370 1684.120 ;
        RECT 1911.370 1631.900 1911.690 1631.960 ;
        RECT 1917.350 1631.900 1917.670 1631.960 ;
        RECT 1911.370 1631.760 1917.670 1631.900 ;
        RECT 1911.370 1631.700 1911.690 1631.760 ;
        RECT 1917.350 1631.700 1917.670 1631.760 ;
      LAYER via ;
        RECT 1911.400 1684.060 1911.660 1684.320 ;
        RECT 1915.080 1684.060 1915.340 1684.320 ;
        RECT 1911.400 1631.700 1911.660 1631.960 ;
        RECT 1917.380 1631.700 1917.640 1631.960 ;
      LAYER met2 ;
        RECT 1915.070 1700.000 1915.350 1704.000 ;
        RECT 1915.140 1684.350 1915.280 1700.000 ;
        RECT 1911.400 1684.030 1911.660 1684.350 ;
        RECT 1915.080 1684.030 1915.340 1684.350 ;
        RECT 1911.460 1631.990 1911.600 1684.030 ;
        RECT 1911.400 1631.670 1911.660 1631.990 ;
        RECT 1917.380 1631.670 1917.640 1631.990 ;
        RECT 1917.440 40.645 1917.580 1631.670 ;
        RECT 1917.370 40.275 1917.650 40.645 ;
        RECT 2833.690 40.275 2833.970 40.645 ;
        RECT 2833.760 2.400 2833.900 40.275 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
      LAYER via2 ;
        RECT 1917.370 40.320 1917.650 40.600 ;
        RECT 2833.690 40.320 2833.970 40.600 ;
      LAYER met3 ;
        RECT 1917.345 40.610 1917.675 40.625 ;
        RECT 2833.665 40.610 2833.995 40.625 ;
        RECT 1917.345 40.310 2833.995 40.610 ;
        RECT 1917.345 40.295 1917.675 40.310 ;
        RECT 2833.665 40.295 2833.995 40.310 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1919.650 1677.460 1919.970 1677.520 ;
        RECT 1923.330 1677.460 1923.650 1677.520 ;
        RECT 1919.650 1677.320 1923.650 1677.460 ;
        RECT 1919.650 1677.260 1919.970 1677.320 ;
        RECT 1923.330 1677.260 1923.650 1677.320 ;
      LAYER via ;
        RECT 1919.680 1677.260 1919.940 1677.520 ;
        RECT 1923.360 1677.260 1923.620 1677.520 ;
      LAYER met2 ;
        RECT 1919.670 1700.000 1919.950 1704.000 ;
        RECT 1919.740 1677.550 1919.880 1700.000 ;
        RECT 1919.680 1677.230 1919.940 1677.550 ;
        RECT 1923.360 1677.230 1923.620 1677.550 ;
        RECT 1923.420 39.965 1923.560 1677.230 ;
        RECT 1923.350 39.595 1923.630 39.965 ;
        RECT 2851.170 39.595 2851.450 39.965 ;
        RECT 2851.240 2.400 2851.380 39.595 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
      LAYER via2 ;
        RECT 1923.350 39.640 1923.630 39.920 ;
        RECT 2851.170 39.640 2851.450 39.920 ;
      LAYER met3 ;
        RECT 1923.325 39.930 1923.655 39.945 ;
        RECT 2851.145 39.930 2851.475 39.945 ;
        RECT 1923.325 39.630 2851.475 39.930 ;
        RECT 1923.325 39.615 1923.655 39.630 ;
        RECT 2851.145 39.615 2851.475 39.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2868.970 -4.800 2869.530 0.300 ;
=======
        RECT 1924.730 1700.410 1925.010 1704.000 ;
        RECT 1923.420 1700.270 1925.010 1700.410 ;
        RECT 1923.420 1677.970 1923.560 1700.270 ;
        RECT 1924.730 1700.000 1925.010 1700.270 ;
        RECT 1922.960 1677.830 1923.560 1677.970 ;
        RECT 1922.960 39.285 1923.100 1677.830 ;
        RECT 1922.890 38.915 1923.170 39.285 ;
        RECT 2869.110 38.915 2869.390 39.285 ;
        RECT 2869.180 2.400 2869.320 38.915 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
      LAYER via2 ;
        RECT 1922.890 38.960 1923.170 39.240 ;
        RECT 2869.110 38.960 2869.390 39.240 ;
      LAYER met3 ;
        RECT 1922.865 39.250 1923.195 39.265 ;
        RECT 2869.085 39.250 2869.415 39.265 ;
        RECT 1922.865 38.950 2869.415 39.250 ;
        RECT 1922.865 38.935 1923.195 38.950 ;
        RECT 2869.085 38.935 2869.415 38.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2886.910 -4.800 2887.470 0.300 ;
=======
        RECT 1929.330 1700.410 1929.610 1704.000 ;
        RECT 1929.330 1700.270 1930.920 1700.410 ;
        RECT 1929.330 1700.000 1929.610 1700.270 ;
        RECT 1930.780 38.605 1930.920 1700.270 ;
        RECT 1930.710 38.235 1930.990 38.605 ;
        RECT 2887.050 38.235 2887.330 38.605 ;
        RECT 2887.120 2.400 2887.260 38.235 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
      LAYER via2 ;
        RECT 1930.710 38.280 1930.990 38.560 ;
        RECT 2887.050 38.280 2887.330 38.560 ;
      LAYER met3 ;
        RECT 1930.685 38.570 1931.015 38.585 ;
        RECT 2887.025 38.570 2887.355 38.585 ;
        RECT 1930.685 38.270 2887.355 38.570 ;
        RECT 1930.685 38.255 1931.015 38.270 ;
        RECT 2887.025 38.255 2887.355 38.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1934.370 1684.260 1934.690 1684.320 ;
        RECT 1938.050 1684.260 1938.370 1684.320 ;
        RECT 1934.370 1684.120 1938.370 1684.260 ;
        RECT 1934.370 1684.060 1934.690 1684.120 ;
        RECT 1938.050 1684.060 1938.370 1684.120 ;
      LAYER via ;
        RECT 1934.400 1684.060 1934.660 1684.320 ;
        RECT 1938.080 1684.060 1938.340 1684.320 ;
      LAYER met2 ;
        RECT 1934.390 1700.000 1934.670 1704.000 ;
        RECT 1934.460 1684.350 1934.600 1700.000 ;
        RECT 1934.400 1684.030 1934.660 1684.350 ;
        RECT 1938.080 1684.030 1938.340 1684.350 ;
        RECT 1938.140 37.925 1938.280 1684.030 ;
        RECT 1938.070 37.555 1938.350 37.925 ;
        RECT 2904.990 37.555 2905.270 37.925 ;
        RECT 2905.060 2.400 2905.200 37.555 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 1938.070 37.600 1938.350 37.880 ;
        RECT 2904.990 37.600 2905.270 37.880 ;
      LAYER met3 ;
        RECT 1938.045 37.890 1938.375 37.905 ;
        RECT 2904.965 37.890 2905.295 37.905 ;
        RECT 1938.045 37.590 2905.295 37.890 ;
        RECT 1938.045 37.575 1938.375 37.590 ;
        RECT 2904.965 37.575 2905.295 37.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 0.300 ;
=======
      LAYER met1 ;
        RECT 852.910 32.540 853.230 32.600 ;
        RECT 1380.530 32.540 1380.850 32.600 ;
        RECT 852.910 32.400 1380.850 32.540 ;
        RECT 852.910 32.340 853.230 32.400 ;
        RECT 1380.530 32.340 1380.850 32.400 ;
      LAYER via ;
        RECT 852.940 32.340 853.200 32.600 ;
        RECT 1380.560 32.340 1380.820 32.600 ;
      LAYER met2 ;
        RECT 1380.090 1700.410 1380.370 1704.000 ;
        RECT 1380.090 1700.270 1380.760 1700.410 ;
        RECT 1380.090 1700.000 1380.370 1700.270 ;
        RECT 1380.620 32.630 1380.760 1700.270 ;
        RECT 852.940 32.310 853.200 32.630 ;
        RECT 1380.560 32.310 1380.820 32.630 ;
        RECT 853.000 2.400 853.140 32.310 ;
        RECT 852.790 -4.800 853.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1380.990 1678.140 1381.310 1678.200 ;
        RECT 1383.750 1678.140 1384.070 1678.200 ;
        RECT 1380.990 1678.000 1384.070 1678.140 ;
        RECT 1380.990 1677.940 1381.310 1678.000 ;
        RECT 1383.750 1677.940 1384.070 1678.000 ;
        RECT 870.850 32.880 871.170 32.940 ;
        RECT 1380.990 32.880 1381.310 32.940 ;
        RECT 870.850 32.740 1381.310 32.880 ;
        RECT 870.850 32.680 871.170 32.740 ;
        RECT 1380.990 32.680 1381.310 32.740 ;
      LAYER via ;
        RECT 1381.020 1677.940 1381.280 1678.200 ;
        RECT 1383.780 1677.940 1384.040 1678.200 ;
        RECT 870.880 32.680 871.140 32.940 ;
        RECT 1381.020 32.680 1381.280 32.940 ;
      LAYER met2 ;
        RECT 1384.690 1700.410 1384.970 1704.000 ;
        RECT 1383.840 1700.270 1384.970 1700.410 ;
        RECT 1383.840 1678.230 1383.980 1700.270 ;
        RECT 1384.690 1700.000 1384.970 1700.270 ;
        RECT 1381.020 1677.910 1381.280 1678.230 ;
        RECT 1383.780 1677.910 1384.040 1678.230 ;
        RECT 1381.080 32.970 1381.220 1677.910 ;
        RECT 870.880 32.650 871.140 32.970 ;
        RECT 1381.020 32.650 1381.280 32.970 ;
        RECT 870.940 2.400 871.080 32.650 ;
        RECT 870.730 -4.800 871.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 0.300 ;
=======
      LAYER met1 ;
        RECT 888.790 33.220 889.110 33.280 ;
        RECT 1388.810 33.220 1389.130 33.280 ;
        RECT 888.790 33.080 1389.130 33.220 ;
        RECT 888.790 33.020 889.110 33.080 ;
        RECT 1388.810 33.020 1389.130 33.080 ;
      LAYER via ;
        RECT 888.820 33.020 889.080 33.280 ;
        RECT 1388.840 33.020 1389.100 33.280 ;
      LAYER met2 ;
        RECT 1389.750 1700.410 1390.030 1704.000 ;
        RECT 1388.900 1700.270 1390.030 1700.410 ;
        RECT 1388.900 33.310 1389.040 1700.270 ;
        RECT 1389.750 1700.000 1390.030 1700.270 ;
        RECT 888.820 32.990 889.080 33.310 ;
        RECT 1388.840 32.990 1389.100 33.310 ;
        RECT 888.880 2.400 889.020 32.990 ;
        RECT 888.670 -4.800 889.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 0.300 ;
=======
      LAYER met1 ;
        RECT 906.730 33.560 907.050 33.620 ;
        RECT 1394.330 33.560 1394.650 33.620 ;
        RECT 906.730 33.420 1394.650 33.560 ;
        RECT 906.730 33.360 907.050 33.420 ;
        RECT 1394.330 33.360 1394.650 33.420 ;
      LAYER via ;
        RECT 906.760 33.360 907.020 33.620 ;
        RECT 1394.360 33.360 1394.620 33.620 ;
      LAYER met2 ;
        RECT 1394.350 1700.000 1394.630 1704.000 ;
        RECT 1394.420 33.650 1394.560 1700.000 ;
        RECT 906.760 33.330 907.020 33.650 ;
        RECT 1394.360 33.330 1394.620 33.650 ;
        RECT 906.820 2.400 906.960 33.330 ;
        RECT 906.610 -4.800 907.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1394.790 1678.140 1395.110 1678.200 ;
        RECT 1398.010 1678.140 1398.330 1678.200 ;
        RECT 1394.790 1678.000 1398.330 1678.140 ;
        RECT 1394.790 1677.940 1395.110 1678.000 ;
        RECT 1398.010 1677.940 1398.330 1678.000 ;
        RECT 924.210 33.900 924.530 33.960 ;
        RECT 1394.790 33.900 1395.110 33.960 ;
        RECT 924.210 33.760 1395.110 33.900 ;
        RECT 924.210 33.700 924.530 33.760 ;
        RECT 1394.790 33.700 1395.110 33.760 ;
      LAYER via ;
        RECT 1394.820 1677.940 1395.080 1678.200 ;
        RECT 1398.040 1677.940 1398.300 1678.200 ;
        RECT 924.240 33.700 924.500 33.960 ;
        RECT 1394.820 33.700 1395.080 33.960 ;
      LAYER met2 ;
        RECT 1399.410 1700.410 1399.690 1704.000 ;
        RECT 1398.100 1700.270 1399.690 1700.410 ;
        RECT 1398.100 1678.230 1398.240 1700.270 ;
        RECT 1399.410 1700.000 1399.690 1700.270 ;
        RECT 1394.820 1677.910 1395.080 1678.230 ;
        RECT 1398.040 1677.910 1398.300 1678.230 ;
        RECT 1394.880 33.990 1395.020 1677.910 ;
        RECT 924.240 33.670 924.500 33.990 ;
        RECT 1394.820 33.670 1395.080 33.990 ;
        RECT 924.300 2.400 924.440 33.670 ;
        RECT 924.090 -4.800 924.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1401.230 1675.080 1401.550 1675.140 ;
        RECT 1403.070 1675.080 1403.390 1675.140 ;
        RECT 1401.230 1674.940 1403.390 1675.080 ;
        RECT 1401.230 1674.880 1401.550 1674.940 ;
        RECT 1403.070 1674.880 1403.390 1674.940 ;
        RECT 942.150 34.240 942.470 34.300 ;
        RECT 1401.230 34.240 1401.550 34.300 ;
        RECT 942.150 34.100 1401.550 34.240 ;
        RECT 942.150 34.040 942.470 34.100 ;
        RECT 1401.230 34.040 1401.550 34.100 ;
      LAYER via ;
        RECT 1401.260 1674.880 1401.520 1675.140 ;
        RECT 1403.100 1674.880 1403.360 1675.140 ;
        RECT 942.180 34.040 942.440 34.300 ;
        RECT 1401.260 34.040 1401.520 34.300 ;
      LAYER met2 ;
        RECT 1404.010 1700.410 1404.290 1704.000 ;
        RECT 1403.160 1700.270 1404.290 1700.410 ;
        RECT 1403.160 1675.170 1403.300 1700.270 ;
        RECT 1404.010 1700.000 1404.290 1700.270 ;
        RECT 1401.260 1674.850 1401.520 1675.170 ;
        RECT 1403.100 1674.850 1403.360 1675.170 ;
        RECT 1401.320 34.330 1401.460 1674.850 ;
        RECT 942.180 34.010 942.440 34.330 ;
        RECT 1401.260 34.010 1401.520 34.330 ;
        RECT 942.240 2.400 942.380 34.010 ;
        RECT 942.030 -4.800 942.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 0.300 ;
=======
      LAYER met1 ;
        RECT 960.090 30.500 960.410 30.560 ;
        RECT 1408.130 30.500 1408.450 30.560 ;
        RECT 960.090 30.360 1408.450 30.500 ;
        RECT 960.090 30.300 960.410 30.360 ;
        RECT 1408.130 30.300 1408.450 30.360 ;
      LAYER via ;
        RECT 960.120 30.300 960.380 30.560 ;
        RECT 1408.160 30.300 1408.420 30.560 ;
      LAYER met2 ;
        RECT 1409.070 1700.410 1409.350 1704.000 ;
        RECT 1408.220 1700.270 1409.350 1700.410 ;
        RECT 1408.220 30.590 1408.360 1700.270 ;
        RECT 1409.070 1700.000 1409.350 1700.270 ;
        RECT 960.120 30.270 960.380 30.590 ;
        RECT 1408.160 30.270 1408.420 30.590 ;
        RECT 960.180 2.400 960.320 30.270 ;
        RECT 959.970 -4.800 960.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 0.300 ;
=======
      LAYER met1 ;
        RECT 1408.590 1678.140 1408.910 1678.200 ;
        RECT 1412.730 1678.140 1413.050 1678.200 ;
        RECT 1408.590 1678.000 1413.050 1678.140 ;
        RECT 1408.590 1677.940 1408.910 1678.000 ;
        RECT 1412.730 1677.940 1413.050 1678.000 ;
        RECT 978.030 30.160 978.350 30.220 ;
        RECT 1408.590 30.160 1408.910 30.220 ;
        RECT 978.030 30.020 1408.910 30.160 ;
        RECT 978.030 29.960 978.350 30.020 ;
        RECT 1408.590 29.960 1408.910 30.020 ;
      LAYER via ;
        RECT 1408.620 1677.940 1408.880 1678.200 ;
        RECT 1412.760 1677.940 1413.020 1678.200 ;
        RECT 978.060 29.960 978.320 30.220 ;
        RECT 1408.620 29.960 1408.880 30.220 ;
      LAYER met2 ;
        RECT 1413.670 1700.410 1413.950 1704.000 ;
        RECT 1412.820 1700.270 1413.950 1700.410 ;
        RECT 1412.820 1678.230 1412.960 1700.270 ;
        RECT 1413.670 1700.000 1413.950 1700.270 ;
        RECT 1408.620 1677.910 1408.880 1678.230 ;
        RECT 1412.760 1677.910 1413.020 1678.230 ;
        RECT 1408.680 30.250 1408.820 1677.910 ;
        RECT 978.060 29.930 978.320 30.250 ;
        RECT 1408.620 29.930 1408.880 30.250 ;
        RECT 978.120 2.400 978.260 29.930 ;
        RECT 977.910 -4.800 978.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 656.830 -4.800 657.390 0.300 ;
=======
        RECT 1327.190 1700.410 1327.470 1704.000 ;
        RECT 1325.880 1700.270 1327.470 1700.410 ;
        RECT 1325.880 33.845 1326.020 1700.270 ;
        RECT 1327.190 1700.000 1327.470 1700.270 ;
        RECT 656.970 33.475 657.250 33.845 ;
        RECT 1325.810 33.475 1326.090 33.845 ;
        RECT 657.040 2.400 657.180 33.475 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 656.970 33.520 657.250 33.800 ;
        RECT 1325.810 33.520 1326.090 33.800 ;
      LAYER met3 ;
        RECT 656.945 33.810 657.275 33.825 ;
        RECT 1325.785 33.810 1326.115 33.825 ;
        RECT 656.945 33.510 1326.115 33.810 ;
        RECT 656.945 33.495 657.275 33.510 ;
        RECT 1325.785 33.495 1326.115 33.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1415.030 1678.480 1415.350 1678.540 ;
        RECT 1417.330 1678.480 1417.650 1678.540 ;
        RECT 1415.030 1678.340 1417.650 1678.480 ;
        RECT 1415.030 1678.280 1415.350 1678.340 ;
        RECT 1417.330 1678.280 1417.650 1678.340 ;
        RECT 995.970 29.820 996.290 29.880 ;
        RECT 1415.030 29.820 1415.350 29.880 ;
        RECT 995.970 29.680 1415.350 29.820 ;
        RECT 995.970 29.620 996.290 29.680 ;
        RECT 1415.030 29.620 1415.350 29.680 ;
      LAYER via ;
        RECT 1415.060 1678.280 1415.320 1678.540 ;
        RECT 1417.360 1678.280 1417.620 1678.540 ;
        RECT 996.000 29.620 996.260 29.880 ;
        RECT 1415.060 29.620 1415.320 29.880 ;
      LAYER met2 ;
        RECT 1418.730 1700.410 1419.010 1704.000 ;
        RECT 1417.420 1700.270 1419.010 1700.410 ;
        RECT 1417.420 1678.570 1417.560 1700.270 ;
        RECT 1418.730 1700.000 1419.010 1700.270 ;
        RECT 1415.060 1678.250 1415.320 1678.570 ;
        RECT 1417.360 1678.250 1417.620 1678.570 ;
        RECT 1415.120 29.910 1415.260 1678.250 ;
        RECT 996.000 29.590 996.260 29.910 ;
        RECT 1415.060 29.590 1415.320 29.910 ;
        RECT 996.060 2.400 996.200 29.590 ;
        RECT 995.850 -4.800 996.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 0.300 ;
=======
      LAYER met1 ;
        RECT 1013.450 29.480 1013.770 29.540 ;
        RECT 1422.390 29.480 1422.710 29.540 ;
        RECT 1013.450 29.340 1422.710 29.480 ;
        RECT 1013.450 29.280 1013.770 29.340 ;
        RECT 1422.390 29.280 1422.710 29.340 ;
      LAYER via ;
        RECT 1013.480 29.280 1013.740 29.540 ;
        RECT 1422.420 29.280 1422.680 29.540 ;
      LAYER met2 ;
        RECT 1423.330 1700.410 1423.610 1704.000 ;
        RECT 1422.480 1700.270 1423.610 1700.410 ;
        RECT 1422.480 29.570 1422.620 1700.270 ;
        RECT 1423.330 1700.000 1423.610 1700.270 ;
        RECT 1013.480 29.250 1013.740 29.570 ;
        RECT 1422.420 29.250 1422.680 29.570 ;
        RECT 1013.540 2.400 1013.680 29.250 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 0.300 ;
=======
      LAYER met1 ;
        RECT 1031.390 29.140 1031.710 29.200 ;
        RECT 1429.290 29.140 1429.610 29.200 ;
        RECT 1031.390 29.000 1429.610 29.140 ;
        RECT 1031.390 28.940 1031.710 29.000 ;
        RECT 1429.290 28.940 1429.610 29.000 ;
      LAYER via ;
        RECT 1031.420 28.940 1031.680 29.200 ;
        RECT 1429.320 28.940 1429.580 29.200 ;
      LAYER met2 ;
        RECT 1428.390 1700.410 1428.670 1704.000 ;
        RECT 1428.390 1700.270 1429.520 1700.410 ;
        RECT 1428.390 1700.000 1428.670 1700.270 ;
        RECT 1429.380 29.230 1429.520 1700.270 ;
        RECT 1031.420 28.910 1031.680 29.230 ;
        RECT 1429.320 28.910 1429.580 29.230 ;
        RECT 1031.480 2.400 1031.620 28.910 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1428.830 1678.480 1429.150 1678.540 ;
        RECT 1432.050 1678.480 1432.370 1678.540 ;
        RECT 1428.830 1678.340 1432.370 1678.480 ;
        RECT 1428.830 1678.280 1429.150 1678.340 ;
        RECT 1432.050 1678.280 1432.370 1678.340 ;
        RECT 1049.330 28.800 1049.650 28.860 ;
        RECT 1428.830 28.800 1429.150 28.860 ;
        RECT 1049.330 28.660 1429.150 28.800 ;
        RECT 1049.330 28.600 1049.650 28.660 ;
        RECT 1428.830 28.600 1429.150 28.660 ;
      LAYER via ;
        RECT 1428.860 1678.280 1429.120 1678.540 ;
        RECT 1432.080 1678.280 1432.340 1678.540 ;
        RECT 1049.360 28.600 1049.620 28.860 ;
        RECT 1428.860 28.600 1429.120 28.860 ;
      LAYER met2 ;
        RECT 1432.990 1700.410 1433.270 1704.000 ;
        RECT 1432.140 1700.270 1433.270 1700.410 ;
        RECT 1432.140 1678.570 1432.280 1700.270 ;
        RECT 1432.990 1700.000 1433.270 1700.270 ;
        RECT 1428.860 1678.250 1429.120 1678.570 ;
        RECT 1432.080 1678.250 1432.340 1678.570 ;
        RECT 1428.920 28.890 1429.060 1678.250 ;
        RECT 1049.360 28.570 1049.620 28.890 ;
        RECT 1428.860 28.570 1429.120 28.890 ;
        RECT 1049.420 2.400 1049.560 28.570 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 0.300 ;
=======
      LAYER met1 ;
        RECT 1067.270 28.460 1067.590 28.520 ;
        RECT 1437.110 28.460 1437.430 28.520 ;
        RECT 1067.270 28.320 1437.430 28.460 ;
        RECT 1067.270 28.260 1067.590 28.320 ;
        RECT 1437.110 28.260 1437.430 28.320 ;
      LAYER via ;
        RECT 1067.300 28.260 1067.560 28.520 ;
        RECT 1437.140 28.260 1437.400 28.520 ;
      LAYER met2 ;
        RECT 1438.050 1700.410 1438.330 1704.000 ;
        RECT 1437.200 1700.270 1438.330 1700.410 ;
        RECT 1437.200 28.550 1437.340 1700.270 ;
        RECT 1438.050 1700.000 1438.330 1700.270 ;
        RECT 1067.300 28.230 1067.560 28.550 ;
        RECT 1437.140 28.230 1437.400 28.550 ;
        RECT 1067.360 2.400 1067.500 28.230 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1085.210 28.120 1085.530 28.180 ;
        RECT 1443.090 28.120 1443.410 28.180 ;
        RECT 1085.210 27.980 1443.410 28.120 ;
        RECT 1085.210 27.920 1085.530 27.980 ;
        RECT 1443.090 27.920 1443.410 27.980 ;
      LAYER via ;
        RECT 1085.240 27.920 1085.500 28.180 ;
        RECT 1443.120 27.920 1443.380 28.180 ;
      LAYER met2 ;
        RECT 1442.650 1700.410 1442.930 1704.000 ;
        RECT 1442.650 1700.270 1443.320 1700.410 ;
        RECT 1442.650 1700.000 1442.930 1700.270 ;
        RECT 1443.180 28.210 1443.320 1700.270 ;
        RECT 1085.240 27.890 1085.500 28.210 ;
        RECT 1443.120 27.890 1443.380 28.210 ;
        RECT 1085.300 2.400 1085.440 27.890 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 0.300 ;
=======
      LAYER li1 ;
        RECT 1445.005 1545.045 1445.175 1587.035 ;
        RECT 1446.845 1048.645 1447.015 1089.955 ;
        RECT 1445.005 783.105 1445.175 807.075 ;
        RECT 1444.545 620.925 1444.715 628.235 ;
        RECT 1444.545 434.265 1444.715 475.915 ;
        RECT 1444.545 227.885 1444.715 275.995 ;
        RECT 1445.005 131.325 1445.175 159.035 ;
        RECT 1444.085 27.625 1444.255 36.295 ;
      LAYER mcon ;
        RECT 1445.005 1586.865 1445.175 1587.035 ;
        RECT 1446.845 1089.785 1447.015 1089.955 ;
        RECT 1445.005 806.905 1445.175 807.075 ;
        RECT 1444.545 628.065 1444.715 628.235 ;
        RECT 1444.545 475.745 1444.715 475.915 ;
        RECT 1444.545 275.825 1444.715 275.995 ;
        RECT 1445.005 158.865 1445.175 159.035 ;
        RECT 1444.085 36.125 1444.255 36.295 ;
      LAYER met1 ;
        RECT 1444.930 1587.020 1445.250 1587.080 ;
        RECT 1444.735 1586.880 1445.250 1587.020 ;
        RECT 1444.930 1586.820 1445.250 1586.880 ;
        RECT 1444.945 1545.200 1445.235 1545.245 ;
        RECT 1445.390 1545.200 1445.710 1545.260 ;
        RECT 1444.945 1545.060 1445.710 1545.200 ;
        RECT 1444.945 1545.015 1445.235 1545.060 ;
        RECT 1445.390 1545.000 1445.710 1545.060 ;
        RECT 1444.930 1497.600 1445.250 1497.660 ;
        RECT 1445.390 1497.600 1445.710 1497.660 ;
        RECT 1444.930 1497.460 1445.710 1497.600 ;
        RECT 1444.930 1497.400 1445.250 1497.460 ;
        RECT 1445.390 1497.400 1445.710 1497.460 ;
        RECT 1444.930 1463.260 1445.250 1463.320 ;
        RECT 1444.560 1463.120 1445.250 1463.260 ;
        RECT 1444.560 1462.640 1444.700 1463.120 ;
        RECT 1444.930 1463.060 1445.250 1463.120 ;
        RECT 1444.470 1462.380 1444.790 1462.640 ;
        RECT 1444.470 1400.700 1444.790 1400.760 ;
        RECT 1444.930 1400.700 1445.250 1400.760 ;
        RECT 1444.470 1400.560 1445.250 1400.700 ;
        RECT 1444.470 1400.500 1444.790 1400.560 ;
        RECT 1444.930 1400.500 1445.250 1400.560 ;
        RECT 1444.470 1352.560 1444.790 1352.820 ;
        RECT 1444.560 1352.080 1444.700 1352.560 ;
        RECT 1444.930 1352.080 1445.250 1352.140 ;
        RECT 1444.560 1351.940 1445.250 1352.080 ;
        RECT 1444.930 1351.880 1445.250 1351.940 ;
        RECT 1444.470 1249.060 1444.790 1249.120 ;
        RECT 1444.930 1249.060 1445.250 1249.120 ;
        RECT 1444.470 1248.920 1445.250 1249.060 ;
        RECT 1444.470 1248.860 1444.790 1248.920 ;
        RECT 1444.930 1248.860 1445.250 1248.920 ;
        RECT 1444.930 1159.640 1445.250 1159.700 ;
        RECT 1444.560 1159.500 1445.250 1159.640 ;
        RECT 1444.560 1159.360 1444.700 1159.500 ;
        RECT 1444.930 1159.440 1445.250 1159.500 ;
        RECT 1444.470 1159.100 1444.790 1159.360 ;
        RECT 1444.010 1145.360 1444.330 1145.420 ;
        RECT 1444.470 1145.360 1444.790 1145.420 ;
        RECT 1444.010 1145.220 1444.790 1145.360 ;
        RECT 1444.010 1145.160 1444.330 1145.220 ;
        RECT 1444.470 1145.160 1444.790 1145.220 ;
        RECT 1444.930 1097.080 1445.250 1097.140 ;
        RECT 1446.770 1097.080 1447.090 1097.140 ;
        RECT 1444.930 1096.940 1447.090 1097.080 ;
        RECT 1444.930 1096.880 1445.250 1096.940 ;
        RECT 1446.770 1096.880 1447.090 1096.940 ;
        RECT 1446.770 1089.940 1447.090 1090.000 ;
        RECT 1446.575 1089.800 1447.090 1089.940 ;
        RECT 1446.770 1089.740 1447.090 1089.800 ;
        RECT 1446.770 1048.800 1447.090 1048.860 ;
        RECT 1446.575 1048.660 1447.090 1048.800 ;
        RECT 1446.770 1048.600 1447.090 1048.660 ;
        RECT 1444.470 862.820 1444.790 862.880 ;
        RECT 1445.390 862.820 1445.710 862.880 ;
        RECT 1444.470 862.680 1445.710 862.820 ;
        RECT 1444.470 862.620 1444.790 862.680 ;
        RECT 1445.390 862.620 1445.710 862.680 ;
        RECT 1444.930 807.060 1445.250 807.120 ;
        RECT 1444.735 806.920 1445.250 807.060 ;
        RECT 1444.930 806.860 1445.250 806.920 ;
        RECT 1444.930 783.260 1445.250 783.320 ;
        RECT 1444.735 783.120 1445.250 783.260 ;
        RECT 1444.930 783.060 1445.250 783.120 ;
        RECT 1444.930 724.440 1445.250 724.500 ;
        RECT 1445.390 724.440 1445.710 724.500 ;
        RECT 1444.930 724.300 1445.710 724.440 ;
        RECT 1444.930 724.240 1445.250 724.300 ;
        RECT 1445.390 724.240 1445.710 724.300 ;
        RECT 1444.470 676.160 1444.790 676.220 ;
        RECT 1445.390 676.160 1445.710 676.220 ;
        RECT 1444.470 676.020 1445.710 676.160 ;
        RECT 1444.470 675.960 1444.790 676.020 ;
        RECT 1445.390 675.960 1445.710 676.020 ;
        RECT 1444.485 628.220 1444.775 628.265 ;
        RECT 1445.390 628.220 1445.710 628.280 ;
        RECT 1444.485 628.080 1445.710 628.220 ;
        RECT 1444.485 628.035 1444.775 628.080 ;
        RECT 1445.390 628.020 1445.710 628.080 ;
        RECT 1444.470 621.080 1444.790 621.140 ;
        RECT 1444.275 620.940 1444.790 621.080 ;
        RECT 1444.470 620.880 1444.790 620.940 ;
        RECT 1444.470 572.800 1444.790 572.860 ;
        RECT 1445.390 572.800 1445.710 572.860 ;
        RECT 1444.470 572.660 1445.710 572.800 ;
        RECT 1444.470 572.600 1444.790 572.660 ;
        RECT 1445.390 572.600 1445.710 572.660 ;
        RECT 1444.470 475.900 1444.790 475.960 ;
        RECT 1444.275 475.760 1444.790 475.900 ;
        RECT 1444.470 475.700 1444.790 475.760 ;
        RECT 1444.485 434.420 1444.775 434.465 ;
        RECT 1444.930 434.420 1445.250 434.480 ;
        RECT 1444.485 434.280 1445.250 434.420 ;
        RECT 1444.485 434.235 1444.775 434.280 ;
        RECT 1444.930 434.220 1445.250 434.280 ;
        RECT 1444.470 379.680 1444.790 379.740 ;
        RECT 1444.930 379.680 1445.250 379.740 ;
        RECT 1444.470 379.540 1445.250 379.680 ;
        RECT 1444.470 379.480 1444.790 379.540 ;
        RECT 1444.930 379.480 1445.250 379.540 ;
        RECT 1444.470 275.980 1444.790 276.040 ;
        RECT 1444.275 275.840 1444.790 275.980 ;
        RECT 1444.470 275.780 1444.790 275.840 ;
        RECT 1444.470 228.040 1444.790 228.100 ;
        RECT 1444.275 227.900 1444.790 228.040 ;
        RECT 1444.470 227.840 1444.790 227.900 ;
        RECT 1444.930 159.020 1445.250 159.080 ;
        RECT 1444.735 158.880 1445.250 159.020 ;
        RECT 1444.930 158.820 1445.250 158.880 ;
        RECT 1444.930 131.480 1445.250 131.540 ;
        RECT 1444.735 131.340 1445.250 131.480 ;
        RECT 1444.930 131.280 1445.250 131.340 ;
        RECT 1444.010 83.200 1444.330 83.260 ;
        RECT 1444.930 83.200 1445.250 83.260 ;
        RECT 1444.010 83.060 1445.250 83.200 ;
        RECT 1444.010 83.000 1444.330 83.060 ;
        RECT 1444.930 83.000 1445.250 83.060 ;
        RECT 1444.010 36.280 1444.330 36.340 ;
        RECT 1443.815 36.140 1444.330 36.280 ;
        RECT 1444.010 36.080 1444.330 36.140 ;
        RECT 1102.690 27.780 1103.010 27.840 ;
        RECT 1444.025 27.780 1444.315 27.825 ;
        RECT 1102.690 27.640 1444.315 27.780 ;
        RECT 1102.690 27.580 1103.010 27.640 ;
        RECT 1444.025 27.595 1444.315 27.640 ;
      LAYER via ;
        RECT 1444.960 1586.820 1445.220 1587.080 ;
        RECT 1445.420 1545.000 1445.680 1545.260 ;
        RECT 1444.960 1497.400 1445.220 1497.660 ;
        RECT 1445.420 1497.400 1445.680 1497.660 ;
        RECT 1444.960 1463.060 1445.220 1463.320 ;
        RECT 1444.500 1462.380 1444.760 1462.640 ;
        RECT 1444.500 1400.500 1444.760 1400.760 ;
        RECT 1444.960 1400.500 1445.220 1400.760 ;
        RECT 1444.500 1352.560 1444.760 1352.820 ;
        RECT 1444.960 1351.880 1445.220 1352.140 ;
        RECT 1444.500 1248.860 1444.760 1249.120 ;
        RECT 1444.960 1248.860 1445.220 1249.120 ;
        RECT 1444.960 1159.440 1445.220 1159.700 ;
        RECT 1444.500 1159.100 1444.760 1159.360 ;
        RECT 1444.040 1145.160 1444.300 1145.420 ;
        RECT 1444.500 1145.160 1444.760 1145.420 ;
        RECT 1444.960 1096.880 1445.220 1097.140 ;
        RECT 1446.800 1096.880 1447.060 1097.140 ;
        RECT 1446.800 1089.740 1447.060 1090.000 ;
        RECT 1446.800 1048.600 1447.060 1048.860 ;
        RECT 1444.500 862.620 1444.760 862.880 ;
        RECT 1445.420 862.620 1445.680 862.880 ;
        RECT 1444.960 806.860 1445.220 807.120 ;
        RECT 1444.960 783.060 1445.220 783.320 ;
        RECT 1444.960 724.240 1445.220 724.500 ;
        RECT 1445.420 724.240 1445.680 724.500 ;
        RECT 1444.500 675.960 1444.760 676.220 ;
        RECT 1445.420 675.960 1445.680 676.220 ;
        RECT 1445.420 628.020 1445.680 628.280 ;
        RECT 1444.500 620.880 1444.760 621.140 ;
        RECT 1444.500 572.600 1444.760 572.860 ;
        RECT 1445.420 572.600 1445.680 572.860 ;
        RECT 1444.500 475.700 1444.760 475.960 ;
        RECT 1444.960 434.220 1445.220 434.480 ;
        RECT 1444.500 379.480 1444.760 379.740 ;
        RECT 1444.960 379.480 1445.220 379.740 ;
        RECT 1444.500 275.780 1444.760 276.040 ;
        RECT 1444.500 227.840 1444.760 228.100 ;
        RECT 1444.960 158.820 1445.220 159.080 ;
        RECT 1444.960 131.280 1445.220 131.540 ;
        RECT 1444.040 83.000 1444.300 83.260 ;
        RECT 1444.960 83.000 1445.220 83.260 ;
        RECT 1444.040 36.080 1444.300 36.340 ;
        RECT 1102.720 27.580 1102.980 27.840 ;
      LAYER met2 ;
        RECT 1447.710 1700.410 1447.990 1704.000 ;
        RECT 1446.860 1700.270 1447.990 1700.410 ;
        RECT 1446.860 1656.210 1447.000 1700.270 ;
        RECT 1447.710 1700.000 1447.990 1700.270 ;
        RECT 1445.020 1656.070 1447.000 1656.210 ;
        RECT 1445.020 1587.110 1445.160 1656.070 ;
        RECT 1444.960 1586.790 1445.220 1587.110 ;
        RECT 1445.420 1544.970 1445.680 1545.290 ;
        RECT 1445.480 1497.690 1445.620 1544.970 ;
        RECT 1444.960 1497.370 1445.220 1497.690 ;
        RECT 1445.420 1497.370 1445.680 1497.690 ;
        RECT 1445.020 1463.350 1445.160 1497.370 ;
        RECT 1444.960 1463.030 1445.220 1463.350 ;
        RECT 1444.500 1462.350 1444.760 1462.670 ;
        RECT 1444.560 1425.010 1444.700 1462.350 ;
        RECT 1444.560 1424.870 1445.160 1425.010 ;
        RECT 1445.020 1400.790 1445.160 1424.870 ;
        RECT 1444.500 1400.470 1444.760 1400.790 ;
        RECT 1444.960 1400.470 1445.220 1400.790 ;
        RECT 1444.560 1352.850 1444.700 1400.470 ;
        RECT 1444.500 1352.530 1444.760 1352.850 ;
        RECT 1444.960 1351.850 1445.220 1352.170 ;
        RECT 1445.020 1304.650 1445.160 1351.850 ;
        RECT 1444.560 1304.510 1445.160 1304.650 ;
        RECT 1444.560 1249.150 1444.700 1304.510 ;
        RECT 1444.500 1248.830 1444.760 1249.150 ;
        RECT 1444.960 1248.830 1445.220 1249.150 ;
        RECT 1445.020 1159.730 1445.160 1248.830 ;
        RECT 1444.960 1159.410 1445.220 1159.730 ;
        RECT 1444.500 1159.070 1444.760 1159.390 ;
        RECT 1444.560 1145.450 1444.700 1159.070 ;
        RECT 1444.040 1145.130 1444.300 1145.450 ;
        RECT 1444.500 1145.130 1444.760 1145.450 ;
        RECT 1444.100 1097.365 1444.240 1145.130 ;
        RECT 1444.030 1096.995 1444.310 1097.365 ;
        RECT 1444.950 1096.995 1445.230 1097.365 ;
        RECT 1444.960 1096.850 1445.220 1096.995 ;
        RECT 1446.800 1096.850 1447.060 1097.170 ;
        RECT 1446.860 1090.030 1447.000 1096.850 ;
        RECT 1446.800 1089.710 1447.060 1090.030 ;
        RECT 1446.800 1048.570 1447.060 1048.890 ;
        RECT 1446.860 1000.805 1447.000 1048.570 ;
        RECT 1445.410 1000.435 1445.690 1000.805 ;
        RECT 1446.790 1000.435 1447.070 1000.805 ;
        RECT 1445.480 953.205 1445.620 1000.435 ;
        RECT 1445.410 952.835 1445.690 953.205 ;
        RECT 1444.490 952.155 1444.770 952.525 ;
        RECT 1444.560 917.900 1444.700 952.155 ;
        RECT 1444.560 917.760 1445.160 917.900 ;
        RECT 1445.020 883.730 1445.160 917.760 ;
        RECT 1445.020 883.590 1445.620 883.730 ;
        RECT 1445.480 862.910 1445.620 883.590 ;
        RECT 1444.500 862.590 1444.760 862.910 ;
        RECT 1445.420 862.590 1445.680 862.910 ;
        RECT 1444.560 814.370 1444.700 862.590 ;
        RECT 1444.560 814.230 1445.160 814.370 ;
        RECT 1445.020 807.150 1445.160 814.230 ;
        RECT 1444.960 806.830 1445.220 807.150 ;
        RECT 1444.960 783.030 1445.220 783.350 ;
        RECT 1445.020 724.530 1445.160 783.030 ;
        RECT 1444.960 724.210 1445.220 724.530 ;
        RECT 1445.420 724.210 1445.680 724.530 ;
        RECT 1445.480 676.445 1445.620 724.210 ;
        RECT 1444.490 676.075 1444.770 676.445 ;
        RECT 1445.410 676.075 1445.690 676.445 ;
        RECT 1444.500 675.930 1444.760 676.075 ;
        RECT 1445.420 675.930 1445.680 676.075 ;
        RECT 1445.480 628.310 1445.620 675.930 ;
        RECT 1445.420 627.990 1445.680 628.310 ;
        RECT 1444.500 620.850 1444.760 621.170 ;
        RECT 1444.560 572.890 1444.700 620.850 ;
        RECT 1444.500 572.570 1444.760 572.890 ;
        RECT 1445.420 572.570 1445.680 572.890 ;
        RECT 1445.480 537.610 1445.620 572.570 ;
        RECT 1445.480 537.470 1446.080 537.610 ;
        RECT 1445.940 530.810 1446.080 537.470 ;
        RECT 1445.480 530.670 1446.080 530.810 ;
        RECT 1445.480 483.890 1445.620 530.670 ;
        RECT 1445.480 483.750 1446.080 483.890 ;
        RECT 1445.940 476.525 1446.080 483.750 ;
        RECT 1444.950 476.410 1445.230 476.525 ;
        RECT 1444.560 476.270 1445.230 476.410 ;
        RECT 1444.560 475.990 1444.700 476.270 ;
        RECT 1444.950 476.155 1445.230 476.270 ;
        RECT 1445.870 476.155 1446.150 476.525 ;
        RECT 1444.500 475.670 1444.760 475.990 ;
        RECT 1444.960 434.190 1445.220 434.510 ;
        RECT 1445.020 379.770 1445.160 434.190 ;
        RECT 1444.500 379.450 1444.760 379.770 ;
        RECT 1444.960 379.450 1445.220 379.770 ;
        RECT 1444.560 276.070 1444.700 379.450 ;
        RECT 1444.500 275.750 1444.760 276.070 ;
        RECT 1444.500 227.810 1444.760 228.130 ;
        RECT 1444.560 196.250 1444.700 227.810 ;
        RECT 1444.560 196.110 1445.160 196.250 ;
        RECT 1445.020 159.110 1445.160 196.110 ;
        RECT 1444.960 158.790 1445.220 159.110 ;
        RECT 1444.960 131.250 1445.220 131.570 ;
        RECT 1445.020 83.290 1445.160 131.250 ;
        RECT 1444.040 82.970 1444.300 83.290 ;
        RECT 1444.960 82.970 1445.220 83.290 ;
        RECT 1444.100 36.370 1444.240 82.970 ;
        RECT 1444.040 36.050 1444.300 36.370 ;
        RECT 1102.720 27.550 1102.980 27.870 ;
        RECT 1102.780 2.400 1102.920 27.550 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
      LAYER via2 ;
        RECT 1444.030 1097.040 1444.310 1097.320 ;
        RECT 1444.950 1097.040 1445.230 1097.320 ;
        RECT 1445.410 1000.480 1445.690 1000.760 ;
        RECT 1446.790 1000.480 1447.070 1000.760 ;
        RECT 1445.410 952.880 1445.690 953.160 ;
        RECT 1444.490 952.200 1444.770 952.480 ;
        RECT 1444.490 676.120 1444.770 676.400 ;
        RECT 1445.410 676.120 1445.690 676.400 ;
        RECT 1444.950 476.200 1445.230 476.480 ;
        RECT 1445.870 476.200 1446.150 476.480 ;
      LAYER met3 ;
        RECT 1444.005 1097.330 1444.335 1097.345 ;
        RECT 1444.925 1097.330 1445.255 1097.345 ;
        RECT 1444.005 1097.030 1445.255 1097.330 ;
        RECT 1444.005 1097.015 1444.335 1097.030 ;
        RECT 1444.925 1097.015 1445.255 1097.030 ;
        RECT 1445.385 1000.770 1445.715 1000.785 ;
        RECT 1446.765 1000.770 1447.095 1000.785 ;
        RECT 1445.385 1000.470 1447.095 1000.770 ;
        RECT 1445.385 1000.455 1445.715 1000.470 ;
        RECT 1446.765 1000.455 1447.095 1000.470 ;
        RECT 1445.385 953.170 1445.715 953.185 ;
        RECT 1443.790 952.870 1445.715 953.170 ;
        RECT 1443.790 952.490 1444.090 952.870 ;
        RECT 1445.385 952.855 1445.715 952.870 ;
        RECT 1444.465 952.490 1444.795 952.505 ;
        RECT 1443.790 952.190 1444.795 952.490 ;
        RECT 1444.465 952.175 1444.795 952.190 ;
        RECT 1444.465 676.410 1444.795 676.425 ;
        RECT 1445.385 676.410 1445.715 676.425 ;
        RECT 1444.465 676.110 1445.715 676.410 ;
        RECT 1444.465 676.095 1444.795 676.110 ;
        RECT 1445.385 676.095 1445.715 676.110 ;
        RECT 1444.925 476.490 1445.255 476.505 ;
        RECT 1445.845 476.490 1446.175 476.505 ;
        RECT 1444.925 476.190 1446.175 476.490 ;
        RECT 1444.925 476.175 1445.255 476.190 ;
        RECT 1445.845 476.175 1446.175 476.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 0.300 ;
=======
      LAYER li1 ;
        RECT 1450.985 923.525 1451.155 965.855 ;
      LAYER mcon ;
        RECT 1450.985 965.685 1451.155 965.855 ;
      LAYER met1 ;
        RECT 1450.910 965.840 1451.230 965.900 ;
        RECT 1450.715 965.700 1451.230 965.840 ;
        RECT 1450.910 965.640 1451.230 965.700 ;
        RECT 1450.910 923.680 1451.230 923.740 ;
        RECT 1450.715 923.540 1451.230 923.680 ;
        RECT 1450.910 923.480 1451.230 923.540 ;
        RECT 1124.310 48.860 1124.630 48.920 ;
        RECT 1450.910 48.860 1451.230 48.920 ;
        RECT 1124.310 48.720 1451.230 48.860 ;
        RECT 1124.310 48.660 1124.630 48.720 ;
        RECT 1450.910 48.660 1451.230 48.720 ;
      LAYER via ;
        RECT 1450.940 965.640 1451.200 965.900 ;
        RECT 1450.940 923.480 1451.200 923.740 ;
        RECT 1124.340 48.660 1124.600 48.920 ;
        RECT 1450.940 48.660 1451.200 48.920 ;
      LAYER met2 ;
        RECT 1452.310 1700.410 1452.590 1704.000 ;
        RECT 1451.000 1700.270 1452.590 1700.410 ;
        RECT 1451.000 965.930 1451.140 1700.270 ;
        RECT 1452.310 1700.000 1452.590 1700.270 ;
        RECT 1450.940 965.610 1451.200 965.930 ;
        RECT 1450.940 923.450 1451.200 923.770 ;
        RECT 1451.000 48.950 1451.140 923.450 ;
        RECT 1124.340 48.630 1124.600 48.950 ;
        RECT 1450.940 48.630 1451.200 48.950 ;
        RECT 1124.400 16.050 1124.540 48.630 ;
        RECT 1120.720 15.910 1124.540 16.050 ;
        RECT 1120.720 2.400 1120.860 15.910 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1145.010 48.520 1145.330 48.580 ;
        RECT 1457.350 48.520 1457.670 48.580 ;
        RECT 1145.010 48.380 1457.670 48.520 ;
        RECT 1145.010 48.320 1145.330 48.380 ;
        RECT 1457.350 48.320 1457.670 48.380 ;
        RECT 1138.570 13.840 1138.890 13.900 ;
        RECT 1145.010 13.840 1145.330 13.900 ;
        RECT 1138.570 13.700 1145.330 13.840 ;
        RECT 1138.570 13.640 1138.890 13.700 ;
        RECT 1145.010 13.640 1145.330 13.700 ;
      LAYER via ;
        RECT 1145.040 48.320 1145.300 48.580 ;
        RECT 1457.380 48.320 1457.640 48.580 ;
        RECT 1138.600 13.640 1138.860 13.900 ;
        RECT 1145.040 13.640 1145.300 13.900 ;
      LAYER met2 ;
        RECT 1456.910 1700.410 1457.190 1704.000 ;
        RECT 1456.910 1700.270 1457.580 1700.410 ;
        RECT 1456.910 1700.000 1457.190 1700.270 ;
        RECT 1457.440 48.610 1457.580 1700.270 ;
        RECT 1145.040 48.290 1145.300 48.610 ;
        RECT 1457.380 48.290 1457.640 48.610 ;
        RECT 1145.100 13.930 1145.240 48.290 ;
        RECT 1138.600 13.610 1138.860 13.930 ;
        RECT 1145.040 13.610 1145.300 13.930 ;
        RECT 1138.660 2.400 1138.800 13.610 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 0.300 ;
=======
      LAYER met1 ;
        RECT 1455.970 1678.480 1456.290 1678.540 ;
        RECT 1460.570 1678.480 1460.890 1678.540 ;
        RECT 1455.970 1678.340 1460.890 1678.480 ;
        RECT 1455.970 1678.280 1456.290 1678.340 ;
        RECT 1460.570 1678.280 1460.890 1678.340 ;
        RECT 1156.510 24.720 1156.830 24.780 ;
        RECT 1455.970 24.720 1456.290 24.780 ;
        RECT 1156.510 24.580 1456.290 24.720 ;
        RECT 1156.510 24.520 1156.830 24.580 ;
        RECT 1455.970 24.520 1456.290 24.580 ;
      LAYER via ;
        RECT 1456.000 1678.280 1456.260 1678.540 ;
        RECT 1460.600 1678.280 1460.860 1678.540 ;
        RECT 1156.540 24.520 1156.800 24.780 ;
        RECT 1456.000 24.520 1456.260 24.780 ;
      LAYER met2 ;
        RECT 1461.970 1700.410 1462.250 1704.000 ;
        RECT 1460.660 1700.270 1462.250 1700.410 ;
        RECT 1460.660 1678.570 1460.800 1700.270 ;
        RECT 1461.970 1700.000 1462.250 1700.270 ;
        RECT 1456.000 1678.250 1456.260 1678.570 ;
        RECT 1460.600 1678.250 1460.860 1678.570 ;
        RECT 1456.060 24.810 1456.200 1678.250 ;
        RECT 1156.540 24.490 1156.800 24.810 ;
        RECT 1456.000 24.490 1456.260 24.810 ;
        RECT 1156.600 2.400 1156.740 24.490 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 674.310 -4.800 674.870 0.300 ;
=======
        RECT 1331.790 1700.410 1332.070 1704.000 ;
        RECT 1331.790 1700.270 1332.460 1700.410 ;
        RECT 1331.790 1700.000 1332.070 1700.270 ;
        RECT 1332.320 34.525 1332.460 1700.270 ;
        RECT 674.450 34.155 674.730 34.525 ;
        RECT 1332.250 34.155 1332.530 34.525 ;
        RECT 674.520 2.400 674.660 34.155 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 674.450 34.200 674.730 34.480 ;
        RECT 1332.250 34.200 1332.530 34.480 ;
      LAYER met3 ;
        RECT 674.425 34.490 674.755 34.505 ;
        RECT 1332.225 34.490 1332.555 34.505 ;
        RECT 674.425 34.190 1332.555 34.490 ;
        RECT 674.425 34.175 674.755 34.190 ;
        RECT 1332.225 34.175 1332.555 34.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1462.870 1678.140 1463.190 1678.200 ;
        RECT 1465.630 1678.140 1465.950 1678.200 ;
        RECT 1462.870 1678.000 1465.950 1678.140 ;
        RECT 1462.870 1677.940 1463.190 1678.000 ;
        RECT 1465.630 1677.940 1465.950 1678.000 ;
      LAYER via ;
        RECT 1462.900 1677.940 1463.160 1678.200 ;
        RECT 1465.660 1677.940 1465.920 1678.200 ;
      LAYER met2 ;
        RECT 1466.570 1700.410 1466.850 1704.000 ;
        RECT 1465.720 1700.270 1466.850 1700.410 ;
        RECT 1465.720 1678.230 1465.860 1700.270 ;
        RECT 1466.570 1700.000 1466.850 1700.270 ;
        RECT 1462.900 1677.910 1463.160 1678.230 ;
        RECT 1465.660 1677.910 1465.920 1678.230 ;
        RECT 1462.960 17.525 1463.100 1677.910 ;
        RECT 1174.010 17.155 1174.290 17.525 ;
        RECT 1462.890 17.155 1463.170 17.525 ;
        RECT 1174.080 2.400 1174.220 17.155 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
      LAYER via2 ;
        RECT 1174.010 17.200 1174.290 17.480 ;
        RECT 1462.890 17.200 1463.170 17.480 ;
      LAYER met3 ;
        RECT 1173.985 17.490 1174.315 17.505 ;
        RECT 1462.865 17.490 1463.195 17.505 ;
        RECT 1173.985 17.190 1463.195 17.490 ;
        RECT 1173.985 17.175 1174.315 17.190 ;
        RECT 1462.865 17.175 1463.195 17.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1191.810 -4.800 1192.370 0.300 ;
=======
        RECT 1471.630 1700.410 1471.910 1704.000 ;
        RECT 1470.320 1700.270 1471.910 1700.410 ;
        RECT 1470.320 18.205 1470.460 1700.270 ;
        RECT 1471.630 1700.000 1471.910 1700.270 ;
        RECT 1191.950 17.835 1192.230 18.205 ;
        RECT 1470.250 17.835 1470.530 18.205 ;
        RECT 1192.020 2.400 1192.160 17.835 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
      LAYER via2 ;
        RECT 1191.950 17.880 1192.230 18.160 ;
        RECT 1470.250 17.880 1470.530 18.160 ;
      LAYER met3 ;
        RECT 1191.925 18.170 1192.255 18.185 ;
        RECT 1470.225 18.170 1470.555 18.185 ;
        RECT 1191.925 17.870 1470.555 18.170 ;
        RECT 1191.925 17.855 1192.255 17.870 ;
        RECT 1470.225 17.855 1470.555 17.870 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1471.150 1678.480 1471.470 1678.540 ;
        RECT 1475.290 1678.480 1475.610 1678.540 ;
        RECT 1471.150 1678.340 1475.610 1678.480 ;
        RECT 1471.150 1678.280 1471.470 1678.340 ;
        RECT 1475.290 1678.280 1475.610 1678.340 ;
        RECT 1209.870 17.580 1210.190 17.640 ;
        RECT 1471.150 17.580 1471.470 17.640 ;
        RECT 1209.870 17.440 1471.470 17.580 ;
        RECT 1209.870 17.380 1210.190 17.440 ;
        RECT 1471.150 17.380 1471.470 17.440 ;
      LAYER via ;
        RECT 1471.180 1678.280 1471.440 1678.540 ;
        RECT 1475.320 1678.280 1475.580 1678.540 ;
        RECT 1209.900 17.380 1210.160 17.640 ;
        RECT 1471.180 17.380 1471.440 17.640 ;
      LAYER met2 ;
        RECT 1476.230 1700.410 1476.510 1704.000 ;
        RECT 1475.380 1700.270 1476.510 1700.410 ;
        RECT 1475.380 1678.570 1475.520 1700.270 ;
        RECT 1476.230 1700.000 1476.510 1700.270 ;
        RECT 1471.180 1678.250 1471.440 1678.570 ;
        RECT 1475.320 1678.250 1475.580 1678.570 ;
        RECT 1471.240 17.670 1471.380 1678.250 ;
        RECT 1209.900 17.350 1210.160 17.670 ;
        RECT 1471.180 17.350 1471.440 17.670 ;
        RECT 1209.960 2.400 1210.100 17.350 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1477.130 1678.140 1477.450 1678.200 ;
        RECT 1479.890 1678.140 1480.210 1678.200 ;
        RECT 1477.130 1678.000 1480.210 1678.140 ;
        RECT 1477.130 1677.940 1477.450 1678.000 ;
        RECT 1479.890 1677.940 1480.210 1678.000 ;
        RECT 1227.810 18.260 1228.130 18.320 ;
        RECT 1477.130 18.260 1477.450 18.320 ;
        RECT 1227.810 18.120 1423.540 18.260 ;
        RECT 1227.810 18.060 1228.130 18.120 ;
        RECT 1423.400 17.920 1423.540 18.120 ;
        RECT 1464.800 18.120 1477.450 18.260 ;
        RECT 1464.800 17.920 1464.940 18.120 ;
        RECT 1477.130 18.060 1477.450 18.120 ;
        RECT 1423.400 17.780 1464.940 17.920 ;
      LAYER via ;
        RECT 1477.160 1677.940 1477.420 1678.200 ;
        RECT 1479.920 1677.940 1480.180 1678.200 ;
        RECT 1227.840 18.060 1228.100 18.320 ;
        RECT 1477.160 18.060 1477.420 18.320 ;
      LAYER met2 ;
        RECT 1481.290 1700.410 1481.570 1704.000 ;
        RECT 1479.980 1700.270 1481.570 1700.410 ;
        RECT 1479.980 1678.230 1480.120 1700.270 ;
        RECT 1481.290 1700.000 1481.570 1700.270 ;
        RECT 1477.160 1677.910 1477.420 1678.230 ;
        RECT 1479.920 1677.910 1480.180 1678.230 ;
        RECT 1477.220 18.350 1477.360 1677.910 ;
        RECT 1227.840 18.030 1228.100 18.350 ;
        RECT 1477.160 18.030 1477.420 18.350 ;
        RECT 1227.900 2.400 1228.040 18.030 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1245.750 37.980 1246.070 38.040 ;
        RECT 1485.410 37.980 1485.730 38.040 ;
        RECT 1245.750 37.840 1485.730 37.980 ;
        RECT 1245.750 37.780 1246.070 37.840 ;
        RECT 1485.410 37.780 1485.730 37.840 ;
      LAYER via ;
        RECT 1245.780 37.780 1246.040 38.040 ;
        RECT 1485.440 37.780 1485.700 38.040 ;
      LAYER met2 ;
        RECT 1485.890 1700.410 1486.170 1704.000 ;
        RECT 1485.500 1700.270 1486.170 1700.410 ;
        RECT 1485.500 38.070 1485.640 1700.270 ;
        RECT 1485.890 1700.000 1486.170 1700.270 ;
        RECT 1245.780 37.750 1246.040 38.070 ;
        RECT 1485.440 37.750 1485.700 38.070 ;
        RECT 1245.840 2.400 1245.980 37.750 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1263.230 38.320 1263.550 38.380 ;
        RECT 1490.930 38.320 1491.250 38.380 ;
        RECT 1263.230 38.180 1491.250 38.320 ;
        RECT 1263.230 38.120 1263.550 38.180 ;
        RECT 1490.930 38.120 1491.250 38.180 ;
      LAYER via ;
        RECT 1263.260 38.120 1263.520 38.380 ;
        RECT 1490.960 38.120 1491.220 38.380 ;
      LAYER met2 ;
        RECT 1490.950 1700.000 1491.230 1704.000 ;
        RECT 1491.020 38.410 1491.160 1700.000 ;
        RECT 1263.260 38.090 1263.520 38.410 ;
        RECT 1490.960 38.090 1491.220 38.410 ;
        RECT 1263.320 2.400 1263.460 38.090 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1491.390 1678.140 1491.710 1678.200 ;
        RECT 1494.610 1678.140 1494.930 1678.200 ;
        RECT 1491.390 1678.000 1494.930 1678.140 ;
        RECT 1491.390 1677.940 1491.710 1678.000 ;
        RECT 1494.610 1677.940 1494.930 1678.000 ;
        RECT 1281.170 38.660 1281.490 38.720 ;
        RECT 1491.390 38.660 1491.710 38.720 ;
        RECT 1281.170 38.520 1491.710 38.660 ;
        RECT 1281.170 38.460 1281.490 38.520 ;
        RECT 1491.390 38.460 1491.710 38.520 ;
      LAYER via ;
        RECT 1491.420 1677.940 1491.680 1678.200 ;
        RECT 1494.640 1677.940 1494.900 1678.200 ;
        RECT 1281.200 38.460 1281.460 38.720 ;
        RECT 1491.420 38.460 1491.680 38.720 ;
      LAYER met2 ;
        RECT 1495.550 1700.410 1495.830 1704.000 ;
        RECT 1494.700 1700.270 1495.830 1700.410 ;
        RECT 1494.700 1678.230 1494.840 1700.270 ;
        RECT 1495.550 1700.000 1495.830 1700.270 ;
        RECT 1491.420 1677.910 1491.680 1678.230 ;
        RECT 1494.640 1677.910 1494.900 1678.230 ;
        RECT 1491.480 38.750 1491.620 1677.910 ;
        RECT 1281.200 38.430 1281.460 38.750 ;
        RECT 1491.420 38.430 1491.680 38.750 ;
        RECT 1281.260 2.400 1281.400 38.430 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1307.390 1688.000 1307.710 1688.060 ;
        RECT 1500.590 1688.000 1500.910 1688.060 ;
        RECT 1307.390 1687.860 1500.910 1688.000 ;
        RECT 1307.390 1687.800 1307.710 1687.860 ;
        RECT 1500.590 1687.800 1500.910 1687.860 ;
        RECT 1299.110 16.560 1299.430 16.620 ;
        RECT 1306.470 16.560 1306.790 16.620 ;
        RECT 1299.110 16.420 1306.790 16.560 ;
        RECT 1299.110 16.360 1299.430 16.420 ;
        RECT 1306.470 16.360 1306.790 16.420 ;
      LAYER via ;
        RECT 1307.420 1687.800 1307.680 1688.060 ;
        RECT 1500.620 1687.800 1500.880 1688.060 ;
        RECT 1299.140 16.360 1299.400 16.620 ;
        RECT 1306.500 16.360 1306.760 16.620 ;
      LAYER met2 ;
        RECT 1500.610 1700.000 1500.890 1704.000 ;
        RECT 1500.680 1688.090 1500.820 1700.000 ;
        RECT 1307.420 1687.770 1307.680 1688.090 ;
        RECT 1500.620 1687.770 1500.880 1688.090 ;
        RECT 1307.480 34.410 1307.620 1687.770 ;
        RECT 1306.560 34.270 1307.620 34.410 ;
        RECT 1306.560 16.650 1306.700 34.270 ;
        RECT 1299.140 16.330 1299.400 16.650 ;
        RECT 1306.500 16.330 1306.760 16.650 ;
        RECT 1299.200 2.400 1299.340 16.330 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 0.300 ;
=======
      LAYER li1 ;
        RECT 1317.125 1435.225 1317.295 1442.195 ;
        RECT 1317.585 1104.065 1317.755 1189.915 ;
        RECT 1317.585 766.105 1317.755 814.215 ;
        RECT 1317.585 427.805 1317.755 475.915 ;
        RECT 1317.585 372.725 1317.755 420.835 ;
        RECT 1316.665 34.425 1316.835 124.015 ;
      LAYER mcon ;
        RECT 1317.125 1442.025 1317.295 1442.195 ;
        RECT 1317.585 1189.745 1317.755 1189.915 ;
        RECT 1317.585 814.045 1317.755 814.215 ;
        RECT 1317.585 475.745 1317.755 475.915 ;
        RECT 1317.585 420.665 1317.755 420.835 ;
        RECT 1316.665 123.845 1316.835 124.015 ;
      LAYER met1 ;
        RECT 1317.510 1688.340 1317.830 1688.400 ;
        RECT 1505.190 1688.340 1505.510 1688.400 ;
        RECT 1317.510 1688.200 1505.510 1688.340 ;
        RECT 1317.510 1688.140 1317.830 1688.200 ;
        RECT 1505.190 1688.140 1505.510 1688.200 ;
        RECT 1317.050 1642.100 1317.370 1642.160 ;
        RECT 1317.510 1642.100 1317.830 1642.160 ;
        RECT 1317.050 1641.960 1317.830 1642.100 ;
        RECT 1317.050 1641.900 1317.370 1641.960 ;
        RECT 1317.510 1641.900 1317.830 1641.960 ;
        RECT 1316.130 1580.220 1316.450 1580.280 ;
        RECT 1317.510 1580.220 1317.830 1580.280 ;
        RECT 1316.130 1580.080 1317.830 1580.220 ;
        RECT 1316.130 1580.020 1316.450 1580.080 ;
        RECT 1317.510 1580.020 1317.830 1580.080 ;
        RECT 1316.590 1490.800 1316.910 1490.860 ;
        RECT 1317.510 1490.800 1317.830 1490.860 ;
        RECT 1316.590 1490.660 1317.830 1490.800 ;
        RECT 1316.590 1490.600 1316.910 1490.660 ;
        RECT 1317.510 1490.600 1317.830 1490.660 ;
        RECT 1317.050 1442.180 1317.370 1442.240 ;
        RECT 1316.855 1442.040 1317.370 1442.180 ;
        RECT 1317.050 1441.980 1317.370 1442.040 ;
        RECT 1317.050 1435.380 1317.370 1435.440 ;
        RECT 1316.855 1435.240 1317.370 1435.380 ;
        RECT 1317.050 1435.180 1317.370 1435.240 ;
        RECT 1317.050 1393.900 1317.370 1393.960 ;
        RECT 1317.510 1393.900 1317.830 1393.960 ;
        RECT 1317.050 1393.760 1317.830 1393.900 ;
        RECT 1317.050 1393.700 1317.370 1393.760 ;
        RECT 1317.510 1393.700 1317.830 1393.760 ;
        RECT 1316.590 1249.060 1316.910 1249.120 ;
        RECT 1317.510 1249.060 1317.830 1249.120 ;
        RECT 1316.590 1248.920 1317.830 1249.060 ;
        RECT 1316.590 1248.860 1316.910 1248.920 ;
        RECT 1317.510 1248.860 1317.830 1248.920 ;
        RECT 1316.590 1189.900 1316.910 1189.960 ;
        RECT 1317.525 1189.900 1317.815 1189.945 ;
        RECT 1316.590 1189.760 1317.815 1189.900 ;
        RECT 1316.590 1189.700 1316.910 1189.760 ;
        RECT 1317.525 1189.715 1317.815 1189.760 ;
        RECT 1317.510 1104.220 1317.830 1104.280 ;
        RECT 1317.315 1104.080 1317.830 1104.220 ;
        RECT 1317.510 1104.020 1317.830 1104.080 ;
        RECT 1317.050 959.720 1317.370 959.780 ;
        RECT 1317.510 959.720 1317.830 959.780 ;
        RECT 1317.050 959.580 1317.830 959.720 ;
        RECT 1317.050 959.520 1317.370 959.580 ;
        RECT 1317.510 959.520 1317.830 959.580 ;
        RECT 1316.590 959.040 1316.910 959.100 ;
        RECT 1317.510 959.040 1317.830 959.100 ;
        RECT 1316.590 958.900 1317.830 959.040 ;
        RECT 1316.590 958.840 1316.910 958.900 ;
        RECT 1317.510 958.840 1317.830 958.900 ;
        RECT 1316.590 910.760 1316.910 910.820 ;
        RECT 1317.510 910.760 1317.830 910.820 ;
        RECT 1316.590 910.620 1317.830 910.760 ;
        RECT 1316.590 910.560 1316.910 910.620 ;
        RECT 1317.510 910.560 1317.830 910.620 ;
        RECT 1317.050 821.340 1317.370 821.400 ;
        RECT 1317.510 821.340 1317.830 821.400 ;
        RECT 1317.050 821.200 1317.830 821.340 ;
        RECT 1317.050 821.140 1317.370 821.200 ;
        RECT 1317.510 821.140 1317.830 821.200 ;
        RECT 1317.510 814.200 1317.830 814.260 ;
        RECT 1317.315 814.060 1317.830 814.200 ;
        RECT 1317.510 814.000 1317.830 814.060 ;
        RECT 1317.510 766.260 1317.830 766.320 ;
        RECT 1317.315 766.120 1317.830 766.260 ;
        RECT 1317.510 766.060 1317.830 766.120 ;
        RECT 1316.590 717.640 1316.910 717.700 ;
        RECT 1317.510 717.640 1317.830 717.700 ;
        RECT 1316.590 717.500 1317.830 717.640 ;
        RECT 1316.590 717.440 1316.910 717.500 ;
        RECT 1317.510 717.440 1317.830 717.500 ;
        RECT 1317.510 475.900 1317.830 475.960 ;
        RECT 1317.315 475.760 1317.830 475.900 ;
        RECT 1317.510 475.700 1317.830 475.760 ;
        RECT 1317.510 427.960 1317.830 428.020 ;
        RECT 1317.315 427.820 1317.830 427.960 ;
        RECT 1317.510 427.760 1317.830 427.820 ;
        RECT 1317.510 420.820 1317.830 420.880 ;
        RECT 1317.315 420.680 1317.830 420.820 ;
        RECT 1317.510 420.620 1317.830 420.680 ;
        RECT 1317.510 372.880 1317.830 372.940 ;
        RECT 1317.315 372.740 1317.830 372.880 ;
        RECT 1317.510 372.680 1317.830 372.740 ;
        RECT 1317.510 331.740 1317.830 331.800 ;
        RECT 1317.140 331.600 1317.830 331.740 ;
        RECT 1317.140 331.460 1317.280 331.600 ;
        RECT 1317.510 331.540 1317.830 331.600 ;
        RECT 1317.050 331.200 1317.370 331.460 ;
        RECT 1317.050 283.120 1317.370 283.180 ;
        RECT 1317.510 283.120 1317.830 283.180 ;
        RECT 1317.050 282.980 1317.830 283.120 ;
        RECT 1317.050 282.920 1317.370 282.980 ;
        RECT 1317.510 282.920 1317.830 282.980 ;
        RECT 1317.050 234.840 1317.370 234.900 ;
        RECT 1317.510 234.840 1317.830 234.900 ;
        RECT 1317.050 234.700 1317.830 234.840 ;
        RECT 1317.050 234.640 1317.370 234.700 ;
        RECT 1317.510 234.640 1317.830 234.700 ;
        RECT 1317.050 186.560 1317.370 186.620 ;
        RECT 1317.510 186.560 1317.830 186.620 ;
        RECT 1317.050 186.420 1317.830 186.560 ;
        RECT 1317.050 186.360 1317.370 186.420 ;
        RECT 1317.510 186.360 1317.830 186.420 ;
        RECT 1316.590 131.140 1316.910 131.200 ;
        RECT 1317.510 131.140 1317.830 131.200 ;
        RECT 1316.590 131.000 1317.830 131.140 ;
        RECT 1316.590 130.940 1316.910 131.000 ;
        RECT 1317.510 130.940 1317.830 131.000 ;
        RECT 1316.590 124.000 1316.910 124.060 ;
        RECT 1316.395 123.860 1316.910 124.000 ;
        RECT 1316.590 123.800 1316.910 123.860 ;
        RECT 1316.605 34.580 1316.895 34.625 ;
        RECT 1317.050 34.580 1317.370 34.640 ;
        RECT 1316.605 34.440 1317.370 34.580 ;
        RECT 1316.605 34.395 1316.895 34.440 ;
        RECT 1317.050 34.380 1317.370 34.440 ;
      LAYER via ;
        RECT 1317.540 1688.140 1317.800 1688.400 ;
        RECT 1505.220 1688.140 1505.480 1688.400 ;
        RECT 1317.080 1641.900 1317.340 1642.160 ;
        RECT 1317.540 1641.900 1317.800 1642.160 ;
        RECT 1316.160 1580.020 1316.420 1580.280 ;
        RECT 1317.540 1580.020 1317.800 1580.280 ;
        RECT 1316.620 1490.600 1316.880 1490.860 ;
        RECT 1317.540 1490.600 1317.800 1490.860 ;
        RECT 1317.080 1441.980 1317.340 1442.240 ;
        RECT 1317.080 1435.180 1317.340 1435.440 ;
        RECT 1317.080 1393.700 1317.340 1393.960 ;
        RECT 1317.540 1393.700 1317.800 1393.960 ;
        RECT 1316.620 1248.860 1316.880 1249.120 ;
        RECT 1317.540 1248.860 1317.800 1249.120 ;
        RECT 1316.620 1189.700 1316.880 1189.960 ;
        RECT 1317.540 1104.020 1317.800 1104.280 ;
        RECT 1317.080 959.520 1317.340 959.780 ;
        RECT 1317.540 959.520 1317.800 959.780 ;
        RECT 1316.620 958.840 1316.880 959.100 ;
        RECT 1317.540 958.840 1317.800 959.100 ;
        RECT 1316.620 910.560 1316.880 910.820 ;
        RECT 1317.540 910.560 1317.800 910.820 ;
        RECT 1317.080 821.140 1317.340 821.400 ;
        RECT 1317.540 821.140 1317.800 821.400 ;
        RECT 1317.540 814.000 1317.800 814.260 ;
        RECT 1317.540 766.060 1317.800 766.320 ;
        RECT 1316.620 717.440 1316.880 717.700 ;
        RECT 1317.540 717.440 1317.800 717.700 ;
        RECT 1317.540 475.700 1317.800 475.960 ;
        RECT 1317.540 427.760 1317.800 428.020 ;
        RECT 1317.540 420.620 1317.800 420.880 ;
        RECT 1317.540 372.680 1317.800 372.940 ;
        RECT 1317.540 331.540 1317.800 331.800 ;
        RECT 1317.080 331.200 1317.340 331.460 ;
        RECT 1317.080 282.920 1317.340 283.180 ;
        RECT 1317.540 282.920 1317.800 283.180 ;
        RECT 1317.080 234.640 1317.340 234.900 ;
        RECT 1317.540 234.640 1317.800 234.900 ;
        RECT 1317.080 186.360 1317.340 186.620 ;
        RECT 1317.540 186.360 1317.800 186.620 ;
        RECT 1316.620 130.940 1316.880 131.200 ;
        RECT 1317.540 130.940 1317.800 131.200 ;
        RECT 1316.620 123.800 1316.880 124.060 ;
        RECT 1317.080 34.380 1317.340 34.640 ;
      LAYER met2 ;
        RECT 1505.210 1700.000 1505.490 1704.000 ;
        RECT 1505.280 1688.430 1505.420 1700.000 ;
        RECT 1317.540 1688.110 1317.800 1688.430 ;
        RECT 1505.220 1688.110 1505.480 1688.430 ;
        RECT 1317.600 1642.190 1317.740 1688.110 ;
        RECT 1317.080 1641.870 1317.340 1642.190 ;
        RECT 1317.540 1641.870 1317.800 1642.190 ;
        RECT 1317.140 1628.445 1317.280 1641.870 ;
        RECT 1316.150 1628.075 1316.430 1628.445 ;
        RECT 1317.070 1628.075 1317.350 1628.445 ;
        RECT 1316.220 1580.310 1316.360 1628.075 ;
        RECT 1316.160 1579.990 1316.420 1580.310 ;
        RECT 1317.540 1579.990 1317.800 1580.310 ;
        RECT 1317.600 1538.570 1317.740 1579.990 ;
        RECT 1316.680 1538.430 1317.740 1538.570 ;
        RECT 1316.680 1490.890 1316.820 1538.430 ;
        RECT 1316.620 1490.570 1316.880 1490.890 ;
        RECT 1317.540 1490.570 1317.800 1490.890 ;
        RECT 1317.600 1483.490 1317.740 1490.570 ;
        RECT 1317.140 1483.350 1317.740 1483.490 ;
        RECT 1317.140 1442.270 1317.280 1483.350 ;
        RECT 1317.080 1441.950 1317.340 1442.270 ;
        RECT 1317.080 1435.150 1317.340 1435.470 ;
        RECT 1317.140 1393.990 1317.280 1435.150 ;
        RECT 1317.080 1393.670 1317.340 1393.990 ;
        RECT 1317.540 1393.670 1317.800 1393.990 ;
        RECT 1317.600 1297.285 1317.740 1393.670 ;
        RECT 1316.610 1296.915 1316.890 1297.285 ;
        RECT 1317.530 1296.915 1317.810 1297.285 ;
        RECT 1316.680 1249.150 1316.820 1296.915 ;
        RECT 1316.620 1248.830 1316.880 1249.150 ;
        RECT 1317.540 1248.830 1317.800 1249.150 ;
        RECT 1317.600 1200.725 1317.740 1248.830 ;
        RECT 1316.610 1200.355 1316.890 1200.725 ;
        RECT 1317.530 1200.355 1317.810 1200.725 ;
        RECT 1316.680 1189.990 1316.820 1200.355 ;
        RECT 1316.620 1189.670 1316.880 1189.990 ;
        RECT 1317.540 1103.990 1317.800 1104.310 ;
        RECT 1317.600 1048.970 1317.740 1103.990 ;
        RECT 1317.140 1048.830 1317.740 1048.970 ;
        RECT 1317.140 1007.605 1317.280 1048.830 ;
        RECT 1317.070 1007.235 1317.350 1007.605 ;
        RECT 1317.070 1006.555 1317.350 1006.925 ;
        RECT 1317.140 959.810 1317.280 1006.555 ;
        RECT 1317.080 959.490 1317.340 959.810 ;
        RECT 1317.540 959.490 1317.800 959.810 ;
        RECT 1317.600 959.130 1317.740 959.490 ;
        RECT 1316.620 958.810 1316.880 959.130 ;
        RECT 1317.540 958.810 1317.800 959.130 ;
        RECT 1316.680 911.045 1316.820 958.810 ;
        RECT 1316.610 910.675 1316.890 911.045 ;
        RECT 1317.530 910.675 1317.810 911.045 ;
        RECT 1316.620 910.530 1316.880 910.675 ;
        RECT 1317.540 910.530 1317.800 910.675 ;
        RECT 1316.680 886.450 1316.820 910.530 ;
        RECT 1316.680 886.310 1317.280 886.450 ;
        RECT 1317.140 821.430 1317.280 886.310 ;
        RECT 1317.080 821.110 1317.340 821.430 ;
        RECT 1317.540 821.110 1317.800 821.430 ;
        RECT 1317.600 814.290 1317.740 821.110 ;
        RECT 1317.540 813.970 1317.800 814.290 ;
        RECT 1317.540 766.030 1317.800 766.350 ;
        RECT 1317.600 717.730 1317.740 766.030 ;
        RECT 1316.620 717.410 1316.880 717.730 ;
        RECT 1317.540 717.410 1317.800 717.730 ;
        RECT 1316.680 669.645 1316.820 717.410 ;
        RECT 1316.610 669.275 1316.890 669.645 ;
        RECT 1317.530 669.275 1317.810 669.645 ;
        RECT 1317.600 475.990 1317.740 669.275 ;
        RECT 1317.540 475.670 1317.800 475.990 ;
        RECT 1317.540 427.730 1317.800 428.050 ;
        RECT 1317.600 420.910 1317.740 427.730 ;
        RECT 1317.540 420.590 1317.800 420.910 ;
        RECT 1317.540 372.650 1317.800 372.970 ;
        RECT 1317.600 331.830 1317.740 372.650 ;
        RECT 1317.540 331.510 1317.800 331.830 ;
        RECT 1317.080 331.170 1317.340 331.490 ;
        RECT 1317.140 283.210 1317.280 331.170 ;
        RECT 1317.080 282.890 1317.340 283.210 ;
        RECT 1317.540 282.890 1317.800 283.210 ;
        RECT 1317.600 234.930 1317.740 282.890 ;
        RECT 1317.080 234.610 1317.340 234.930 ;
        RECT 1317.540 234.610 1317.800 234.930 ;
        RECT 1317.140 186.650 1317.280 234.610 ;
        RECT 1317.080 186.330 1317.340 186.650 ;
        RECT 1317.540 186.330 1317.800 186.650 ;
        RECT 1317.600 131.230 1317.740 186.330 ;
        RECT 1316.620 130.910 1316.880 131.230 ;
        RECT 1317.540 130.910 1317.800 131.230 ;
        RECT 1316.680 124.090 1316.820 130.910 ;
        RECT 1316.620 123.770 1316.880 124.090 ;
        RECT 1317.080 34.350 1317.340 34.670 ;
        RECT 1317.140 2.400 1317.280 34.350 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
      LAYER via2 ;
        RECT 1316.150 1628.120 1316.430 1628.400 ;
        RECT 1317.070 1628.120 1317.350 1628.400 ;
        RECT 1316.610 1296.960 1316.890 1297.240 ;
        RECT 1317.530 1296.960 1317.810 1297.240 ;
        RECT 1316.610 1200.400 1316.890 1200.680 ;
        RECT 1317.530 1200.400 1317.810 1200.680 ;
        RECT 1317.070 1007.280 1317.350 1007.560 ;
        RECT 1317.070 1006.600 1317.350 1006.880 ;
        RECT 1316.610 910.720 1316.890 911.000 ;
        RECT 1317.530 910.720 1317.810 911.000 ;
        RECT 1316.610 669.320 1316.890 669.600 ;
        RECT 1317.530 669.320 1317.810 669.600 ;
      LAYER met3 ;
        RECT 1316.125 1628.410 1316.455 1628.425 ;
        RECT 1317.045 1628.410 1317.375 1628.425 ;
        RECT 1316.125 1628.110 1317.375 1628.410 ;
        RECT 1316.125 1628.095 1316.455 1628.110 ;
        RECT 1317.045 1628.095 1317.375 1628.110 ;
        RECT 1316.585 1297.250 1316.915 1297.265 ;
        RECT 1317.505 1297.250 1317.835 1297.265 ;
        RECT 1316.585 1296.950 1317.835 1297.250 ;
        RECT 1316.585 1296.935 1316.915 1296.950 ;
        RECT 1317.505 1296.935 1317.835 1296.950 ;
        RECT 1316.585 1200.690 1316.915 1200.705 ;
        RECT 1317.505 1200.690 1317.835 1200.705 ;
        RECT 1316.585 1200.390 1317.835 1200.690 ;
        RECT 1316.585 1200.375 1316.915 1200.390 ;
        RECT 1317.505 1200.375 1317.835 1200.390 ;
        RECT 1317.045 1007.570 1317.375 1007.585 ;
        RECT 1317.045 1007.270 1318.050 1007.570 ;
        RECT 1317.045 1007.255 1317.375 1007.270 ;
        RECT 1317.045 1006.890 1317.375 1006.905 ;
        RECT 1317.750 1006.890 1318.050 1007.270 ;
        RECT 1317.045 1006.590 1318.050 1006.890 ;
        RECT 1317.045 1006.575 1317.375 1006.590 ;
        RECT 1316.585 911.010 1316.915 911.025 ;
        RECT 1317.505 911.010 1317.835 911.025 ;
        RECT 1316.585 910.710 1317.835 911.010 ;
        RECT 1316.585 910.695 1316.915 910.710 ;
        RECT 1317.505 910.695 1317.835 910.710 ;
        RECT 1316.585 669.610 1316.915 669.625 ;
        RECT 1317.505 669.610 1317.835 669.625 ;
        RECT 1316.585 669.310 1317.835 669.610 ;
        RECT 1316.585 669.295 1316.915 669.310 ;
        RECT 1317.505 669.295 1317.835 669.310 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1338.210 1689.360 1338.530 1689.420 ;
        RECT 1510.250 1689.360 1510.570 1689.420 ;
        RECT 1338.210 1689.220 1510.570 1689.360 ;
        RECT 1338.210 1689.160 1338.530 1689.220 ;
        RECT 1510.250 1689.160 1510.570 1689.220 ;
        RECT 1334.990 20.640 1335.310 20.700 ;
        RECT 1338.210 20.640 1338.530 20.700 ;
        RECT 1334.990 20.500 1338.530 20.640 ;
        RECT 1334.990 20.440 1335.310 20.500 ;
        RECT 1338.210 20.440 1338.530 20.500 ;
      LAYER via ;
        RECT 1338.240 1689.160 1338.500 1689.420 ;
        RECT 1510.280 1689.160 1510.540 1689.420 ;
        RECT 1335.020 20.440 1335.280 20.700 ;
        RECT 1338.240 20.440 1338.500 20.700 ;
      LAYER met2 ;
        RECT 1510.270 1700.000 1510.550 1704.000 ;
        RECT 1510.340 1689.450 1510.480 1700.000 ;
        RECT 1338.240 1689.130 1338.500 1689.450 ;
        RECT 1510.280 1689.130 1510.540 1689.450 ;
        RECT 1338.300 20.730 1338.440 1689.130 ;
        RECT 1335.020 20.410 1335.280 20.730 ;
        RECT 1338.240 20.410 1338.500 20.730 ;
        RECT 1335.080 2.400 1335.220 20.410 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1335.910 1642.780 1336.230 1642.840 ;
        RECT 1335.080 1642.640 1336.230 1642.780 ;
        RECT 1335.080 1642.500 1335.220 1642.640 ;
        RECT 1335.910 1642.580 1336.230 1642.640 ;
        RECT 1334.990 1642.240 1335.310 1642.500 ;
        RECT 696.510 54.640 696.830 54.700 ;
        RECT 1334.990 54.640 1335.310 54.700 ;
        RECT 696.510 54.500 1335.310 54.640 ;
        RECT 696.510 54.440 696.830 54.500 ;
        RECT 1334.990 54.440 1335.310 54.500 ;
      LAYER via ;
        RECT 1335.940 1642.580 1336.200 1642.840 ;
        RECT 1335.020 1642.240 1335.280 1642.500 ;
        RECT 696.540 54.440 696.800 54.700 ;
        RECT 1335.020 54.440 1335.280 54.700 ;
      LAYER met2 ;
        RECT 1336.850 1700.410 1337.130 1704.000 ;
        RECT 1336.000 1700.270 1337.130 1700.410 ;
        RECT 1336.000 1642.870 1336.140 1700.270 ;
        RECT 1336.850 1700.000 1337.130 1700.270 ;
        RECT 1335.940 1642.550 1336.200 1642.870 ;
        RECT 1335.020 1642.210 1335.280 1642.530 ;
        RECT 1335.080 54.730 1335.220 1642.210 ;
        RECT 696.540 54.410 696.800 54.730 ;
        RECT 1335.020 54.410 1335.280 54.730 ;
        RECT 696.600 17.410 696.740 54.410 ;
        RECT 692.460 17.270 696.740 17.410 ;
        RECT 692.460 2.400 692.600 17.270 ;
        RECT 692.250 -4.800 692.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 0.300 ;
=======
      LAYER li1 ;
        RECT 1410.965 16.065 1411.135 20.315 ;
      LAYER mcon ;
        RECT 1410.965 20.145 1411.135 20.315 ;
      LAYER met1 ;
        RECT 1410.905 20.300 1411.195 20.345 ;
        RECT 1512.090 20.300 1512.410 20.360 ;
        RECT 1410.905 20.160 1512.410 20.300 ;
        RECT 1410.905 20.115 1411.195 20.160 ;
        RECT 1512.090 20.100 1512.410 20.160 ;
        RECT 1352.470 16.220 1352.790 16.280 ;
        RECT 1410.905 16.220 1411.195 16.265 ;
        RECT 1352.470 16.080 1411.195 16.220 ;
        RECT 1352.470 16.020 1352.790 16.080 ;
        RECT 1410.905 16.035 1411.195 16.080 ;
      LAYER via ;
        RECT 1512.120 20.100 1512.380 20.360 ;
        RECT 1352.500 16.020 1352.760 16.280 ;
      LAYER met2 ;
        RECT 1514.870 1700.410 1515.150 1704.000 ;
        RECT 1514.020 1700.270 1515.150 1700.410 ;
        RECT 1514.020 1675.930 1514.160 1700.270 ;
        RECT 1514.870 1700.000 1515.150 1700.270 ;
        RECT 1512.640 1675.790 1514.160 1675.930 ;
        RECT 1512.640 20.810 1512.780 1675.790 ;
        RECT 1512.180 20.670 1512.780 20.810 ;
        RECT 1512.180 20.390 1512.320 20.670 ;
        RECT 1512.120 20.070 1512.380 20.390 ;
        RECT 1352.500 15.990 1352.760 16.310 ;
        RECT 1352.560 2.400 1352.700 15.990 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1393.960 20.500 1512.780 20.640 ;
        RECT 1370.410 20.300 1370.730 20.360 ;
        RECT 1393.960 20.300 1394.100 20.500 ;
        RECT 1370.410 20.160 1394.100 20.300 ;
        RECT 1512.640 20.300 1512.780 20.500 ;
        RECT 1519.450 20.300 1519.770 20.360 ;
        RECT 1512.640 20.160 1519.770 20.300 ;
        RECT 1370.410 20.100 1370.730 20.160 ;
        RECT 1519.450 20.100 1519.770 20.160 ;
      LAYER via ;
        RECT 1370.440 20.100 1370.700 20.360 ;
        RECT 1519.480 20.100 1519.740 20.360 ;
      LAYER met2 ;
        RECT 1519.930 1700.410 1520.210 1704.000 ;
        RECT 1519.540 1700.270 1520.210 1700.410 ;
        RECT 1519.540 20.390 1519.680 1700.270 ;
        RECT 1519.930 1700.000 1520.210 1700.270 ;
        RECT 1370.440 20.070 1370.700 20.390 ;
        RECT 1519.480 20.070 1519.740 20.390 ;
        RECT 1370.500 2.400 1370.640 20.070 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 0.300 ;
=======
      LAYER li1 ;
        RECT 1438.105 15.045 1438.275 16.575 ;
        RECT 1486.405 16.405 1486.575 18.955 ;
      LAYER mcon ;
        RECT 1486.405 18.785 1486.575 18.955 ;
        RECT 1438.105 16.405 1438.275 16.575 ;
      LAYER met1 ;
        RECT 1518.990 1678.140 1519.310 1678.200 ;
        RECT 1523.590 1678.140 1523.910 1678.200 ;
        RECT 1518.990 1678.000 1523.910 1678.140 ;
        RECT 1518.990 1677.940 1519.310 1678.000 ;
        RECT 1523.590 1677.940 1523.910 1678.000 ;
        RECT 1486.345 18.940 1486.635 18.985 ;
        RECT 1518.530 18.940 1518.850 19.000 ;
        RECT 1486.345 18.800 1518.850 18.940 ;
        RECT 1486.345 18.755 1486.635 18.800 ;
        RECT 1518.530 18.740 1518.850 18.800 ;
        RECT 1438.045 16.560 1438.335 16.605 ;
        RECT 1486.345 16.560 1486.635 16.605 ;
        RECT 1438.045 16.420 1486.635 16.560 ;
        RECT 1438.045 16.375 1438.335 16.420 ;
        RECT 1486.345 16.375 1486.635 16.420 ;
        RECT 1388.350 15.200 1388.670 15.260 ;
        RECT 1438.045 15.200 1438.335 15.245 ;
        RECT 1388.350 15.060 1438.335 15.200 ;
        RECT 1388.350 15.000 1388.670 15.060 ;
        RECT 1438.045 15.015 1438.335 15.060 ;
      LAYER via ;
        RECT 1519.020 1677.940 1519.280 1678.200 ;
        RECT 1523.620 1677.940 1523.880 1678.200 ;
        RECT 1518.560 18.740 1518.820 19.000 ;
        RECT 1388.380 15.000 1388.640 15.260 ;
      LAYER met2 ;
        RECT 1524.530 1700.410 1524.810 1704.000 ;
        RECT 1523.680 1700.270 1524.810 1700.410 ;
        RECT 1523.680 1678.230 1523.820 1700.270 ;
        RECT 1524.530 1700.000 1524.810 1700.270 ;
        RECT 1519.020 1677.910 1519.280 1678.230 ;
        RECT 1523.620 1677.910 1523.880 1678.230 ;
        RECT 1519.080 20.130 1519.220 1677.910 ;
        RECT 1518.620 19.990 1519.220 20.130 ;
        RECT 1518.620 19.030 1518.760 19.990 ;
        RECT 1518.560 18.710 1518.820 19.030 ;
        RECT 1388.380 14.970 1388.640 15.290 ;
        RECT 1388.440 2.400 1388.580 14.970 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 0.300 ;
=======
      LAYER li1 ;
        RECT 1479.505 1684.445 1479.675 1685.635 ;
      LAYER mcon ;
        RECT 1479.505 1685.465 1479.675 1685.635 ;
      LAYER met1 ;
        RECT 1407.210 1685.620 1407.530 1685.680 ;
        RECT 1479.445 1685.620 1479.735 1685.665 ;
        RECT 1407.210 1685.480 1479.735 1685.620 ;
        RECT 1407.210 1685.420 1407.530 1685.480 ;
        RECT 1479.445 1685.435 1479.735 1685.480 ;
        RECT 1479.445 1684.600 1479.735 1684.645 ;
        RECT 1529.570 1684.600 1529.890 1684.660 ;
        RECT 1479.445 1684.460 1529.890 1684.600 ;
        RECT 1479.445 1684.415 1479.735 1684.460 ;
        RECT 1529.570 1684.400 1529.890 1684.460 ;
        RECT 1406.290 2.960 1406.610 3.020 ;
        RECT 1407.210 2.960 1407.530 3.020 ;
        RECT 1406.290 2.820 1407.530 2.960 ;
        RECT 1406.290 2.760 1406.610 2.820 ;
        RECT 1407.210 2.760 1407.530 2.820 ;
      LAYER via ;
        RECT 1407.240 1685.420 1407.500 1685.680 ;
        RECT 1529.600 1684.400 1529.860 1684.660 ;
        RECT 1406.320 2.760 1406.580 3.020 ;
        RECT 1407.240 2.760 1407.500 3.020 ;
      LAYER met2 ;
        RECT 1529.590 1700.000 1529.870 1704.000 ;
        RECT 1407.240 1685.390 1407.500 1685.710 ;
        RECT 1407.300 3.050 1407.440 1685.390 ;
        RECT 1529.660 1684.690 1529.800 1700.000 ;
        RECT 1529.600 1684.370 1529.860 1684.690 ;
        RECT 1406.320 2.730 1406.580 3.050 ;
        RECT 1407.240 2.730 1407.500 3.050 ;
        RECT 1406.380 2.400 1406.520 2.730 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 0.300 ;
=======
      LAYER met1 ;
        RECT 1427.910 1685.280 1428.230 1685.340 ;
        RECT 1534.170 1685.280 1534.490 1685.340 ;
        RECT 1427.910 1685.140 1534.490 1685.280 ;
        RECT 1427.910 1685.080 1428.230 1685.140 ;
        RECT 1534.170 1685.080 1534.490 1685.140 ;
        RECT 1427.910 318.960 1428.230 319.220 ;
        RECT 1428.000 318.540 1428.140 318.960 ;
        RECT 1427.910 318.280 1428.230 318.540 ;
        RECT 1423.770 18.260 1424.090 18.320 ;
        RECT 1427.910 18.260 1428.230 18.320 ;
        RECT 1423.770 18.120 1428.230 18.260 ;
        RECT 1423.770 18.060 1424.090 18.120 ;
        RECT 1427.910 18.060 1428.230 18.120 ;
      LAYER via ;
        RECT 1427.940 1685.080 1428.200 1685.340 ;
        RECT 1534.200 1685.080 1534.460 1685.340 ;
        RECT 1427.940 318.960 1428.200 319.220 ;
        RECT 1427.940 318.280 1428.200 318.540 ;
        RECT 1423.800 18.060 1424.060 18.320 ;
        RECT 1427.940 18.060 1428.200 18.320 ;
      LAYER met2 ;
        RECT 1534.190 1700.000 1534.470 1704.000 ;
        RECT 1534.260 1685.370 1534.400 1700.000 ;
        RECT 1427.940 1685.050 1428.200 1685.370 ;
        RECT 1534.200 1685.050 1534.460 1685.370 ;
        RECT 1428.000 319.250 1428.140 1685.050 ;
        RECT 1427.940 318.930 1428.200 319.250 ;
        RECT 1427.940 318.250 1428.200 318.570 ;
        RECT 1428.000 18.350 1428.140 318.250 ;
        RECT 1423.800 18.030 1424.060 18.350 ;
        RECT 1427.940 18.030 1428.200 18.350 ;
        RECT 1423.860 2.400 1424.000 18.030 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 0.300 ;
=======
      LAYER met1 ;
        RECT 1441.710 1684.940 1442.030 1685.000 ;
        RECT 1539.230 1684.940 1539.550 1685.000 ;
        RECT 1441.710 1684.800 1539.550 1684.940 ;
        RECT 1441.710 1684.740 1442.030 1684.800 ;
        RECT 1539.230 1684.740 1539.550 1684.800 ;
      LAYER via ;
        RECT 1441.740 1684.740 1442.000 1685.000 ;
        RECT 1539.260 1684.740 1539.520 1685.000 ;
      LAYER met2 ;
        RECT 1539.250 1700.000 1539.530 1704.000 ;
        RECT 1539.320 1685.030 1539.460 1700.000 ;
        RECT 1441.740 1684.710 1442.000 1685.030 ;
        RECT 1539.260 1684.710 1539.520 1685.030 ;
        RECT 1441.800 2.400 1441.940 1684.710 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1539.690 1669.640 1540.010 1669.700 ;
        RECT 1542.910 1669.640 1543.230 1669.700 ;
        RECT 1539.690 1669.500 1543.230 1669.640 ;
        RECT 1539.690 1669.440 1540.010 1669.500 ;
        RECT 1542.910 1669.440 1543.230 1669.500 ;
        RECT 1459.650 14.520 1459.970 14.580 ;
        RECT 1539.690 14.520 1540.010 14.580 ;
        RECT 1459.650 14.380 1540.010 14.520 ;
        RECT 1459.650 14.320 1459.970 14.380 ;
        RECT 1539.690 14.320 1540.010 14.380 ;
      LAYER via ;
        RECT 1539.720 1669.440 1539.980 1669.700 ;
        RECT 1542.940 1669.440 1543.200 1669.700 ;
        RECT 1459.680 14.320 1459.940 14.580 ;
        RECT 1539.720 14.320 1539.980 14.580 ;
      LAYER met2 ;
        RECT 1543.850 1700.410 1544.130 1704.000 ;
        RECT 1543.000 1700.270 1544.130 1700.410 ;
        RECT 1543.000 1669.730 1543.140 1700.270 ;
        RECT 1543.850 1700.000 1544.130 1700.270 ;
        RECT 1539.720 1669.410 1539.980 1669.730 ;
        RECT 1542.940 1669.410 1543.200 1669.730 ;
        RECT 1539.780 14.610 1539.920 1669.410 ;
        RECT 1459.680 14.290 1459.940 14.610 ;
        RECT 1539.720 14.290 1539.980 14.610 ;
        RECT 1459.740 2.400 1459.880 14.290 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1477.590 17.580 1477.910 17.640 ;
        RECT 1547.510 17.580 1547.830 17.640 ;
        RECT 1477.590 17.440 1547.830 17.580 ;
        RECT 1477.590 17.380 1477.910 17.440 ;
        RECT 1547.510 17.380 1547.830 17.440 ;
      LAYER via ;
        RECT 1477.620 17.380 1477.880 17.640 ;
        RECT 1547.540 17.380 1547.800 17.640 ;
      LAYER met2 ;
        RECT 1548.910 1700.410 1549.190 1704.000 ;
        RECT 1547.600 1700.270 1549.190 1700.410 ;
        RECT 1547.600 17.670 1547.740 1700.270 ;
        RECT 1548.910 1700.000 1549.190 1700.270 ;
        RECT 1477.620 17.350 1477.880 17.670 ;
        RECT 1547.540 17.350 1547.800 17.670 ;
        RECT 1477.680 2.400 1477.820 17.350 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 0.300 ;
=======
      LAYER li1 ;
        RECT 1514.465 1655.545 1514.635 1687.675 ;
      LAYER mcon ;
        RECT 1514.465 1687.505 1514.635 1687.675 ;
      LAYER met1 ;
        RECT 1514.405 1687.660 1514.695 1687.705 ;
        RECT 1553.490 1687.660 1553.810 1687.720 ;
        RECT 1514.405 1687.520 1553.810 1687.660 ;
        RECT 1514.405 1687.475 1514.695 1687.520 ;
        RECT 1553.490 1687.460 1553.810 1687.520 ;
        RECT 1514.390 1655.700 1514.710 1655.760 ;
        RECT 1514.195 1655.560 1514.710 1655.700 ;
        RECT 1514.390 1655.500 1514.710 1655.560 ;
        RECT 1495.530 16.220 1495.850 16.280 ;
        RECT 1514.390 16.220 1514.710 16.280 ;
        RECT 1495.530 16.080 1514.710 16.220 ;
        RECT 1495.530 16.020 1495.850 16.080 ;
        RECT 1514.390 16.020 1514.710 16.080 ;
      LAYER via ;
        RECT 1553.520 1687.460 1553.780 1687.720 ;
        RECT 1514.420 1655.500 1514.680 1655.760 ;
        RECT 1495.560 16.020 1495.820 16.280 ;
        RECT 1514.420 16.020 1514.680 16.280 ;
      LAYER met2 ;
        RECT 1553.510 1700.000 1553.790 1704.000 ;
        RECT 1553.580 1687.750 1553.720 1700.000 ;
        RECT 1553.520 1687.430 1553.780 1687.750 ;
        RECT 1514.420 1655.470 1514.680 1655.790 ;
        RECT 1514.480 16.310 1514.620 1655.470 ;
        RECT 1495.560 15.990 1495.820 16.310 ;
        RECT 1514.420 15.990 1514.680 16.310 ;
        RECT 1495.620 2.400 1495.760 15.990 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1521.290 1686.980 1521.610 1687.040 ;
        RECT 1558.090 1686.980 1558.410 1687.040 ;
        RECT 1521.290 1686.840 1558.410 1686.980 ;
        RECT 1521.290 1686.780 1521.610 1686.840 ;
        RECT 1558.090 1686.780 1558.410 1686.840 ;
        RECT 1513.010 20.640 1513.330 20.700 ;
        RECT 1521.290 20.640 1521.610 20.700 ;
        RECT 1513.010 20.500 1521.610 20.640 ;
        RECT 1513.010 20.440 1513.330 20.500 ;
        RECT 1521.290 20.440 1521.610 20.500 ;
      LAYER via ;
        RECT 1521.320 1686.780 1521.580 1687.040 ;
        RECT 1558.120 1686.780 1558.380 1687.040 ;
        RECT 1513.040 20.440 1513.300 20.700 ;
        RECT 1521.320 20.440 1521.580 20.700 ;
      LAYER met2 ;
        RECT 1558.110 1700.000 1558.390 1704.000 ;
        RECT 1558.180 1687.070 1558.320 1700.000 ;
        RECT 1521.320 1686.750 1521.580 1687.070 ;
        RECT 1558.120 1686.750 1558.380 1687.070 ;
        RECT 1521.380 20.730 1521.520 1686.750 ;
        RECT 1513.040 20.410 1513.300 20.730 ;
        RECT 1521.320 20.410 1521.580 20.730 ;
        RECT 1513.100 2.400 1513.240 20.410 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1338.670 1678.140 1338.990 1678.200 ;
        RECT 1340.510 1678.140 1340.830 1678.200 ;
        RECT 1338.670 1678.000 1340.830 1678.140 ;
        RECT 1338.670 1677.940 1338.990 1678.000 ;
        RECT 1340.510 1677.940 1340.830 1678.000 ;
        RECT 709.850 39.340 710.170 39.400 ;
        RECT 1338.670 39.340 1338.990 39.400 ;
        RECT 709.850 39.200 1338.990 39.340 ;
        RECT 709.850 39.140 710.170 39.200 ;
        RECT 1338.670 39.140 1338.990 39.200 ;
      LAYER via ;
        RECT 1338.700 1677.940 1338.960 1678.200 ;
        RECT 1340.540 1677.940 1340.800 1678.200 ;
        RECT 709.880 39.140 710.140 39.400 ;
        RECT 1338.700 39.140 1338.960 39.400 ;
      LAYER met2 ;
        RECT 1341.450 1700.410 1341.730 1704.000 ;
        RECT 1340.600 1700.270 1341.730 1700.410 ;
        RECT 1340.600 1678.230 1340.740 1700.270 ;
        RECT 1341.450 1700.000 1341.730 1700.270 ;
        RECT 1338.700 1677.910 1338.960 1678.230 ;
        RECT 1340.540 1677.910 1340.800 1678.230 ;
        RECT 1338.760 39.430 1338.900 1677.910 ;
        RECT 709.880 39.110 710.140 39.430 ;
        RECT 1338.700 39.110 1338.960 39.430 ;
        RECT 709.940 17.410 710.080 39.110 ;
        RECT 709.940 17.270 710.540 17.410 ;
        RECT 710.400 2.400 710.540 17.270 ;
        RECT 710.190 -4.800 710.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1531.410 1689.700 1531.730 1689.760 ;
        RECT 1563.150 1689.700 1563.470 1689.760 ;
        RECT 1531.410 1689.560 1563.470 1689.700 ;
        RECT 1531.410 1689.500 1531.730 1689.560 ;
        RECT 1563.150 1689.500 1563.470 1689.560 ;
      LAYER via ;
        RECT 1531.440 1689.500 1531.700 1689.760 ;
        RECT 1563.180 1689.500 1563.440 1689.760 ;
      LAYER met2 ;
        RECT 1563.170 1700.000 1563.450 1704.000 ;
        RECT 1563.240 1689.790 1563.380 1700.000 ;
        RECT 1531.440 1689.470 1531.700 1689.790 ;
        RECT 1563.180 1689.470 1563.440 1689.790 ;
        RECT 1531.500 3.130 1531.640 1689.470 ;
        RECT 1531.040 2.990 1531.640 3.130 ;
        RECT 1531.040 2.400 1531.180 2.990 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1552.110 1689.020 1552.430 1689.080 ;
        RECT 1567.750 1689.020 1568.070 1689.080 ;
        RECT 1552.110 1688.880 1568.070 1689.020 ;
        RECT 1552.110 1688.820 1552.430 1688.880 ;
        RECT 1567.750 1688.820 1568.070 1688.880 ;
        RECT 1548.890 20.640 1549.210 20.700 ;
        RECT 1552.110 20.640 1552.430 20.700 ;
        RECT 1548.890 20.500 1552.430 20.640 ;
        RECT 1548.890 20.440 1549.210 20.500 ;
        RECT 1552.110 20.440 1552.430 20.500 ;
      LAYER via ;
        RECT 1552.140 1688.820 1552.400 1689.080 ;
        RECT 1567.780 1688.820 1568.040 1689.080 ;
        RECT 1548.920 20.440 1549.180 20.700 ;
        RECT 1552.140 20.440 1552.400 20.700 ;
      LAYER met2 ;
        RECT 1567.770 1700.000 1568.050 1704.000 ;
        RECT 1567.840 1689.110 1567.980 1700.000 ;
        RECT 1552.140 1688.790 1552.400 1689.110 ;
        RECT 1567.780 1688.790 1568.040 1689.110 ;
        RECT 1552.200 20.730 1552.340 1688.790 ;
        RECT 1548.920 20.410 1549.180 20.730 ;
        RECT 1552.140 20.410 1552.400 20.730 ;
        RECT 1548.980 2.400 1549.120 20.410 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1567.290 1678.140 1567.610 1678.200 ;
        RECT 1571.890 1678.140 1572.210 1678.200 ;
        RECT 1567.290 1678.000 1572.210 1678.140 ;
        RECT 1567.290 1677.940 1567.610 1678.000 ;
        RECT 1571.890 1677.940 1572.210 1678.000 ;
      LAYER via ;
        RECT 1567.320 1677.940 1567.580 1678.200 ;
        RECT 1571.920 1677.940 1572.180 1678.200 ;
      LAYER met2 ;
        RECT 1572.830 1700.410 1573.110 1704.000 ;
        RECT 1571.980 1700.270 1573.110 1700.410 ;
        RECT 1571.980 1678.230 1572.120 1700.270 ;
        RECT 1572.830 1700.000 1573.110 1700.270 ;
        RECT 1567.320 1677.910 1567.580 1678.230 ;
        RECT 1571.920 1677.910 1572.180 1678.230 ;
        RECT 1567.380 3.130 1567.520 1677.910 ;
        RECT 1566.920 2.990 1567.520 3.130 ;
        RECT 1566.920 2.400 1567.060 2.990 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 0.300 ;
=======
      LAYER met1 ;
        RECT 1577.410 1683.920 1577.730 1683.980 ;
        RECT 1580.630 1683.920 1580.950 1683.980 ;
        RECT 1577.410 1683.780 1580.950 1683.920 ;
        RECT 1577.410 1683.720 1577.730 1683.780 ;
        RECT 1580.630 1683.720 1580.950 1683.780 ;
        RECT 1580.630 2.960 1580.950 3.020 ;
        RECT 1584.770 2.960 1585.090 3.020 ;
        RECT 1580.630 2.820 1585.090 2.960 ;
        RECT 1580.630 2.760 1580.950 2.820 ;
        RECT 1584.770 2.760 1585.090 2.820 ;
      LAYER via ;
        RECT 1577.440 1683.720 1577.700 1683.980 ;
        RECT 1580.660 1683.720 1580.920 1683.980 ;
        RECT 1580.660 2.760 1580.920 3.020 ;
        RECT 1584.800 2.760 1585.060 3.020 ;
      LAYER met2 ;
        RECT 1577.430 1700.000 1577.710 1704.000 ;
        RECT 1577.500 1684.010 1577.640 1700.000 ;
        RECT 1577.440 1683.690 1577.700 1684.010 ;
        RECT 1580.660 1683.690 1580.920 1684.010 ;
        RECT 1580.720 3.050 1580.860 1683.690 ;
        RECT 1580.660 2.730 1580.920 3.050 ;
        RECT 1584.800 2.730 1585.060 3.050 ;
        RECT 1584.860 2.400 1585.000 2.730 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1582.470 1683.920 1582.790 1683.980 ;
        RECT 1586.610 1683.920 1586.930 1683.980 ;
        RECT 1582.470 1683.780 1586.930 1683.920 ;
        RECT 1582.470 1683.720 1582.790 1683.780 ;
        RECT 1586.610 1683.720 1586.930 1683.780 ;
        RECT 1586.610 20.300 1586.930 20.360 ;
        RECT 1602.250 20.300 1602.570 20.360 ;
        RECT 1586.610 20.160 1602.570 20.300 ;
        RECT 1586.610 20.100 1586.930 20.160 ;
        RECT 1602.250 20.100 1602.570 20.160 ;
      LAYER via ;
        RECT 1582.500 1683.720 1582.760 1683.980 ;
        RECT 1586.640 1683.720 1586.900 1683.980 ;
        RECT 1586.640 20.100 1586.900 20.360 ;
        RECT 1602.280 20.100 1602.540 20.360 ;
      LAYER met2 ;
        RECT 1582.490 1700.000 1582.770 1704.000 ;
        RECT 1582.560 1684.010 1582.700 1700.000 ;
        RECT 1582.500 1683.690 1582.760 1684.010 ;
        RECT 1586.640 1683.690 1586.900 1684.010 ;
        RECT 1586.700 20.390 1586.840 1683.690 ;
        RECT 1586.640 20.070 1586.900 20.390 ;
        RECT 1602.280 20.070 1602.540 20.390 ;
        RECT 1602.340 2.400 1602.480 20.070 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 0.300 ;
=======
      LAYER met1 ;
        RECT 1587.070 1684.940 1587.390 1685.000 ;
        RECT 1604.090 1684.940 1604.410 1685.000 ;
        RECT 1587.070 1684.800 1604.410 1684.940 ;
        RECT 1587.070 1684.740 1587.390 1684.800 ;
        RECT 1604.090 1684.740 1604.410 1684.800 ;
        RECT 1604.090 16.560 1604.410 16.620 ;
        RECT 1620.190 16.560 1620.510 16.620 ;
        RECT 1604.090 16.420 1620.510 16.560 ;
        RECT 1604.090 16.360 1604.410 16.420 ;
        RECT 1620.190 16.360 1620.510 16.420 ;
      LAYER via ;
        RECT 1587.100 1684.740 1587.360 1685.000 ;
        RECT 1604.120 1684.740 1604.380 1685.000 ;
        RECT 1604.120 16.360 1604.380 16.620 ;
        RECT 1620.220 16.360 1620.480 16.620 ;
      LAYER met2 ;
        RECT 1587.090 1700.000 1587.370 1704.000 ;
        RECT 1587.160 1685.030 1587.300 1700.000 ;
        RECT 1587.100 1684.710 1587.360 1685.030 ;
        RECT 1604.120 1684.710 1604.380 1685.030 ;
        RECT 1604.180 16.650 1604.320 1684.710 ;
        RECT 1604.120 16.330 1604.380 16.650 ;
        RECT 1620.220 16.330 1620.480 16.650 ;
        RECT 1620.280 2.400 1620.420 16.330 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1592.130 1686.980 1592.450 1687.040 ;
        RECT 1617.890 1686.980 1618.210 1687.040 ;
        RECT 1592.130 1686.840 1618.210 1686.980 ;
        RECT 1592.130 1686.780 1592.450 1686.840 ;
        RECT 1617.890 1686.780 1618.210 1686.840 ;
        RECT 1617.890 15.200 1618.210 15.260 ;
        RECT 1638.130 15.200 1638.450 15.260 ;
        RECT 1617.890 15.060 1638.450 15.200 ;
        RECT 1617.890 15.000 1618.210 15.060 ;
        RECT 1638.130 15.000 1638.450 15.060 ;
      LAYER via ;
        RECT 1592.160 1686.780 1592.420 1687.040 ;
        RECT 1617.920 1686.780 1618.180 1687.040 ;
        RECT 1617.920 15.000 1618.180 15.260 ;
        RECT 1638.160 15.000 1638.420 15.260 ;
      LAYER met2 ;
        RECT 1592.150 1700.000 1592.430 1704.000 ;
        RECT 1592.220 1687.070 1592.360 1700.000 ;
        RECT 1592.160 1686.750 1592.420 1687.070 ;
        RECT 1617.920 1686.750 1618.180 1687.070 ;
        RECT 1617.980 15.290 1618.120 1686.750 ;
        RECT 1617.920 14.970 1618.180 15.290 ;
        RECT 1638.160 14.970 1638.420 15.290 ;
        RECT 1638.220 2.400 1638.360 14.970 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 0.300 ;
=======
      LAYER li1 ;
        RECT 1621.645 16.745 1621.815 18.275 ;
      LAYER mcon ;
        RECT 1621.645 18.105 1621.815 18.275 ;
      LAYER met1 ;
        RECT 1596.730 1683.920 1597.050 1683.980 ;
        RECT 1600.410 1683.920 1600.730 1683.980 ;
        RECT 1596.730 1683.780 1600.730 1683.920 ;
        RECT 1596.730 1683.720 1597.050 1683.780 ;
        RECT 1600.410 1683.720 1600.730 1683.780 ;
        RECT 1600.410 18.260 1600.730 18.320 ;
        RECT 1621.585 18.260 1621.875 18.305 ;
        RECT 1600.410 18.120 1621.875 18.260 ;
        RECT 1600.410 18.060 1600.730 18.120 ;
        RECT 1621.585 18.075 1621.875 18.120 ;
        RECT 1621.585 16.900 1621.875 16.945 ;
        RECT 1656.070 16.900 1656.390 16.960 ;
        RECT 1621.585 16.760 1656.390 16.900 ;
        RECT 1621.585 16.715 1621.875 16.760 ;
        RECT 1656.070 16.700 1656.390 16.760 ;
      LAYER via ;
        RECT 1596.760 1683.720 1597.020 1683.980 ;
        RECT 1600.440 1683.720 1600.700 1683.980 ;
        RECT 1600.440 18.060 1600.700 18.320 ;
        RECT 1656.100 16.700 1656.360 16.960 ;
      LAYER met2 ;
        RECT 1596.750 1700.000 1597.030 1704.000 ;
        RECT 1596.820 1684.010 1596.960 1700.000 ;
        RECT 1596.760 1683.690 1597.020 1684.010 ;
        RECT 1600.440 1683.690 1600.700 1684.010 ;
        RECT 1600.500 18.350 1600.640 1683.690 ;
        RECT 1600.440 18.030 1600.700 18.350 ;
        RECT 1656.100 16.670 1656.360 16.990 ;
        RECT 1656.160 2.400 1656.300 16.670 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 0.300 ;
=======
      LAYER li1 ;
        RECT 1628.545 1686.485 1628.715 1688.015 ;
      LAYER mcon ;
        RECT 1628.545 1687.845 1628.715 1688.015 ;
      LAYER met1 ;
        RECT 1601.790 1688.000 1602.110 1688.060 ;
        RECT 1628.485 1688.000 1628.775 1688.045 ;
        RECT 1601.790 1687.860 1628.775 1688.000 ;
        RECT 1601.790 1687.800 1602.110 1687.860 ;
        RECT 1628.485 1687.815 1628.775 1687.860 ;
        RECT 1628.485 1686.640 1628.775 1686.685 ;
        RECT 1666.190 1686.640 1666.510 1686.700 ;
        RECT 1628.485 1686.500 1666.510 1686.640 ;
        RECT 1628.485 1686.455 1628.775 1686.500 ;
        RECT 1666.190 1686.440 1666.510 1686.500 ;
        RECT 1666.190 17.580 1666.510 17.640 ;
        RECT 1673.550 17.580 1673.870 17.640 ;
        RECT 1666.190 17.440 1673.870 17.580 ;
        RECT 1666.190 17.380 1666.510 17.440 ;
        RECT 1673.550 17.380 1673.870 17.440 ;
      LAYER via ;
        RECT 1601.820 1687.800 1602.080 1688.060 ;
        RECT 1666.220 1686.440 1666.480 1686.700 ;
        RECT 1666.220 17.380 1666.480 17.640 ;
        RECT 1673.580 17.380 1673.840 17.640 ;
      LAYER met2 ;
        RECT 1601.810 1700.000 1602.090 1704.000 ;
        RECT 1601.880 1688.090 1602.020 1700.000 ;
        RECT 1601.820 1687.770 1602.080 1688.090 ;
        RECT 1666.220 1686.410 1666.480 1686.730 ;
        RECT 1666.280 17.670 1666.420 1686.410 ;
        RECT 1666.220 17.350 1666.480 17.670 ;
        RECT 1673.580 17.350 1673.840 17.670 ;
        RECT 1673.640 2.400 1673.780 17.350 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1607.310 19.620 1607.630 19.680 ;
        RECT 1691.490 19.620 1691.810 19.680 ;
        RECT 1607.310 19.480 1691.810 19.620 ;
        RECT 1607.310 19.420 1607.630 19.480 ;
        RECT 1691.490 19.420 1691.810 19.480 ;
      LAYER via ;
        RECT 1607.340 19.420 1607.600 19.680 ;
        RECT 1691.520 19.420 1691.780 19.680 ;
      LAYER met2 ;
        RECT 1606.410 1700.410 1606.690 1704.000 ;
        RECT 1606.410 1700.270 1607.540 1700.410 ;
        RECT 1606.410 1700.000 1606.690 1700.270 ;
        RECT 1607.400 19.710 1607.540 1700.270 ;
        RECT 1607.340 19.390 1607.600 19.710 ;
        RECT 1691.520 19.390 1691.780 19.710 ;
        RECT 1691.580 2.400 1691.720 19.390 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 0.300 ;
=======
      LAYER met1 ;
        RECT 728.250 39.680 728.570 39.740 ;
        RECT 1346.490 39.680 1346.810 39.740 ;
        RECT 728.250 39.540 1346.810 39.680 ;
        RECT 728.250 39.480 728.570 39.540 ;
        RECT 1346.490 39.480 1346.810 39.540 ;
      LAYER via ;
        RECT 728.280 39.480 728.540 39.740 ;
        RECT 1346.520 39.480 1346.780 39.740 ;
      LAYER met2 ;
        RECT 1346.510 1700.000 1346.790 1704.000 ;
        RECT 1346.580 39.770 1346.720 1700.000 ;
        RECT 728.280 39.450 728.540 39.770 ;
        RECT 1346.520 39.450 1346.780 39.770 ;
        RECT 728.340 2.400 728.480 39.450 ;
        RECT 728.130 -4.800 728.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 0.300 ;
=======
      LAYER met1 ;
        RECT 1611.450 1688.680 1611.770 1688.740 ;
        RECT 1614.210 1688.680 1614.530 1688.740 ;
        RECT 1611.450 1688.540 1614.530 1688.680 ;
        RECT 1611.450 1688.480 1611.770 1688.540 ;
        RECT 1614.210 1688.480 1614.530 1688.540 ;
        RECT 1614.210 18.600 1614.530 18.660 ;
        RECT 1709.430 18.600 1709.750 18.660 ;
        RECT 1614.210 18.460 1709.750 18.600 ;
        RECT 1614.210 18.400 1614.530 18.460 ;
        RECT 1709.430 18.400 1709.750 18.460 ;
      LAYER via ;
        RECT 1611.480 1688.480 1611.740 1688.740 ;
        RECT 1614.240 1688.480 1614.500 1688.740 ;
        RECT 1614.240 18.400 1614.500 18.660 ;
        RECT 1709.460 18.400 1709.720 18.660 ;
      LAYER met2 ;
        RECT 1611.470 1700.000 1611.750 1704.000 ;
        RECT 1611.540 1688.770 1611.680 1700.000 ;
        RECT 1611.480 1688.450 1611.740 1688.770 ;
        RECT 1614.240 1688.450 1614.500 1688.770 ;
        RECT 1614.300 18.690 1614.440 1688.450 ;
        RECT 1614.240 18.370 1614.500 18.690 ;
        RECT 1709.460 18.370 1709.720 18.690 ;
        RECT 1709.520 2.400 1709.660 18.370 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1616.050 1685.280 1616.370 1685.340 ;
        RECT 1621.110 1685.280 1621.430 1685.340 ;
        RECT 1616.050 1685.140 1621.430 1685.280 ;
        RECT 1616.050 1685.080 1616.370 1685.140 ;
        RECT 1621.110 1685.080 1621.430 1685.140 ;
        RECT 1621.110 17.920 1621.430 17.980 ;
        RECT 1727.370 17.920 1727.690 17.980 ;
        RECT 1621.110 17.780 1727.690 17.920 ;
        RECT 1621.110 17.720 1621.430 17.780 ;
        RECT 1727.370 17.720 1727.690 17.780 ;
      LAYER via ;
        RECT 1616.080 1685.080 1616.340 1685.340 ;
        RECT 1621.140 1685.080 1621.400 1685.340 ;
        RECT 1621.140 17.720 1621.400 17.980 ;
        RECT 1727.400 17.720 1727.660 17.980 ;
      LAYER met2 ;
        RECT 1616.070 1700.000 1616.350 1704.000 ;
        RECT 1616.140 1685.370 1616.280 1700.000 ;
        RECT 1616.080 1685.050 1616.340 1685.370 ;
        RECT 1621.140 1685.050 1621.400 1685.370 ;
        RECT 1621.200 18.010 1621.340 1685.050 ;
        RECT 1621.140 17.690 1621.400 18.010 ;
        RECT 1727.400 17.690 1727.660 18.010 ;
        RECT 1727.460 2.400 1727.600 17.690 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 0.300 ;
=======
      LAYER li1 ;
        RECT 1638.665 15.045 1638.835 16.235 ;
        RECT 1653.385 15.215 1653.555 16.575 ;
        RECT 1652.005 15.045 1653.555 15.215 ;
        RECT 1675.465 14.365 1675.635 16.575 ;
        RECT 1732.965 14.365 1734.515 14.535 ;
      LAYER mcon ;
        RECT 1653.385 16.405 1653.555 16.575 ;
        RECT 1638.665 16.065 1638.835 16.235 ;
        RECT 1675.465 16.405 1675.635 16.575 ;
        RECT 1734.345 14.365 1734.515 14.535 ;
      LAYER met1 ;
        RECT 1621.570 1684.940 1621.890 1685.000 ;
        RECT 1631.690 1684.940 1632.010 1685.000 ;
        RECT 1621.570 1684.800 1632.010 1684.940 ;
        RECT 1621.570 1684.740 1621.890 1684.800 ;
        RECT 1631.690 1684.740 1632.010 1684.800 ;
        RECT 1631.690 19.960 1632.010 20.020 ;
        RECT 1633.070 19.960 1633.390 20.020 ;
        RECT 1631.690 19.820 1633.390 19.960 ;
        RECT 1631.690 19.760 1632.010 19.820 ;
        RECT 1633.070 19.760 1633.390 19.820 ;
        RECT 1653.325 16.560 1653.615 16.605 ;
        RECT 1675.405 16.560 1675.695 16.605 ;
        RECT 1653.325 16.420 1675.695 16.560 ;
        RECT 1653.325 16.375 1653.615 16.420 ;
        RECT 1675.405 16.375 1675.695 16.420 ;
        RECT 1633.070 16.220 1633.390 16.280 ;
        RECT 1638.605 16.220 1638.895 16.265 ;
        RECT 1633.070 16.080 1638.895 16.220 ;
        RECT 1633.070 16.020 1633.390 16.080 ;
        RECT 1638.605 16.035 1638.895 16.080 ;
        RECT 1638.605 15.200 1638.895 15.245 ;
        RECT 1651.945 15.200 1652.235 15.245 ;
        RECT 1638.605 15.060 1652.235 15.200 ;
        RECT 1638.605 15.015 1638.895 15.060 ;
        RECT 1651.945 15.015 1652.235 15.060 ;
        RECT 1675.405 14.520 1675.695 14.565 ;
        RECT 1732.905 14.520 1733.195 14.565 ;
        RECT 1675.405 14.380 1733.195 14.520 ;
        RECT 1675.405 14.335 1675.695 14.380 ;
        RECT 1732.905 14.335 1733.195 14.380 ;
        RECT 1734.285 14.520 1734.575 14.565 ;
        RECT 1745.310 14.520 1745.630 14.580 ;
        RECT 1734.285 14.380 1745.630 14.520 ;
        RECT 1734.285 14.335 1734.575 14.380 ;
        RECT 1745.310 14.320 1745.630 14.380 ;
      LAYER via ;
        RECT 1621.600 1684.740 1621.860 1685.000 ;
        RECT 1631.720 1684.740 1631.980 1685.000 ;
        RECT 1631.720 19.760 1631.980 20.020 ;
        RECT 1633.100 19.760 1633.360 20.020 ;
        RECT 1633.100 16.020 1633.360 16.280 ;
        RECT 1745.340 14.320 1745.600 14.580 ;
      LAYER met2 ;
        RECT 1621.130 1700.000 1621.410 1704.000 ;
        RECT 1621.200 1686.130 1621.340 1700.000 ;
        RECT 1621.200 1685.990 1621.800 1686.130 ;
        RECT 1621.660 1685.030 1621.800 1685.990 ;
        RECT 1621.600 1684.710 1621.860 1685.030 ;
        RECT 1631.720 1684.710 1631.980 1685.030 ;
        RECT 1631.780 20.050 1631.920 1684.710 ;
        RECT 1631.720 19.730 1631.980 20.050 ;
        RECT 1633.100 19.730 1633.360 20.050 ;
        RECT 1633.160 16.310 1633.300 19.730 ;
        RECT 1633.100 15.990 1633.360 16.310 ;
        RECT 1745.340 14.290 1745.600 14.610 ;
        RECT 1745.400 2.400 1745.540 14.290 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 0.300 ;
=======
      LAYER met1 ;
        RECT 1625.710 1688.680 1626.030 1688.740 ;
        RECT 1628.010 1688.680 1628.330 1688.740 ;
        RECT 1625.710 1688.540 1628.330 1688.680 ;
        RECT 1625.710 1688.480 1626.030 1688.540 ;
        RECT 1628.010 1688.480 1628.330 1688.540 ;
        RECT 1628.010 15.540 1628.330 15.600 ;
        RECT 1628.010 15.400 1652.620 15.540 ;
        RECT 1628.010 15.340 1628.330 15.400 ;
        RECT 1652.480 15.200 1652.620 15.400 ;
        RECT 1762.790 15.200 1763.110 15.260 ;
        RECT 1652.480 15.060 1763.110 15.200 ;
        RECT 1762.790 15.000 1763.110 15.060 ;
      LAYER via ;
        RECT 1625.740 1688.480 1626.000 1688.740 ;
        RECT 1628.040 1688.480 1628.300 1688.740 ;
        RECT 1628.040 15.340 1628.300 15.600 ;
        RECT 1762.820 15.000 1763.080 15.260 ;
      LAYER met2 ;
        RECT 1625.730 1700.000 1626.010 1704.000 ;
        RECT 1625.800 1688.770 1625.940 1700.000 ;
        RECT 1625.740 1688.450 1626.000 1688.770 ;
        RECT 1628.040 1688.450 1628.300 1688.770 ;
        RECT 1628.100 15.630 1628.240 1688.450 ;
        RECT 1628.040 15.310 1628.300 15.630 ;
        RECT 1762.820 14.970 1763.080 15.290 ;
        RECT 1762.880 2.400 1763.020 14.970 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 0.300 ;
=======
      LAYER li1 ;
        RECT 1644.645 17.425 1644.815 19.975 ;
        RECT 1656.605 16.745 1656.775 17.595 ;
      LAYER mcon ;
        RECT 1644.645 19.805 1644.815 19.975 ;
        RECT 1656.605 17.425 1656.775 17.595 ;
      LAYER met1 ;
        RECT 1630.770 1688.340 1631.090 1688.400 ;
        RECT 1634.910 1688.340 1635.230 1688.400 ;
        RECT 1630.770 1688.200 1635.230 1688.340 ;
        RECT 1630.770 1688.140 1631.090 1688.200 ;
        RECT 1634.910 1688.140 1635.230 1688.200 ;
        RECT 1634.910 19.960 1635.230 20.020 ;
        RECT 1644.585 19.960 1644.875 20.005 ;
        RECT 1634.910 19.820 1644.875 19.960 ;
        RECT 1634.910 19.760 1635.230 19.820 ;
        RECT 1644.585 19.775 1644.875 19.820 ;
        RECT 1644.585 17.580 1644.875 17.625 ;
        RECT 1656.545 17.580 1656.835 17.625 ;
        RECT 1644.585 17.440 1656.835 17.580 ;
        RECT 1644.585 17.395 1644.875 17.440 ;
        RECT 1656.545 17.395 1656.835 17.440 ;
        RECT 1656.545 16.900 1656.835 16.945 ;
        RECT 1780.730 16.900 1781.050 16.960 ;
        RECT 1656.545 16.760 1781.050 16.900 ;
        RECT 1656.545 16.715 1656.835 16.760 ;
        RECT 1780.730 16.700 1781.050 16.760 ;
      LAYER via ;
        RECT 1630.800 1688.140 1631.060 1688.400 ;
        RECT 1634.940 1688.140 1635.200 1688.400 ;
        RECT 1634.940 19.760 1635.200 20.020 ;
        RECT 1780.760 16.700 1781.020 16.960 ;
      LAYER met2 ;
        RECT 1630.790 1700.000 1631.070 1704.000 ;
        RECT 1630.860 1688.430 1631.000 1700.000 ;
        RECT 1630.800 1688.110 1631.060 1688.430 ;
        RECT 1634.940 1688.110 1635.200 1688.430 ;
        RECT 1635.000 20.050 1635.140 1688.110 ;
        RECT 1634.940 19.730 1635.200 20.050 ;
        RECT 1780.760 16.670 1781.020 16.990 ;
        RECT 1780.820 2.400 1780.960 16.670 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1635.370 1689.020 1635.690 1689.080 ;
        RECT 1640.890 1689.020 1641.210 1689.080 ;
        RECT 1635.370 1688.880 1641.210 1689.020 ;
        RECT 1635.370 1688.820 1635.690 1688.880 ;
        RECT 1640.890 1688.820 1641.210 1688.880 ;
        RECT 1640.890 22.000 1641.210 22.060 ;
        RECT 1798.670 22.000 1798.990 22.060 ;
        RECT 1640.890 21.860 1798.990 22.000 ;
        RECT 1640.890 21.800 1641.210 21.860 ;
        RECT 1798.670 21.800 1798.990 21.860 ;
      LAYER via ;
        RECT 1635.400 1688.820 1635.660 1689.080 ;
        RECT 1640.920 1688.820 1641.180 1689.080 ;
        RECT 1640.920 21.800 1641.180 22.060 ;
        RECT 1798.700 21.800 1798.960 22.060 ;
      LAYER met2 ;
        RECT 1635.390 1700.000 1635.670 1704.000 ;
        RECT 1635.460 1689.110 1635.600 1700.000 ;
        RECT 1635.400 1688.790 1635.660 1689.110 ;
        RECT 1640.920 1688.790 1641.180 1689.110 ;
        RECT 1640.980 22.090 1641.120 1688.790 ;
        RECT 1640.920 21.770 1641.180 22.090 ;
        RECT 1798.700 21.770 1798.960 22.090 ;
        RECT 1798.760 2.400 1798.900 21.770 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1816.610 23.360 1816.930 23.420 ;
        RECT 1801.980 23.220 1816.930 23.360 ;
        RECT 1639.970 23.020 1640.290 23.080 ;
        RECT 1801.980 23.020 1802.120 23.220 ;
        RECT 1816.610 23.160 1816.930 23.220 ;
        RECT 1639.970 22.880 1802.120 23.020 ;
        RECT 1639.970 22.820 1640.290 22.880 ;
      LAYER via ;
        RECT 1640.000 22.820 1640.260 23.080 ;
        RECT 1816.640 23.160 1816.900 23.420 ;
      LAYER met2 ;
        RECT 1640.450 1700.410 1640.730 1704.000 ;
        RECT 1640.060 1700.270 1640.730 1700.410 ;
        RECT 1640.060 23.110 1640.200 1700.270 ;
        RECT 1640.450 1700.000 1640.730 1700.270 ;
        RECT 1816.640 23.130 1816.900 23.450 ;
        RECT 1640.000 22.790 1640.260 23.110 ;
        RECT 1816.700 2.400 1816.840 23.130 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 0.300 ;
=======
      LAYER li1 ;
        RECT 1801.505 22.185 1801.675 23.375 ;
      LAYER mcon ;
        RECT 1801.505 23.205 1801.675 23.375 ;
      LAYER met1 ;
        RECT 1645.030 1688.340 1645.350 1688.400 ;
        RECT 1648.250 1688.340 1648.570 1688.400 ;
        RECT 1645.030 1688.200 1648.570 1688.340 ;
        RECT 1645.030 1688.140 1645.350 1688.200 ;
        RECT 1648.250 1688.140 1648.570 1688.200 ;
        RECT 1648.250 23.360 1648.570 23.420 ;
        RECT 1801.445 23.360 1801.735 23.405 ;
        RECT 1648.250 23.220 1801.735 23.360 ;
        RECT 1648.250 23.160 1648.570 23.220 ;
        RECT 1801.445 23.175 1801.735 23.220 ;
        RECT 1801.445 22.340 1801.735 22.385 ;
        RECT 1834.550 22.340 1834.870 22.400 ;
        RECT 1801.445 22.200 1834.870 22.340 ;
        RECT 1801.445 22.155 1801.735 22.200 ;
        RECT 1834.550 22.140 1834.870 22.200 ;
      LAYER via ;
        RECT 1645.060 1688.140 1645.320 1688.400 ;
        RECT 1648.280 1688.140 1648.540 1688.400 ;
        RECT 1648.280 23.160 1648.540 23.420 ;
        RECT 1834.580 22.140 1834.840 22.400 ;
      LAYER met2 ;
        RECT 1645.050 1700.000 1645.330 1704.000 ;
        RECT 1645.120 1688.430 1645.260 1700.000 ;
        RECT 1645.060 1688.110 1645.320 1688.430 ;
        RECT 1648.280 1688.110 1648.540 1688.430 ;
        RECT 1648.340 23.450 1648.480 1688.110 ;
        RECT 1648.280 23.130 1648.540 23.450 ;
        RECT 1834.580 22.110 1834.840 22.430 ;
        RECT 1834.640 2.400 1834.780 22.110 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 0.300 ;
=======
      LAYER met1 ;
        RECT 1650.090 1688.340 1650.410 1688.400 ;
        RECT 1654.230 1688.340 1654.550 1688.400 ;
        RECT 1650.090 1688.200 1654.550 1688.340 ;
        RECT 1650.090 1688.140 1650.410 1688.200 ;
        RECT 1654.230 1688.140 1654.550 1688.200 ;
        RECT 1654.230 27.100 1654.550 27.160 ;
        RECT 1654.230 26.960 1825.120 27.100 ;
        RECT 1654.230 26.900 1654.550 26.960 ;
        RECT 1824.980 26.760 1825.120 26.960 ;
        RECT 1852.030 26.760 1852.350 26.820 ;
        RECT 1824.980 26.620 1852.350 26.760 ;
        RECT 1852.030 26.560 1852.350 26.620 ;
      LAYER via ;
        RECT 1650.120 1688.140 1650.380 1688.400 ;
        RECT 1654.260 1688.140 1654.520 1688.400 ;
        RECT 1654.260 26.900 1654.520 27.160 ;
        RECT 1852.060 26.560 1852.320 26.820 ;
      LAYER met2 ;
        RECT 1650.110 1700.000 1650.390 1704.000 ;
        RECT 1650.180 1688.430 1650.320 1700.000 ;
        RECT 1650.120 1688.110 1650.380 1688.430 ;
        RECT 1654.260 1688.110 1654.520 1688.430 ;
        RECT 1654.320 27.190 1654.460 1688.110 ;
        RECT 1654.260 26.870 1654.520 27.190 ;
        RECT 1852.060 26.530 1852.320 26.850 ;
        RECT 1852.120 2.400 1852.260 26.530 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1655.150 26.080 1655.470 26.140 ;
        RECT 1869.970 26.080 1870.290 26.140 ;
        RECT 1655.150 25.940 1870.290 26.080 ;
        RECT 1655.150 25.880 1655.470 25.940 ;
        RECT 1869.970 25.880 1870.290 25.940 ;
      LAYER via ;
        RECT 1655.180 25.880 1655.440 26.140 ;
        RECT 1870.000 25.880 1870.260 26.140 ;
      LAYER met2 ;
        RECT 1654.710 1700.410 1654.990 1704.000 ;
        RECT 1654.710 1700.270 1655.380 1700.410 ;
        RECT 1654.710 1700.000 1654.990 1700.270 ;
        RECT 1655.240 26.170 1655.380 1700.270 ;
        RECT 1655.180 25.850 1655.440 26.170 ;
        RECT 1870.000 25.850 1870.260 26.170 ;
        RECT 1870.060 2.400 1870.200 25.850 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 0.300 ;
=======
      LAYER met1 ;
        RECT 1346.030 1666.580 1346.350 1666.640 ;
        RECT 1350.170 1666.580 1350.490 1666.640 ;
        RECT 1346.030 1666.440 1350.490 1666.580 ;
        RECT 1346.030 1666.380 1346.350 1666.440 ;
        RECT 1350.170 1666.380 1350.490 1666.440 ;
        RECT 746.190 40.020 746.510 40.080 ;
        RECT 1346.030 40.020 1346.350 40.080 ;
        RECT 746.190 39.880 1346.350 40.020 ;
        RECT 746.190 39.820 746.510 39.880 ;
        RECT 1346.030 39.820 1346.350 39.880 ;
      LAYER via ;
        RECT 1346.060 1666.380 1346.320 1666.640 ;
        RECT 1350.200 1666.380 1350.460 1666.640 ;
        RECT 746.220 39.820 746.480 40.080 ;
        RECT 1346.060 39.820 1346.320 40.080 ;
      LAYER met2 ;
        RECT 1351.110 1700.410 1351.390 1704.000 ;
        RECT 1350.260 1700.270 1351.390 1700.410 ;
        RECT 1350.260 1666.670 1350.400 1700.270 ;
        RECT 1351.110 1700.000 1351.390 1700.270 ;
        RECT 1346.060 1666.350 1346.320 1666.670 ;
        RECT 1350.200 1666.350 1350.460 1666.670 ;
        RECT 1346.120 40.110 1346.260 1666.350 ;
        RECT 746.220 39.790 746.480 40.110 ;
        RECT 1346.060 39.790 1346.320 40.110 ;
        RECT 746.280 2.400 746.420 39.790 ;
        RECT 746.070 -4.800 746.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1659.290 1688.680 1659.610 1688.740 ;
        RECT 1661.590 1688.680 1661.910 1688.740 ;
        RECT 1659.290 1688.540 1661.910 1688.680 ;
        RECT 1659.290 1688.480 1659.610 1688.540 ;
        RECT 1661.590 1688.480 1661.910 1688.540 ;
        RECT 1887.910 26.080 1888.230 26.140 ;
        RECT 1870.520 25.940 1888.230 26.080 ;
        RECT 1661.590 25.740 1661.910 25.800 ;
        RECT 1870.520 25.740 1870.660 25.940 ;
        RECT 1887.910 25.880 1888.230 25.940 ;
        RECT 1661.590 25.600 1870.660 25.740 ;
        RECT 1661.590 25.540 1661.910 25.600 ;
      LAYER via ;
        RECT 1659.320 1688.480 1659.580 1688.740 ;
        RECT 1661.620 1688.480 1661.880 1688.740 ;
        RECT 1661.620 25.540 1661.880 25.800 ;
        RECT 1887.940 25.880 1888.200 26.140 ;
      LAYER met2 ;
        RECT 1659.310 1700.000 1659.590 1704.000 ;
        RECT 1659.380 1688.770 1659.520 1700.000 ;
        RECT 1659.320 1688.450 1659.580 1688.770 ;
        RECT 1661.620 1688.450 1661.880 1688.770 ;
        RECT 1661.680 25.830 1661.820 1688.450 ;
        RECT 1887.940 25.850 1888.200 26.170 ;
        RECT 1661.620 25.510 1661.880 25.830 ;
        RECT 1888.000 2.400 1888.140 25.850 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1664.350 1688.680 1664.670 1688.740 ;
        RECT 1668.490 1688.680 1668.810 1688.740 ;
        RECT 1664.350 1688.540 1668.810 1688.680 ;
        RECT 1664.350 1688.480 1664.670 1688.540 ;
        RECT 1668.490 1688.480 1668.810 1688.540 ;
        RECT 1905.850 25.740 1906.170 25.800 ;
        RECT 1872.820 25.600 1906.170 25.740 ;
        RECT 1668.490 25.060 1668.810 25.120 ;
        RECT 1872.820 25.060 1872.960 25.600 ;
        RECT 1905.850 25.540 1906.170 25.600 ;
        RECT 1668.490 24.920 1872.960 25.060 ;
        RECT 1668.490 24.860 1668.810 24.920 ;
      LAYER via ;
        RECT 1664.380 1688.480 1664.640 1688.740 ;
        RECT 1668.520 1688.480 1668.780 1688.740 ;
        RECT 1668.520 24.860 1668.780 25.120 ;
        RECT 1905.880 25.540 1906.140 25.800 ;
      LAYER met2 ;
        RECT 1664.370 1700.000 1664.650 1704.000 ;
        RECT 1664.440 1688.770 1664.580 1700.000 ;
        RECT 1664.380 1688.450 1664.640 1688.770 ;
        RECT 1668.520 1688.450 1668.780 1688.770 ;
        RECT 1668.580 25.150 1668.720 1688.450 ;
        RECT 1905.880 25.510 1906.140 25.830 ;
        RECT 1668.520 24.830 1668.780 25.150 ;
        RECT 1905.940 2.400 1906.080 25.510 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1668.030 24.380 1668.350 24.440 ;
        RECT 1668.030 24.240 1918.960 24.380 ;
        RECT 1668.030 24.180 1668.350 24.240 ;
        RECT 1918.820 24.040 1918.960 24.240 ;
        RECT 1923.330 24.040 1923.650 24.100 ;
        RECT 1918.820 23.900 1923.650 24.040 ;
        RECT 1923.330 23.840 1923.650 23.900 ;
      LAYER via ;
        RECT 1668.060 24.180 1668.320 24.440 ;
        RECT 1923.360 23.840 1923.620 24.100 ;
      LAYER met2 ;
        RECT 1668.970 1700.410 1669.250 1704.000 ;
        RECT 1668.120 1700.270 1669.250 1700.410 ;
        RECT 1668.120 24.470 1668.260 1700.270 ;
        RECT 1668.970 1700.000 1669.250 1700.270 ;
        RECT 1668.060 24.150 1668.320 24.470 ;
        RECT 1923.360 23.810 1923.620 24.130 ;
        RECT 1923.420 2.400 1923.560 23.810 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 0.300 ;
=======
      LAYER met1 ;
        RECT 1674.930 34.920 1675.250 34.980 ;
        RECT 1941.270 34.920 1941.590 34.980 ;
        RECT 1674.930 34.780 1941.590 34.920 ;
        RECT 1674.930 34.720 1675.250 34.780 ;
        RECT 1941.270 34.720 1941.590 34.780 ;
      LAYER via ;
        RECT 1674.960 34.720 1675.220 34.980 ;
        RECT 1941.300 34.720 1941.560 34.980 ;
      LAYER met2 ;
        RECT 1674.030 1700.410 1674.310 1704.000 ;
        RECT 1674.030 1700.270 1675.160 1700.410 ;
        RECT 1674.030 1700.000 1674.310 1700.270 ;
        RECT 1675.020 35.010 1675.160 1700.270 ;
        RECT 1674.960 34.690 1675.220 35.010 ;
        RECT 1941.300 34.690 1941.560 35.010 ;
        RECT 1941.360 2.400 1941.500 34.690 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1678.610 1688.680 1678.930 1688.740 ;
        RECT 1682.290 1688.680 1682.610 1688.740 ;
        RECT 1678.610 1688.540 1682.610 1688.680 ;
        RECT 1678.610 1688.480 1678.930 1688.540 ;
        RECT 1682.290 1688.480 1682.610 1688.540 ;
        RECT 1682.290 35.260 1682.610 35.320 ;
        RECT 1959.210 35.260 1959.530 35.320 ;
        RECT 1682.290 35.120 1959.530 35.260 ;
        RECT 1682.290 35.060 1682.610 35.120 ;
        RECT 1959.210 35.060 1959.530 35.120 ;
      LAYER via ;
        RECT 1678.640 1688.480 1678.900 1688.740 ;
        RECT 1682.320 1688.480 1682.580 1688.740 ;
        RECT 1682.320 35.060 1682.580 35.320 ;
        RECT 1959.240 35.060 1959.500 35.320 ;
      LAYER met2 ;
        RECT 1678.630 1700.000 1678.910 1704.000 ;
        RECT 1678.700 1688.770 1678.840 1700.000 ;
        RECT 1678.640 1688.450 1678.900 1688.770 ;
        RECT 1682.320 1688.450 1682.580 1688.770 ;
        RECT 1682.380 35.350 1682.520 1688.450 ;
        RECT 1682.320 35.030 1682.580 35.350 ;
        RECT 1959.240 35.030 1959.500 35.350 ;
        RECT 1959.300 2.400 1959.440 35.030 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1683.670 1684.940 1683.990 1685.000 ;
        RECT 1688.730 1684.940 1689.050 1685.000 ;
        RECT 1683.670 1684.800 1689.050 1684.940 ;
        RECT 1683.670 1684.740 1683.990 1684.800 ;
        RECT 1688.730 1684.740 1689.050 1684.800 ;
        RECT 1688.730 35.600 1689.050 35.660 ;
        RECT 1977.150 35.600 1977.470 35.660 ;
        RECT 1688.730 35.460 1977.470 35.600 ;
        RECT 1688.730 35.400 1689.050 35.460 ;
        RECT 1977.150 35.400 1977.470 35.460 ;
      LAYER via ;
        RECT 1683.700 1684.740 1683.960 1685.000 ;
        RECT 1688.760 1684.740 1689.020 1685.000 ;
        RECT 1688.760 35.400 1689.020 35.660 ;
        RECT 1977.180 35.400 1977.440 35.660 ;
      LAYER met2 ;
        RECT 1683.690 1700.000 1683.970 1704.000 ;
        RECT 1683.760 1685.030 1683.900 1700.000 ;
        RECT 1683.700 1684.710 1683.960 1685.030 ;
        RECT 1688.760 1684.710 1689.020 1685.030 ;
        RECT 1688.820 35.690 1688.960 1684.710 ;
        RECT 1688.760 35.370 1689.020 35.690 ;
        RECT 1977.180 35.370 1977.440 35.690 ;
        RECT 1977.240 2.400 1977.380 35.370 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1689.190 35.940 1689.510 36.000 ;
        RECT 1995.090 35.940 1995.410 36.000 ;
        RECT 1689.190 35.800 1995.410 35.940 ;
        RECT 1689.190 35.740 1689.510 35.800 ;
        RECT 1995.090 35.740 1995.410 35.800 ;
      LAYER via ;
        RECT 1689.220 35.740 1689.480 36.000 ;
        RECT 1995.120 35.740 1995.380 36.000 ;
      LAYER met2 ;
        RECT 1688.290 1700.410 1688.570 1704.000 ;
        RECT 1688.290 1700.270 1689.420 1700.410 ;
        RECT 1688.290 1700.000 1688.570 1700.270 ;
        RECT 1689.280 36.030 1689.420 1700.270 ;
        RECT 1689.220 35.710 1689.480 36.030 ;
        RECT 1995.120 35.710 1995.380 36.030 ;
        RECT 1995.180 2.400 1995.320 35.710 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1693.330 1688.340 1693.650 1688.400 ;
        RECT 1696.550 1688.340 1696.870 1688.400 ;
        RECT 1693.330 1688.200 1696.870 1688.340 ;
        RECT 1693.330 1688.140 1693.650 1688.200 ;
        RECT 1696.550 1688.140 1696.870 1688.200 ;
        RECT 1696.550 36.280 1696.870 36.340 ;
        RECT 2012.570 36.280 2012.890 36.340 ;
        RECT 1696.550 36.140 2012.890 36.280 ;
        RECT 1696.550 36.080 1696.870 36.140 ;
        RECT 2012.570 36.080 2012.890 36.140 ;
      LAYER via ;
        RECT 1693.360 1688.140 1693.620 1688.400 ;
        RECT 1696.580 1688.140 1696.840 1688.400 ;
        RECT 1696.580 36.080 1696.840 36.340 ;
        RECT 2012.600 36.080 2012.860 36.340 ;
      LAYER met2 ;
        RECT 1693.350 1700.000 1693.630 1704.000 ;
        RECT 1693.420 1688.430 1693.560 1700.000 ;
        RECT 1693.360 1688.110 1693.620 1688.430 ;
        RECT 1696.580 1688.110 1696.840 1688.430 ;
        RECT 1696.640 36.370 1696.780 1688.110 ;
        RECT 1696.580 36.050 1696.840 36.370 ;
        RECT 2012.600 36.050 2012.860 36.370 ;
        RECT 2012.660 2.400 2012.800 36.050 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 0.300 ;
=======
      LAYER met1 ;
        RECT 1697.930 1688.340 1698.250 1688.400 ;
        RECT 1702.990 1688.340 1703.310 1688.400 ;
        RECT 1697.930 1688.200 1703.310 1688.340 ;
        RECT 1697.930 1688.140 1698.250 1688.200 ;
        RECT 1702.990 1688.140 1703.310 1688.200 ;
        RECT 1702.990 42.740 1703.310 42.800 ;
        RECT 2030.510 42.740 2030.830 42.800 ;
        RECT 1702.990 42.600 2030.830 42.740 ;
        RECT 1702.990 42.540 1703.310 42.600 ;
        RECT 2030.510 42.540 2030.830 42.600 ;
      LAYER via ;
        RECT 1697.960 1688.140 1698.220 1688.400 ;
        RECT 1703.020 1688.140 1703.280 1688.400 ;
        RECT 1703.020 42.540 1703.280 42.800 ;
        RECT 2030.540 42.540 2030.800 42.800 ;
      LAYER met2 ;
        RECT 1697.950 1700.000 1698.230 1704.000 ;
        RECT 1698.020 1688.430 1698.160 1700.000 ;
        RECT 1697.960 1688.110 1698.220 1688.430 ;
        RECT 1703.020 1688.110 1703.280 1688.430 ;
        RECT 1703.080 42.830 1703.220 1688.110 ;
        RECT 1703.020 42.510 1703.280 42.830 ;
        RECT 2030.540 42.510 2030.800 42.830 ;
        RECT 2030.600 2.400 2030.740 42.510 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 0.300 ;
=======
      LAYER met1 ;
        RECT 1702.530 43.420 1702.850 43.480 ;
        RECT 2048.450 43.420 2048.770 43.480 ;
        RECT 1702.530 43.280 2048.770 43.420 ;
        RECT 1702.530 43.220 1702.850 43.280 ;
        RECT 2048.450 43.220 2048.770 43.280 ;
      LAYER via ;
        RECT 1702.560 43.220 1702.820 43.480 ;
        RECT 2048.480 43.220 2048.740 43.480 ;
      LAYER met2 ;
        RECT 1703.010 1700.410 1703.290 1704.000 ;
        RECT 1702.620 1700.270 1703.290 1700.410 ;
        RECT 1702.620 43.510 1702.760 1700.270 ;
        RECT 1703.010 1700.000 1703.290 1700.270 ;
        RECT 1702.560 43.190 1702.820 43.510 ;
        RECT 2048.480 43.190 2048.740 43.510 ;
        RECT 2048.540 2.400 2048.680 43.190 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 0.300 ;
=======
      LAYER met1 ;
        RECT 763.670 40.360 763.990 40.420 ;
        RECT 1353.390 40.360 1353.710 40.420 ;
        RECT 763.670 40.220 1353.710 40.360 ;
        RECT 763.670 40.160 763.990 40.220 ;
        RECT 1353.390 40.160 1353.710 40.220 ;
      LAYER via ;
        RECT 763.700 40.160 763.960 40.420 ;
        RECT 1353.420 40.160 1353.680 40.420 ;
      LAYER met2 ;
        RECT 1355.710 1700.410 1355.990 1704.000 ;
        RECT 1354.860 1700.270 1355.990 1700.410 ;
        RECT 1354.860 1677.970 1355.000 1700.270 ;
        RECT 1355.710 1700.000 1355.990 1700.270 ;
        RECT 1353.480 1677.830 1355.000 1677.970 ;
        RECT 1353.480 40.450 1353.620 1677.830 ;
        RECT 763.700 40.130 763.960 40.450 ;
        RECT 1353.420 40.130 1353.680 40.450 ;
        RECT 763.760 2.400 763.900 40.130 ;
        RECT 763.550 -4.800 764.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 0.300 ;
=======
      LAYER met1 ;
        RECT 1708.970 43.760 1709.290 43.820 ;
        RECT 2065.930 43.760 2066.250 43.820 ;
        RECT 1708.970 43.620 2066.250 43.760 ;
        RECT 1708.970 43.560 1709.290 43.620 ;
        RECT 2065.930 43.560 2066.250 43.620 ;
      LAYER via ;
        RECT 1709.000 43.560 1709.260 43.820 ;
        RECT 2065.960 43.560 2066.220 43.820 ;
      LAYER met2 ;
        RECT 1707.610 1700.410 1707.890 1704.000 ;
        RECT 1707.610 1700.270 1709.200 1700.410 ;
        RECT 1707.610 1700.000 1707.890 1700.270 ;
        RECT 1709.060 43.850 1709.200 1700.270 ;
        RECT 1709.000 43.530 1709.260 43.850 ;
        RECT 2065.960 43.530 2066.220 43.850 ;
        RECT 2066.020 17.410 2066.160 43.530 ;
        RECT 2066.020 17.270 2066.620 17.410 ;
        RECT 2066.480 2.400 2066.620 17.270 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1712.650 1688.680 1712.970 1688.740 ;
        RECT 1716.790 1688.680 1717.110 1688.740 ;
        RECT 1712.650 1688.540 1717.110 1688.680 ;
        RECT 1712.650 1688.480 1712.970 1688.540 ;
        RECT 1716.790 1688.480 1717.110 1688.540 ;
        RECT 1716.790 44.100 1717.110 44.160 ;
        RECT 2084.330 44.100 2084.650 44.160 ;
        RECT 1716.790 43.960 2084.650 44.100 ;
        RECT 1716.790 43.900 1717.110 43.960 ;
        RECT 2084.330 43.900 2084.650 43.960 ;
      LAYER via ;
        RECT 1712.680 1688.480 1712.940 1688.740 ;
        RECT 1716.820 1688.480 1717.080 1688.740 ;
        RECT 1716.820 43.900 1717.080 44.160 ;
        RECT 2084.360 43.900 2084.620 44.160 ;
      LAYER met2 ;
        RECT 1712.670 1700.000 1712.950 1704.000 ;
        RECT 1712.740 1688.770 1712.880 1700.000 ;
        RECT 1712.680 1688.450 1712.940 1688.770 ;
        RECT 1716.820 1688.450 1717.080 1688.770 ;
        RECT 1716.880 44.190 1717.020 1688.450 ;
        RECT 1716.820 43.870 1717.080 44.190 ;
        RECT 2084.360 43.870 2084.620 44.190 ;
        RECT 2084.420 2.400 2084.560 43.870 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1717.250 44.440 1717.570 44.500 ;
        RECT 2101.810 44.440 2102.130 44.500 ;
        RECT 1717.250 44.300 2102.130 44.440 ;
        RECT 1717.250 44.240 1717.570 44.300 ;
        RECT 2101.810 44.240 2102.130 44.300 ;
      LAYER via ;
        RECT 1717.280 44.240 1717.540 44.500 ;
        RECT 2101.840 44.240 2102.100 44.500 ;
      LAYER met2 ;
        RECT 1717.270 1700.000 1717.550 1704.000 ;
        RECT 1717.340 44.530 1717.480 1700.000 ;
        RECT 1717.280 44.210 1717.540 44.530 ;
        RECT 2101.840 44.210 2102.100 44.530 ;
        RECT 2101.900 2.400 2102.040 44.210 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1722.310 1688.340 1722.630 1688.400 ;
        RECT 1724.150 1688.340 1724.470 1688.400 ;
        RECT 1722.310 1688.200 1724.470 1688.340 ;
        RECT 1722.310 1688.140 1722.630 1688.200 ;
        RECT 1724.150 1688.140 1724.470 1688.200 ;
        RECT 1724.150 48.180 1724.470 48.240 ;
        RECT 2119.750 48.180 2120.070 48.240 ;
        RECT 1724.150 48.040 2120.070 48.180 ;
        RECT 1724.150 47.980 1724.470 48.040 ;
        RECT 2119.750 47.980 2120.070 48.040 ;
      LAYER via ;
        RECT 1722.340 1688.140 1722.600 1688.400 ;
        RECT 1724.180 1688.140 1724.440 1688.400 ;
        RECT 1724.180 47.980 1724.440 48.240 ;
        RECT 2119.780 47.980 2120.040 48.240 ;
      LAYER met2 ;
        RECT 1722.330 1700.000 1722.610 1704.000 ;
        RECT 1722.400 1688.430 1722.540 1700.000 ;
        RECT 1722.340 1688.110 1722.600 1688.430 ;
        RECT 1724.180 1688.110 1724.440 1688.430 ;
        RECT 1724.240 48.270 1724.380 1688.110 ;
        RECT 1724.180 47.950 1724.440 48.270 ;
        RECT 2119.780 47.950 2120.040 48.270 ;
        RECT 2119.840 2.400 2119.980 47.950 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 0.300 ;
=======
      LAYER met1 ;
        RECT 1726.910 1688.340 1727.230 1688.400 ;
        RECT 1730.130 1688.340 1730.450 1688.400 ;
        RECT 1726.910 1688.200 1730.450 1688.340 ;
        RECT 1726.910 1688.140 1727.230 1688.200 ;
        RECT 1730.130 1688.140 1730.450 1688.200 ;
        RECT 1730.130 47.840 1730.450 47.900 ;
        RECT 2137.690 47.840 2138.010 47.900 ;
        RECT 1730.130 47.700 2138.010 47.840 ;
        RECT 1730.130 47.640 1730.450 47.700 ;
        RECT 2137.690 47.640 2138.010 47.700 ;
      LAYER via ;
        RECT 1726.940 1688.140 1727.200 1688.400 ;
        RECT 1730.160 1688.140 1730.420 1688.400 ;
        RECT 1730.160 47.640 1730.420 47.900 ;
        RECT 2137.720 47.640 2137.980 47.900 ;
      LAYER met2 ;
        RECT 1726.930 1700.000 1727.210 1704.000 ;
        RECT 1727.000 1688.430 1727.140 1700.000 ;
        RECT 1726.940 1688.110 1727.200 1688.430 ;
        RECT 1730.160 1688.110 1730.420 1688.430 ;
        RECT 1730.220 47.930 1730.360 1688.110 ;
        RECT 1730.160 47.610 1730.420 47.930 ;
        RECT 2137.720 47.610 2137.980 47.930 ;
        RECT 2137.780 2.400 2137.920 47.610 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 0.300 ;
=======
      LAYER met1 ;
        RECT 1731.970 1688.340 1732.290 1688.400 ;
        RECT 1737.950 1688.340 1738.270 1688.400 ;
        RECT 1731.970 1688.200 1738.270 1688.340 ;
        RECT 1731.970 1688.140 1732.290 1688.200 ;
        RECT 1737.950 1688.140 1738.270 1688.200 ;
        RECT 1737.950 47.500 1738.270 47.560 ;
        RECT 2155.630 47.500 2155.950 47.560 ;
        RECT 1737.950 47.360 2155.950 47.500 ;
        RECT 1737.950 47.300 1738.270 47.360 ;
        RECT 2155.630 47.300 2155.950 47.360 ;
      LAYER via ;
        RECT 1732.000 1688.140 1732.260 1688.400 ;
        RECT 1737.980 1688.140 1738.240 1688.400 ;
        RECT 1737.980 47.300 1738.240 47.560 ;
        RECT 2155.660 47.300 2155.920 47.560 ;
      LAYER met2 ;
        RECT 1731.990 1700.000 1732.270 1704.000 ;
        RECT 1732.060 1688.430 1732.200 1700.000 ;
        RECT 1732.000 1688.110 1732.260 1688.430 ;
        RECT 1737.980 1688.110 1738.240 1688.430 ;
        RECT 1738.040 47.590 1738.180 1688.110 ;
        RECT 1737.980 47.270 1738.240 47.590 ;
        RECT 2155.660 47.270 2155.920 47.590 ;
        RECT 2155.720 2.400 2155.860 47.270 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1737.490 47.160 1737.810 47.220 ;
        RECT 2173.110 47.160 2173.430 47.220 ;
        RECT 1737.490 47.020 2173.430 47.160 ;
        RECT 1737.490 46.960 1737.810 47.020 ;
        RECT 2173.110 46.960 2173.430 47.020 ;
      LAYER via ;
        RECT 1737.520 46.960 1737.780 47.220 ;
        RECT 2173.140 46.960 2173.400 47.220 ;
      LAYER met2 ;
        RECT 1736.590 1700.410 1736.870 1704.000 ;
        RECT 1736.590 1700.270 1737.720 1700.410 ;
        RECT 1736.590 1700.000 1736.870 1700.270 ;
        RECT 1737.580 47.250 1737.720 1700.270 ;
        RECT 1737.520 46.930 1737.780 47.250 ;
        RECT 2173.140 46.930 2173.400 47.250 ;
        RECT 2173.200 2.400 2173.340 46.930 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1741.630 1688.340 1741.950 1688.400 ;
        RECT 1744.390 1688.340 1744.710 1688.400 ;
        RECT 1741.630 1688.200 1744.710 1688.340 ;
        RECT 1741.630 1688.140 1741.950 1688.200 ;
        RECT 1744.390 1688.140 1744.710 1688.200 ;
        RECT 1744.390 46.820 1744.710 46.880 ;
        RECT 2191.050 46.820 2191.370 46.880 ;
        RECT 1744.390 46.680 2191.370 46.820 ;
        RECT 1744.390 46.620 1744.710 46.680 ;
        RECT 2191.050 46.620 2191.370 46.680 ;
      LAYER via ;
        RECT 1741.660 1688.140 1741.920 1688.400 ;
        RECT 1744.420 1688.140 1744.680 1688.400 ;
        RECT 1744.420 46.620 1744.680 46.880 ;
        RECT 2191.080 46.620 2191.340 46.880 ;
      LAYER met2 ;
        RECT 1741.650 1700.000 1741.930 1704.000 ;
        RECT 1741.720 1688.430 1741.860 1700.000 ;
        RECT 1741.660 1688.110 1741.920 1688.430 ;
        RECT 1744.420 1688.110 1744.680 1688.430 ;
        RECT 1744.480 46.910 1744.620 1688.110 ;
        RECT 1744.420 46.590 1744.680 46.910 ;
        RECT 2191.080 46.590 2191.340 46.910 ;
        RECT 2191.140 2.400 2191.280 46.590 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1746.230 1688.340 1746.550 1688.400 ;
        RECT 1750.830 1688.340 1751.150 1688.400 ;
        RECT 1746.230 1688.200 1751.150 1688.340 ;
        RECT 1746.230 1688.140 1746.550 1688.200 ;
        RECT 1750.830 1688.140 1751.150 1688.200 ;
        RECT 1750.830 46.480 1751.150 46.540 ;
        RECT 2208.990 46.480 2209.310 46.540 ;
        RECT 1750.830 46.340 2209.310 46.480 ;
        RECT 1750.830 46.280 1751.150 46.340 ;
        RECT 2208.990 46.280 2209.310 46.340 ;
      LAYER via ;
        RECT 1746.260 1688.140 1746.520 1688.400 ;
        RECT 1750.860 1688.140 1751.120 1688.400 ;
        RECT 1750.860 46.280 1751.120 46.540 ;
        RECT 2209.020 46.280 2209.280 46.540 ;
      LAYER met2 ;
        RECT 1746.250 1700.000 1746.530 1704.000 ;
        RECT 1746.320 1688.430 1746.460 1700.000 ;
        RECT 1746.260 1688.110 1746.520 1688.430 ;
        RECT 1750.860 1688.110 1751.120 1688.430 ;
        RECT 1750.920 46.570 1751.060 1688.110 ;
        RECT 1750.860 46.250 1751.120 46.570 ;
        RECT 2209.020 46.250 2209.280 46.570 ;
        RECT 2209.080 2.400 2209.220 46.250 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 0.300 ;
=======
      LAYER met1 ;
        RECT 1751.290 46.140 1751.610 46.200 ;
        RECT 2226.930 46.140 2227.250 46.200 ;
        RECT 1751.290 46.000 2227.250 46.140 ;
        RECT 1751.290 45.940 1751.610 46.000 ;
        RECT 2226.930 45.940 2227.250 46.000 ;
      LAYER via ;
        RECT 1751.320 45.940 1751.580 46.200 ;
        RECT 2226.960 45.940 2227.220 46.200 ;
      LAYER met2 ;
        RECT 1750.850 1700.410 1751.130 1704.000 ;
        RECT 1750.850 1700.270 1751.520 1700.410 ;
        RECT 1750.850 1700.000 1751.130 1700.270 ;
        RECT 1751.380 46.230 1751.520 1700.270 ;
        RECT 1751.320 45.910 1751.580 46.230 ;
        RECT 2226.960 45.910 2227.220 46.230 ;
        RECT 2227.020 2.400 2227.160 45.910 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 0.300 ;
=======
      LAYER met1 ;
        RECT 781.610 40.700 781.930 40.760 ;
        RECT 1359.370 40.700 1359.690 40.760 ;
        RECT 781.610 40.560 1359.690 40.700 ;
        RECT 781.610 40.500 781.930 40.560 ;
        RECT 1359.370 40.500 1359.690 40.560 ;
      LAYER via ;
        RECT 781.640 40.500 781.900 40.760 ;
        RECT 1359.400 40.500 1359.660 40.760 ;
      LAYER met2 ;
        RECT 1360.770 1700.410 1361.050 1704.000 ;
        RECT 1359.460 1700.270 1361.050 1700.410 ;
        RECT 1359.460 40.790 1359.600 1700.270 ;
        RECT 1360.770 1700.000 1361.050 1700.270 ;
        RECT 781.640 40.470 781.900 40.790 ;
        RECT 1359.400 40.470 1359.660 40.790 ;
        RECT 781.700 2.400 781.840 40.470 ;
        RECT 781.490 -4.800 782.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1755.890 1688.340 1756.210 1688.400 ;
        RECT 1757.730 1688.340 1758.050 1688.400 ;
        RECT 1755.890 1688.200 1758.050 1688.340 ;
        RECT 1755.890 1688.140 1756.210 1688.200 ;
        RECT 1757.730 1688.140 1758.050 1688.200 ;
        RECT 1757.730 45.800 1758.050 45.860 ;
        RECT 2244.870 45.800 2245.190 45.860 ;
        RECT 1757.730 45.660 2245.190 45.800 ;
        RECT 1757.730 45.600 1758.050 45.660 ;
        RECT 2244.870 45.600 2245.190 45.660 ;
      LAYER via ;
        RECT 1755.920 1688.140 1756.180 1688.400 ;
        RECT 1757.760 1688.140 1758.020 1688.400 ;
        RECT 1757.760 45.600 1758.020 45.860 ;
        RECT 2244.900 45.600 2245.160 45.860 ;
      LAYER met2 ;
        RECT 1755.910 1700.000 1756.190 1704.000 ;
        RECT 1755.980 1688.430 1756.120 1700.000 ;
        RECT 1755.920 1688.110 1756.180 1688.430 ;
        RECT 1757.760 1688.110 1758.020 1688.430 ;
        RECT 1757.820 45.890 1757.960 1688.110 ;
        RECT 1757.760 45.570 1758.020 45.890 ;
        RECT 2244.900 45.570 2245.160 45.890 ;
        RECT 2244.960 2.400 2245.100 45.570 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 0.300 ;
=======
      LAYER met1 ;
        RECT 1760.490 1688.680 1760.810 1688.740 ;
        RECT 1765.550 1688.680 1765.870 1688.740 ;
        RECT 1760.490 1688.540 1765.870 1688.680 ;
        RECT 1760.490 1688.480 1760.810 1688.540 ;
        RECT 1765.550 1688.480 1765.870 1688.540 ;
        RECT 1765.550 45.460 1765.870 45.520 ;
        RECT 2262.350 45.460 2262.670 45.520 ;
        RECT 1765.550 45.320 2262.670 45.460 ;
        RECT 1765.550 45.260 1765.870 45.320 ;
        RECT 2262.350 45.260 2262.670 45.320 ;
      LAYER via ;
        RECT 1760.520 1688.480 1760.780 1688.740 ;
        RECT 1765.580 1688.480 1765.840 1688.740 ;
        RECT 1765.580 45.260 1765.840 45.520 ;
        RECT 2262.380 45.260 2262.640 45.520 ;
      LAYER met2 ;
        RECT 1760.510 1700.000 1760.790 1704.000 ;
        RECT 1760.580 1688.770 1760.720 1700.000 ;
        RECT 1760.520 1688.450 1760.780 1688.770 ;
        RECT 1765.580 1688.450 1765.840 1688.770 ;
        RECT 1765.640 45.550 1765.780 1688.450 ;
        RECT 1765.580 45.230 1765.840 45.550 ;
        RECT 2262.380 45.230 2262.640 45.550 ;
        RECT 2262.440 2.400 2262.580 45.230 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1765.090 45.120 1765.410 45.180 ;
        RECT 2280.290 45.120 2280.610 45.180 ;
        RECT 1765.090 44.980 2280.610 45.120 ;
        RECT 1765.090 44.920 1765.410 44.980 ;
        RECT 2280.290 44.920 2280.610 44.980 ;
      LAYER via ;
        RECT 1765.120 44.920 1765.380 45.180 ;
        RECT 2280.320 44.920 2280.580 45.180 ;
      LAYER met2 ;
        RECT 1765.570 1700.410 1765.850 1704.000 ;
        RECT 1765.180 1700.270 1765.850 1700.410 ;
        RECT 1765.180 45.210 1765.320 1700.270 ;
        RECT 1765.570 1700.000 1765.850 1700.270 ;
        RECT 1765.120 44.890 1765.380 45.210 ;
        RECT 2280.320 44.890 2280.580 45.210 ;
        RECT 2280.380 2.400 2280.520 44.890 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1771.990 50.900 1772.310 50.960 ;
        RECT 2298.230 50.900 2298.550 50.960 ;
        RECT 1771.990 50.760 2298.550 50.900 ;
        RECT 1771.990 50.700 1772.310 50.760 ;
        RECT 2298.230 50.700 2298.550 50.760 ;
      LAYER via ;
        RECT 1772.020 50.700 1772.280 50.960 ;
        RECT 2298.260 50.700 2298.520 50.960 ;
      LAYER met2 ;
        RECT 1770.170 1700.410 1770.450 1704.000 ;
        RECT 1770.170 1700.270 1771.300 1700.410 ;
        RECT 1770.170 1700.000 1770.450 1700.270 ;
        RECT 1771.160 1687.490 1771.300 1700.270 ;
        RECT 1771.160 1687.350 1772.220 1687.490 ;
        RECT 1772.080 50.990 1772.220 1687.350 ;
        RECT 1772.020 50.670 1772.280 50.990 ;
        RECT 2298.260 50.670 2298.520 50.990 ;
        RECT 2298.320 2.400 2298.460 50.670 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1775.210 1685.280 1775.530 1685.340 ;
        RECT 1778.430 1685.280 1778.750 1685.340 ;
        RECT 1775.210 1685.140 1778.750 1685.280 ;
        RECT 1775.210 1685.080 1775.530 1685.140 ;
        RECT 1778.430 1685.080 1778.750 1685.140 ;
        RECT 1778.430 51.240 1778.750 51.300 ;
        RECT 2311.570 51.240 2311.890 51.300 ;
        RECT 1778.430 51.100 2311.890 51.240 ;
        RECT 1778.430 51.040 1778.750 51.100 ;
        RECT 2311.570 51.040 2311.890 51.100 ;
      LAYER via ;
        RECT 1775.240 1685.080 1775.500 1685.340 ;
        RECT 1778.460 1685.080 1778.720 1685.340 ;
        RECT 1778.460 51.040 1778.720 51.300 ;
        RECT 2311.600 51.040 2311.860 51.300 ;
      LAYER met2 ;
        RECT 1775.230 1700.000 1775.510 1704.000 ;
        RECT 1775.300 1685.370 1775.440 1700.000 ;
        RECT 1775.240 1685.050 1775.500 1685.370 ;
        RECT 1778.460 1685.050 1778.720 1685.370 ;
        RECT 1778.520 51.330 1778.660 1685.050 ;
        RECT 1778.460 51.010 1778.720 51.330 ;
        RECT 2311.600 51.010 2311.860 51.330 ;
        RECT 2311.660 16.730 2311.800 51.010 ;
        RECT 2311.660 16.590 2316.400 16.730 ;
        RECT 2316.260 2.400 2316.400 16.590 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1777.970 1689.020 1778.290 1689.080 ;
        RECT 1779.810 1689.020 1780.130 1689.080 ;
        RECT 1777.970 1688.880 1780.130 1689.020 ;
        RECT 1777.970 1688.820 1778.290 1688.880 ;
        RECT 1779.810 1688.820 1780.130 1688.880 ;
        RECT 1777.970 54.980 1778.290 55.040 ;
        RECT 2332.270 54.980 2332.590 55.040 ;
        RECT 1777.970 54.840 2332.590 54.980 ;
        RECT 1777.970 54.780 1778.290 54.840 ;
        RECT 2332.270 54.780 2332.590 54.840 ;
      LAYER via ;
        RECT 1778.000 1688.820 1778.260 1689.080 ;
        RECT 1779.840 1688.820 1780.100 1689.080 ;
        RECT 1778.000 54.780 1778.260 55.040 ;
        RECT 2332.300 54.780 2332.560 55.040 ;
      LAYER met2 ;
        RECT 1779.830 1700.000 1780.110 1704.000 ;
        RECT 1779.900 1689.110 1780.040 1700.000 ;
        RECT 1778.000 1688.790 1778.260 1689.110 ;
        RECT 1779.840 1688.790 1780.100 1689.110 ;
        RECT 1778.060 55.070 1778.200 1688.790 ;
        RECT 1778.000 54.750 1778.260 55.070 ;
        RECT 2332.300 54.750 2332.560 55.070 ;
        RECT 2332.360 16.730 2332.500 54.750 ;
        RECT 2332.360 16.590 2334.340 16.730 ;
        RECT 2334.200 2.400 2334.340 16.590 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1785.790 54.640 1786.110 54.700 ;
        RECT 2346.070 54.640 2346.390 54.700 ;
        RECT 1785.790 54.500 2346.390 54.640 ;
        RECT 1785.790 54.440 1786.110 54.500 ;
        RECT 2346.070 54.440 2346.390 54.500 ;
      LAYER via ;
        RECT 1785.820 54.440 1786.080 54.700 ;
        RECT 2346.100 54.440 2346.360 54.700 ;
      LAYER met2 ;
        RECT 1784.890 1700.410 1785.170 1704.000 ;
        RECT 1784.890 1700.270 1786.020 1700.410 ;
        RECT 1784.890 1700.000 1785.170 1700.270 ;
        RECT 1785.880 54.730 1786.020 1700.270 ;
        RECT 1785.820 54.410 1786.080 54.730 ;
        RECT 2346.100 54.410 2346.360 54.730 ;
        RECT 2346.160 16.730 2346.300 54.410 ;
        RECT 2346.160 16.590 2351.820 16.730 ;
        RECT 2351.680 2.400 2351.820 16.590 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 0.300 ;
=======
      LAYER met1 ;
        RECT 1789.470 1684.600 1789.790 1684.660 ;
        RECT 1792.690 1684.600 1793.010 1684.660 ;
        RECT 1789.470 1684.460 1793.010 1684.600 ;
        RECT 1789.470 1684.400 1789.790 1684.460 ;
        RECT 1792.690 1684.400 1793.010 1684.460 ;
        RECT 1792.690 54.300 1793.010 54.360 ;
        RECT 2366.770 54.300 2367.090 54.360 ;
        RECT 1792.690 54.160 2367.090 54.300 ;
        RECT 1792.690 54.100 1793.010 54.160 ;
        RECT 2366.770 54.100 2367.090 54.160 ;
      LAYER via ;
        RECT 1789.500 1684.400 1789.760 1684.660 ;
        RECT 1792.720 1684.400 1792.980 1684.660 ;
        RECT 1792.720 54.100 1792.980 54.360 ;
        RECT 2366.800 54.100 2367.060 54.360 ;
      LAYER met2 ;
        RECT 1789.490 1700.000 1789.770 1704.000 ;
        RECT 1789.560 1684.690 1789.700 1700.000 ;
        RECT 1789.500 1684.370 1789.760 1684.690 ;
        RECT 1792.720 1684.370 1792.980 1684.690 ;
        RECT 1792.780 54.390 1792.920 1684.370 ;
        RECT 1792.720 54.070 1792.980 54.390 ;
        RECT 2366.800 54.070 2367.060 54.390 ;
        RECT 2366.860 16.730 2367.000 54.070 ;
        RECT 2366.860 16.590 2369.760 16.730 ;
        RECT 2369.620 2.400 2369.760 16.590 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1794.530 1687.660 1794.850 1687.720 ;
        RECT 1799.590 1687.660 1799.910 1687.720 ;
        RECT 1794.530 1687.520 1799.910 1687.660 ;
        RECT 1794.530 1687.460 1794.850 1687.520 ;
        RECT 1799.590 1687.460 1799.910 1687.520 ;
        RECT 1799.590 53.960 1799.910 54.020 ;
        RECT 2387.930 53.960 2388.250 54.020 ;
        RECT 1799.590 53.820 2388.250 53.960 ;
        RECT 1799.590 53.760 1799.910 53.820 ;
        RECT 2387.930 53.760 2388.250 53.820 ;
      LAYER via ;
        RECT 1794.560 1687.460 1794.820 1687.720 ;
        RECT 1799.620 1687.460 1799.880 1687.720 ;
        RECT 1799.620 53.760 1799.880 54.020 ;
        RECT 2387.960 53.760 2388.220 54.020 ;
      LAYER met2 ;
        RECT 1794.550 1700.000 1794.830 1704.000 ;
        RECT 1794.620 1687.750 1794.760 1700.000 ;
        RECT 1794.560 1687.430 1794.820 1687.750 ;
        RECT 1799.620 1687.430 1799.880 1687.750 ;
        RECT 1799.680 54.050 1799.820 1687.430 ;
        RECT 1799.620 53.730 1799.880 54.050 ;
        RECT 2387.960 53.730 2388.220 54.050 ;
        RECT 2388.020 17.410 2388.160 53.730 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1799.130 53.620 1799.450 53.680 ;
        RECT 2401.270 53.620 2401.590 53.680 ;
        RECT 1799.130 53.480 2401.590 53.620 ;
        RECT 1799.130 53.420 1799.450 53.480 ;
        RECT 2401.270 53.420 2401.590 53.480 ;
        RECT 2401.270 2.960 2401.590 3.020 ;
        RECT 2405.410 2.960 2405.730 3.020 ;
        RECT 2401.270 2.820 2405.730 2.960 ;
        RECT 2401.270 2.760 2401.590 2.820 ;
        RECT 2405.410 2.760 2405.730 2.820 ;
      LAYER via ;
        RECT 1799.160 53.420 1799.420 53.680 ;
        RECT 2401.300 53.420 2401.560 53.680 ;
        RECT 2401.300 2.760 2401.560 3.020 ;
        RECT 2405.440 2.760 2405.700 3.020 ;
      LAYER met2 ;
        RECT 1799.150 1700.000 1799.430 1704.000 ;
        RECT 1799.220 53.710 1799.360 1700.000 ;
        RECT 1799.160 53.390 1799.420 53.710 ;
        RECT 2401.300 53.390 2401.560 53.710 ;
        RECT 2401.360 3.050 2401.500 53.390 ;
        RECT 2401.300 2.730 2401.560 3.050 ;
        RECT 2405.440 2.730 2405.700 3.050 ;
        RECT 2405.500 2.400 2405.640 2.730 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1359.830 1678.140 1360.150 1678.200 ;
        RECT 1364.430 1678.140 1364.750 1678.200 ;
        RECT 1359.830 1678.000 1364.750 1678.140 ;
        RECT 1359.830 1677.940 1360.150 1678.000 ;
        RECT 1364.430 1677.940 1364.750 1678.000 ;
        RECT 799.550 41.040 799.870 41.100 ;
        RECT 1359.830 41.040 1360.150 41.100 ;
        RECT 799.550 40.900 1360.150 41.040 ;
        RECT 799.550 40.840 799.870 40.900 ;
        RECT 1359.830 40.840 1360.150 40.900 ;
      LAYER via ;
        RECT 1359.860 1677.940 1360.120 1678.200 ;
        RECT 1364.460 1677.940 1364.720 1678.200 ;
        RECT 799.580 40.840 799.840 41.100 ;
        RECT 1359.860 40.840 1360.120 41.100 ;
      LAYER met2 ;
        RECT 1365.370 1700.410 1365.650 1704.000 ;
        RECT 1364.520 1700.270 1365.650 1700.410 ;
        RECT 1364.520 1678.230 1364.660 1700.270 ;
        RECT 1365.370 1700.000 1365.650 1700.270 ;
        RECT 1359.860 1677.910 1360.120 1678.230 ;
        RECT 1364.460 1677.910 1364.720 1678.230 ;
        RECT 1359.920 41.130 1360.060 1677.910 ;
        RECT 799.580 40.810 799.840 41.130 ;
        RECT 1359.860 40.810 1360.120 41.130 ;
        RECT 799.640 2.400 799.780 40.810 ;
        RECT 799.430 -4.800 799.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1320.270 1642.440 1320.590 1642.500 ;
        RECT 1323.030 1642.440 1323.350 1642.500 ;
        RECT 1320.270 1642.300 1323.350 1642.440 ;
        RECT 1320.270 1642.240 1320.590 1642.300 ;
        RECT 1323.030 1642.240 1323.350 1642.300 ;
      LAYER via ;
        RECT 1320.300 1642.240 1320.560 1642.500 ;
        RECT 1323.060 1642.240 1323.320 1642.500 ;
      LAYER met2 ;
        RECT 1323.970 1700.410 1324.250 1704.000 ;
        RECT 1323.120 1700.270 1324.250 1700.410 ;
        RECT 1323.120 1642.530 1323.260 1700.270 ;
        RECT 1323.970 1700.000 1324.250 1700.270 ;
        RECT 1320.300 1642.210 1320.560 1642.530 ;
        RECT 1323.060 1642.210 1323.320 1642.530 ;
        RECT 1320.360 41.325 1320.500 1642.210 ;
        RECT 645.010 40.955 645.290 41.325 ;
        RECT 1320.290 40.955 1320.570 41.325 ;
        RECT 645.080 2.400 645.220 40.955 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 645.010 41.000 645.290 41.280 ;
        RECT 1320.290 41.000 1320.570 41.280 ;
      LAYER met3 ;
        RECT 644.985 41.290 645.315 41.305 ;
        RECT 1320.265 41.290 1320.595 41.305 ;
        RECT 644.985 40.990 1320.595 41.290 ;
        RECT 644.985 40.975 645.315 40.990 ;
        RECT 1320.265 40.975 1320.595 40.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1806.030 53.280 1806.350 53.340 ;
        RECT 2428.870 53.280 2429.190 53.340 ;
        RECT 1806.030 53.140 2429.190 53.280 ;
        RECT 1806.030 53.080 1806.350 53.140 ;
        RECT 2428.870 53.080 2429.190 53.140 ;
      LAYER via ;
        RECT 1806.060 53.080 1806.320 53.340 ;
        RECT 2428.900 53.080 2429.160 53.340 ;
      LAYER met2 ;
        RECT 1805.590 1700.410 1805.870 1704.000 ;
        RECT 1805.590 1700.270 1806.260 1700.410 ;
        RECT 1805.590 1700.000 1805.870 1700.270 ;
        RECT 1806.120 53.370 1806.260 1700.270 ;
        RECT 1806.060 53.050 1806.320 53.370 ;
        RECT 2428.900 53.050 2429.160 53.370 ;
        RECT 2428.960 2.400 2429.100 53.050 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1812.930 52.940 1813.250 53.000 ;
        RECT 2442.670 52.940 2442.990 53.000 ;
        RECT 1812.930 52.800 2442.990 52.940 ;
        RECT 1812.930 52.740 1813.250 52.800 ;
        RECT 2442.670 52.740 2442.990 52.800 ;
        RECT 2442.670 2.960 2442.990 3.020 ;
        RECT 2446.810 2.960 2447.130 3.020 ;
        RECT 2442.670 2.820 2447.130 2.960 ;
        RECT 2442.670 2.760 2442.990 2.820 ;
        RECT 2446.810 2.760 2447.130 2.820 ;
      LAYER via ;
        RECT 1812.960 52.740 1813.220 53.000 ;
        RECT 2442.700 52.740 2442.960 53.000 ;
        RECT 2442.700 2.760 2442.960 3.020 ;
        RECT 2446.840 2.760 2447.100 3.020 ;
      LAYER met2 ;
        RECT 1810.650 1700.410 1810.930 1704.000 ;
        RECT 1810.650 1700.270 1811.320 1700.410 ;
        RECT 1810.650 1700.000 1810.930 1700.270 ;
        RECT 1811.180 1677.970 1811.320 1700.270 ;
        RECT 1811.180 1677.830 1813.160 1677.970 ;
        RECT 1813.020 53.030 1813.160 1677.830 ;
        RECT 1812.960 52.710 1813.220 53.030 ;
        RECT 2442.700 52.710 2442.960 53.030 ;
        RECT 2442.760 3.050 2442.900 52.710 ;
        RECT 2442.700 2.730 2442.960 3.050 ;
        RECT 2446.840 2.730 2447.100 3.050 ;
        RECT 2446.900 2.400 2447.040 2.730 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1815.230 1683.920 1815.550 1683.980 ;
        RECT 1819.370 1683.920 1819.690 1683.980 ;
        RECT 1815.230 1683.780 1819.690 1683.920 ;
        RECT 1815.230 1683.720 1815.550 1683.780 ;
        RECT 1819.370 1683.720 1819.690 1683.780 ;
        RECT 1819.830 52.600 1820.150 52.660 ;
        RECT 2463.370 52.600 2463.690 52.660 ;
        RECT 1819.830 52.460 2463.690 52.600 ;
        RECT 1819.830 52.400 1820.150 52.460 ;
        RECT 2463.370 52.400 2463.690 52.460 ;
        RECT 2463.370 2.960 2463.690 3.020 ;
        RECT 2464.750 2.960 2465.070 3.020 ;
        RECT 2463.370 2.820 2465.070 2.960 ;
        RECT 2463.370 2.760 2463.690 2.820 ;
        RECT 2464.750 2.760 2465.070 2.820 ;
      LAYER via ;
        RECT 1815.260 1683.720 1815.520 1683.980 ;
        RECT 1819.400 1683.720 1819.660 1683.980 ;
        RECT 1819.860 52.400 1820.120 52.660 ;
        RECT 2463.400 52.400 2463.660 52.660 ;
        RECT 2463.400 2.760 2463.660 3.020 ;
        RECT 2464.780 2.760 2465.040 3.020 ;
      LAYER met2 ;
        RECT 1815.250 1700.000 1815.530 1704.000 ;
        RECT 1815.320 1684.010 1815.460 1700.000 ;
        RECT 1815.260 1683.690 1815.520 1684.010 ;
        RECT 1819.400 1683.690 1819.660 1684.010 ;
        RECT 1819.460 1669.810 1819.600 1683.690 ;
        RECT 1819.460 1669.670 1820.060 1669.810 ;
        RECT 1819.920 52.690 1820.060 1669.670 ;
        RECT 1819.860 52.370 1820.120 52.690 ;
        RECT 2463.400 52.370 2463.660 52.690 ;
        RECT 2463.460 3.050 2463.600 52.370 ;
        RECT 2463.400 2.730 2463.660 3.050 ;
        RECT 2464.780 2.730 2465.040 3.050 ;
        RECT 2464.840 2.400 2464.980 2.730 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 0.300 ;
=======
      LAYER li1 ;
        RECT 1825.425 19.125 1825.595 19.975 ;
      LAYER mcon ;
        RECT 1825.425 19.805 1825.595 19.975 ;
      LAYER met1 ;
        RECT 1825.365 19.960 1825.655 20.005 ;
        RECT 2482.690 19.960 2483.010 20.020 ;
        RECT 1825.365 19.820 2483.010 19.960 ;
        RECT 1825.365 19.775 1825.655 19.820 ;
        RECT 2482.690 19.760 2483.010 19.820 ;
        RECT 1821.210 19.280 1821.530 19.340 ;
        RECT 1825.365 19.280 1825.655 19.325 ;
        RECT 1821.210 19.140 1825.655 19.280 ;
        RECT 1821.210 19.080 1821.530 19.140 ;
        RECT 1825.365 19.095 1825.655 19.140 ;
      LAYER via ;
        RECT 2482.720 19.760 2482.980 20.020 ;
        RECT 1821.240 19.080 1821.500 19.340 ;
      LAYER met2 ;
        RECT 1820.310 1700.410 1820.590 1704.000 ;
        RECT 1820.310 1700.270 1821.440 1700.410 ;
        RECT 1820.310 1700.000 1820.590 1700.270 ;
        RECT 1821.300 19.370 1821.440 1700.270 ;
        RECT 2482.720 19.730 2482.980 20.050 ;
        RECT 1821.240 19.050 1821.500 19.370 ;
        RECT 2482.780 2.400 2482.920 19.730 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 0.300 ;
=======
      LAYER met1 ;
        RECT 1824.890 1684.260 1825.210 1684.320 ;
        RECT 1827.650 1684.260 1827.970 1684.320 ;
        RECT 1824.890 1684.120 1827.970 1684.260 ;
        RECT 1824.890 1684.060 1825.210 1684.120 ;
        RECT 1827.650 1684.060 1827.970 1684.120 ;
        RECT 1828.110 19.280 1828.430 19.340 ;
        RECT 2500.630 19.280 2500.950 19.340 ;
        RECT 1828.110 19.140 2500.950 19.280 ;
        RECT 1828.110 19.080 1828.430 19.140 ;
        RECT 2500.630 19.080 2500.950 19.140 ;
      LAYER via ;
        RECT 1824.920 1684.060 1825.180 1684.320 ;
        RECT 1827.680 1684.060 1827.940 1684.320 ;
        RECT 1828.140 19.080 1828.400 19.340 ;
        RECT 2500.660 19.080 2500.920 19.340 ;
      LAYER met2 ;
        RECT 1824.910 1700.000 1825.190 1704.000 ;
        RECT 1824.980 1684.350 1825.120 1700.000 ;
        RECT 1824.920 1684.030 1825.180 1684.350 ;
        RECT 1827.680 1684.030 1827.940 1684.350 ;
        RECT 1827.740 1677.970 1827.880 1684.030 ;
        RECT 1827.740 1677.830 1828.340 1677.970 ;
        RECT 1828.200 19.370 1828.340 1677.830 ;
        RECT 1828.140 19.050 1828.400 19.370 ;
        RECT 2500.660 19.050 2500.920 19.370 ;
        RECT 2500.720 2.400 2500.860 19.050 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 0.300 ;
=======
      LAYER li1 ;
        RECT 1847.965 1684.445 1848.135 1685.635 ;
        RECT 1866.365 1684.445 1869.755 1684.615 ;
        RECT 1869.585 1683.765 1869.755 1684.445 ;
        RECT 1938.585 1683.765 1939.675 1683.935 ;
      LAYER mcon ;
        RECT 1847.965 1685.465 1848.135 1685.635 ;
        RECT 1939.505 1683.765 1939.675 1683.935 ;
      LAYER met1 ;
        RECT 1829.950 1685.620 1830.270 1685.680 ;
        RECT 1847.905 1685.620 1848.195 1685.665 ;
        RECT 1829.950 1685.480 1848.195 1685.620 ;
        RECT 1829.950 1685.420 1830.270 1685.480 ;
        RECT 1847.905 1685.435 1848.195 1685.480 ;
        RECT 1847.905 1684.600 1848.195 1684.645 ;
        RECT 1866.305 1684.600 1866.595 1684.645 ;
        RECT 1847.905 1684.460 1866.595 1684.600 ;
        RECT 1847.905 1684.415 1848.195 1684.460 ;
        RECT 1866.305 1684.415 1866.595 1684.460 ;
        RECT 1869.525 1683.920 1869.815 1683.965 ;
        RECT 1938.525 1683.920 1938.815 1683.965 ;
        RECT 1869.525 1683.780 1938.815 1683.920 ;
        RECT 1869.525 1683.735 1869.815 1683.780 ;
        RECT 1938.525 1683.735 1938.815 1683.780 ;
        RECT 1939.445 1683.920 1939.735 1683.965 ;
        RECT 1969.790 1683.920 1970.110 1683.980 ;
        RECT 1939.445 1683.780 1970.110 1683.920 ;
        RECT 1939.445 1683.735 1939.735 1683.780 ;
        RECT 1969.790 1683.720 1970.110 1683.780 ;
        RECT 1969.790 15.200 1970.110 15.260 ;
        RECT 2518.110 15.200 2518.430 15.260 ;
        RECT 1969.790 15.060 2518.430 15.200 ;
        RECT 1969.790 15.000 1970.110 15.060 ;
        RECT 2518.110 15.000 2518.430 15.060 ;
      LAYER via ;
        RECT 1829.980 1685.420 1830.240 1685.680 ;
        RECT 1969.820 1683.720 1970.080 1683.980 ;
        RECT 1969.820 15.000 1970.080 15.260 ;
        RECT 2518.140 15.000 2518.400 15.260 ;
      LAYER met2 ;
        RECT 1829.970 1700.000 1830.250 1704.000 ;
        RECT 1830.040 1685.710 1830.180 1700.000 ;
        RECT 1829.980 1685.390 1830.240 1685.710 ;
        RECT 1969.820 1683.690 1970.080 1684.010 ;
        RECT 1969.880 15.290 1970.020 1683.690 ;
        RECT 1969.820 14.970 1970.080 15.290 ;
        RECT 2518.140 14.970 2518.400 15.290 ;
        RECT 2518.200 2.400 2518.340 14.970 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2535.930 -4.800 2536.490 0.300 ;
=======
        RECT 1834.570 1700.410 1834.850 1704.000 ;
        RECT 1834.570 1700.270 1835.240 1700.410 ;
        RECT 1834.570 1700.000 1834.850 1700.270 ;
        RECT 1835.100 19.565 1835.240 1700.270 ;
        RECT 1835.030 19.195 1835.310 19.565 ;
        RECT 2536.070 19.195 2536.350 19.565 ;
        RECT 2536.140 2.400 2536.280 19.195 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
      LAYER via2 ;
        RECT 1835.030 19.240 1835.310 19.520 ;
        RECT 2536.070 19.240 2536.350 19.520 ;
      LAYER met3 ;
        RECT 1835.005 19.530 1835.335 19.545 ;
        RECT 2536.045 19.530 2536.375 19.545 ;
        RECT 1835.005 19.230 2536.375 19.530 ;
        RECT 1835.005 19.215 1835.335 19.230 ;
        RECT 2536.045 19.215 2536.375 19.230 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 0.300 ;
=======
      LAYER li1 ;
        RECT 1848.885 1683.765 1849.055 1685.975 ;
        RECT 1870.505 1683.085 1870.675 1684.615 ;
      LAYER mcon ;
        RECT 1848.885 1685.805 1849.055 1685.975 ;
        RECT 1870.505 1684.445 1870.675 1684.615 ;
      LAYER met1 ;
        RECT 1839.610 1685.960 1839.930 1686.020 ;
        RECT 1848.825 1685.960 1849.115 1686.005 ;
        RECT 1839.610 1685.820 1849.115 1685.960 ;
        RECT 1839.610 1685.760 1839.930 1685.820 ;
        RECT 1848.825 1685.775 1849.115 1685.820 ;
        RECT 1870.445 1684.600 1870.735 1684.645 ;
        RECT 2004.290 1684.600 2004.610 1684.660 ;
        RECT 1870.445 1684.460 2004.610 1684.600 ;
        RECT 1870.445 1684.415 1870.735 1684.460 ;
        RECT 2004.290 1684.400 2004.610 1684.460 ;
        RECT 1848.825 1683.920 1849.115 1683.965 ;
        RECT 1848.825 1683.780 1869.280 1683.920 ;
        RECT 1848.825 1683.735 1849.115 1683.780 ;
        RECT 1869.140 1683.240 1869.280 1683.780 ;
        RECT 1870.445 1683.240 1870.735 1683.285 ;
        RECT 1869.140 1683.100 1870.735 1683.240 ;
        RECT 1870.445 1683.055 1870.735 1683.100 ;
        RECT 2004.290 15.540 2004.610 15.600 ;
        RECT 2553.990 15.540 2554.310 15.600 ;
        RECT 2004.290 15.400 2554.310 15.540 ;
        RECT 2004.290 15.340 2004.610 15.400 ;
        RECT 2553.990 15.340 2554.310 15.400 ;
      LAYER via ;
        RECT 1839.640 1685.760 1839.900 1686.020 ;
        RECT 2004.320 1684.400 2004.580 1684.660 ;
        RECT 2004.320 15.340 2004.580 15.600 ;
        RECT 2554.020 15.340 2554.280 15.600 ;
      LAYER met2 ;
        RECT 1839.630 1700.000 1839.910 1704.000 ;
        RECT 1839.700 1686.050 1839.840 1700.000 ;
        RECT 1839.640 1685.730 1839.900 1686.050 ;
        RECT 2004.320 1684.370 2004.580 1684.690 ;
        RECT 2004.380 15.630 2004.520 1684.370 ;
        RECT 2004.320 15.310 2004.580 15.630 ;
        RECT 2554.020 15.310 2554.280 15.630 ;
        RECT 2554.080 2.400 2554.220 15.310 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 0.300 ;
=======
      LAYER met1 ;
        RECT 1844.210 1684.600 1844.530 1684.660 ;
        RECT 1847.430 1684.600 1847.750 1684.660 ;
        RECT 1844.210 1684.460 1847.750 1684.600 ;
        RECT 1844.210 1684.400 1844.530 1684.460 ;
        RECT 1847.430 1684.400 1847.750 1684.460 ;
        RECT 1847.430 52.260 1847.750 52.320 ;
        RECT 2566.870 52.260 2567.190 52.320 ;
        RECT 1847.430 52.120 2567.190 52.260 ;
        RECT 1847.430 52.060 1847.750 52.120 ;
        RECT 2566.870 52.060 2567.190 52.120 ;
      LAYER via ;
        RECT 1844.240 1684.400 1844.500 1684.660 ;
        RECT 1847.460 1684.400 1847.720 1684.660 ;
        RECT 1847.460 52.060 1847.720 52.320 ;
        RECT 2566.900 52.060 2567.160 52.320 ;
      LAYER met2 ;
        RECT 1844.230 1700.000 1844.510 1704.000 ;
        RECT 1844.300 1684.690 1844.440 1700.000 ;
        RECT 1844.240 1684.370 1844.500 1684.690 ;
        RECT 1847.460 1684.370 1847.720 1684.690 ;
        RECT 1847.520 52.350 1847.660 1684.370 ;
        RECT 1847.460 52.030 1847.720 52.350 ;
        RECT 2566.900 52.030 2567.160 52.350 ;
        RECT 2566.960 16.730 2567.100 52.030 ;
        RECT 2566.960 16.590 2572.160 16.730 ;
        RECT 2572.020 2.400 2572.160 16.590 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 0.300 ;
=======
      LAYER li1 ;
        RECT 1867.745 1685.805 1868.835 1685.975 ;
        RECT 1868.665 1684.955 1868.835 1685.805 ;
        RECT 1874.185 1685.465 1874.355 1689.035 ;
        RECT 1868.665 1684.785 1869.755 1684.955 ;
        RECT 1897.645 1683.425 1897.815 1689.035 ;
      LAYER mcon ;
        RECT 1874.185 1688.865 1874.355 1689.035 ;
        RECT 1897.645 1688.865 1897.815 1689.035 ;
        RECT 1869.585 1684.785 1869.755 1684.955 ;
      LAYER met1 ;
        RECT 1874.125 1689.020 1874.415 1689.065 ;
        RECT 1897.585 1689.020 1897.875 1689.065 ;
        RECT 1874.125 1688.880 1897.875 1689.020 ;
        RECT 1874.125 1688.835 1874.415 1688.880 ;
        RECT 1897.585 1688.835 1897.875 1688.880 ;
        RECT 1867.685 1685.960 1867.975 1686.005 ;
        RECT 1856.720 1685.820 1867.975 1685.960 ;
        RECT 1849.270 1685.280 1849.590 1685.340 ;
        RECT 1856.720 1685.280 1856.860 1685.820 ;
        RECT 1867.685 1685.775 1867.975 1685.820 ;
        RECT 1874.125 1685.620 1874.415 1685.665 ;
        RECT 1870.060 1685.480 1874.415 1685.620 ;
        RECT 1870.060 1685.280 1870.200 1685.480 ;
        RECT 1874.125 1685.435 1874.415 1685.480 ;
        RECT 1849.270 1685.140 1856.860 1685.280 ;
        RECT 1869.600 1685.140 1870.200 1685.280 ;
        RECT 1849.270 1685.080 1849.590 1685.140 ;
        RECT 1869.600 1684.985 1869.740 1685.140 ;
        RECT 1869.525 1684.755 1869.815 1684.985 ;
        RECT 2004.750 1684.260 2005.070 1684.320 ;
        RECT 1939.060 1684.120 2005.070 1684.260 ;
        RECT 1897.585 1683.580 1897.875 1683.625 ;
        RECT 1939.060 1683.580 1939.200 1684.120 ;
        RECT 2004.750 1684.060 2005.070 1684.120 ;
        RECT 1897.585 1683.440 1939.200 1683.580 ;
        RECT 1897.585 1683.395 1897.875 1683.440 ;
        RECT 2004.750 16.220 2005.070 16.280 ;
        RECT 2589.410 16.220 2589.730 16.280 ;
        RECT 2004.750 16.080 2589.730 16.220 ;
        RECT 2004.750 16.020 2005.070 16.080 ;
        RECT 2589.410 16.020 2589.730 16.080 ;
      LAYER via ;
        RECT 1849.300 1685.080 1849.560 1685.340 ;
        RECT 2004.780 1684.060 2005.040 1684.320 ;
        RECT 2004.780 16.020 2005.040 16.280 ;
        RECT 2589.440 16.020 2589.700 16.280 ;
      LAYER met2 ;
        RECT 1849.290 1700.000 1849.570 1704.000 ;
        RECT 1849.360 1685.370 1849.500 1700.000 ;
        RECT 1849.300 1685.050 1849.560 1685.370 ;
        RECT 2004.780 1684.030 2005.040 1684.350 ;
        RECT 2004.840 16.310 2004.980 1684.030 ;
        RECT 2004.780 15.990 2005.040 16.310 ;
        RECT 2589.440 15.990 2589.700 16.310 ;
        RECT 2589.500 2.400 2589.640 15.990 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1366.730 1678.480 1367.050 1678.540 ;
        RECT 1370.870 1678.480 1371.190 1678.540 ;
        RECT 1366.730 1678.340 1371.190 1678.480 ;
        RECT 1366.730 1678.280 1367.050 1678.340 ;
        RECT 1370.870 1678.280 1371.190 1678.340 ;
        RECT 823.470 41.380 823.790 41.440 ;
        RECT 1200.670 41.380 1200.990 41.440 ;
        RECT 823.470 41.240 1200.990 41.380 ;
        RECT 823.470 41.180 823.790 41.240 ;
        RECT 1200.670 41.180 1200.990 41.240 ;
        RECT 1203.430 41.380 1203.750 41.440 ;
        RECT 1366.730 41.380 1367.050 41.440 ;
        RECT 1203.430 41.240 1367.050 41.380 ;
        RECT 1203.430 41.180 1203.750 41.240 ;
        RECT 1366.730 41.180 1367.050 41.240 ;
      LAYER via ;
        RECT 1366.760 1678.280 1367.020 1678.540 ;
        RECT 1370.900 1678.280 1371.160 1678.540 ;
        RECT 823.500 41.180 823.760 41.440 ;
        RECT 1200.700 41.180 1200.960 41.440 ;
        RECT 1203.460 41.180 1203.720 41.440 ;
        RECT 1366.760 41.180 1367.020 41.440 ;
      LAYER met2 ;
        RECT 1371.810 1700.410 1372.090 1704.000 ;
        RECT 1370.960 1700.270 1372.090 1700.410 ;
        RECT 1370.960 1678.570 1371.100 1700.270 ;
        RECT 1371.810 1700.000 1372.090 1700.270 ;
        RECT 1366.760 1678.250 1367.020 1678.570 ;
        RECT 1370.900 1678.250 1371.160 1678.570 ;
        RECT 1366.820 41.470 1366.960 1678.250 ;
        RECT 823.500 41.150 823.760 41.470 ;
        RECT 1200.700 41.150 1200.960 41.470 ;
        RECT 1203.460 41.150 1203.720 41.470 ;
        RECT 1366.760 41.150 1367.020 41.470 ;
        RECT 823.560 2.400 823.700 41.150 ;
        RECT 1200.760 40.645 1200.900 41.150 ;
        RECT 1203.520 40.645 1203.660 41.150 ;
        RECT 1200.690 40.275 1200.970 40.645 ;
        RECT 1203.450 40.275 1203.730 40.645 ;
        RECT 823.350 -4.800 823.910 2.400 ;
      LAYER via2 ;
        RECT 1200.690 40.320 1200.970 40.600 ;
        RECT 1203.450 40.320 1203.730 40.600 ;
      LAYER met3 ;
        RECT 1200.665 40.610 1200.995 40.625 ;
        RECT 1203.425 40.610 1203.755 40.625 ;
        RECT 1200.665 40.310 1203.755 40.610 ;
        RECT 1200.665 40.295 1200.995 40.310 ;
        RECT 1203.425 40.295 1203.755 40.310 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 0.300 ;
=======
      LAYER li1 ;
        RECT 1858.545 17.085 1858.715 18.955 ;
      LAYER mcon ;
        RECT 1858.545 18.785 1858.715 18.955 ;
      LAYER met1 ;
        RECT 1853.870 1686.640 1854.190 1686.700 ;
        RECT 1855.710 1686.640 1856.030 1686.700 ;
        RECT 1853.870 1686.500 1856.030 1686.640 ;
        RECT 1853.870 1686.440 1854.190 1686.500 ;
        RECT 1855.710 1686.440 1856.030 1686.500 ;
        RECT 1855.710 18.940 1856.030 19.000 ;
        RECT 1858.485 18.940 1858.775 18.985 ;
        RECT 1855.710 18.800 1858.775 18.940 ;
        RECT 1855.710 18.740 1856.030 18.800 ;
        RECT 1858.485 18.755 1858.775 18.800 ;
        RECT 2607.350 17.580 2607.670 17.640 ;
        RECT 1873.740 17.440 2607.670 17.580 ;
        RECT 1858.485 17.240 1858.775 17.285 ;
        RECT 1873.740 17.240 1873.880 17.440 ;
        RECT 2607.350 17.380 2607.670 17.440 ;
        RECT 1858.485 17.100 1873.880 17.240 ;
        RECT 1858.485 17.055 1858.775 17.100 ;
      LAYER via ;
        RECT 1853.900 1686.440 1854.160 1686.700 ;
        RECT 1855.740 1686.440 1856.000 1686.700 ;
        RECT 1855.740 18.740 1856.000 19.000 ;
        RECT 2607.380 17.380 2607.640 17.640 ;
      LAYER met2 ;
        RECT 1853.890 1700.000 1854.170 1704.000 ;
        RECT 1853.960 1686.730 1854.100 1700.000 ;
        RECT 1853.900 1686.410 1854.160 1686.730 ;
        RECT 1855.740 1686.410 1856.000 1686.730 ;
        RECT 1855.800 19.030 1855.940 1686.410 ;
        RECT 1855.740 18.710 1856.000 19.030 ;
        RECT 2607.380 17.350 2607.640 17.670 ;
        RECT 2607.440 2.400 2607.580 17.350 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 0.300 ;
=======
      LAYER li1 ;
        RECT 1869.125 1685.125 1869.295 1686.655 ;
        RECT 1870.505 1685.125 1870.675 1686.655 ;
        RECT 2087.165 16.405 2087.335 18.615 ;
      LAYER mcon ;
        RECT 1869.125 1686.485 1869.295 1686.655 ;
        RECT 1870.505 1686.485 1870.675 1686.655 ;
        RECT 2087.165 18.445 2087.335 18.615 ;
      LAYER met1 ;
        RECT 1869.065 1686.640 1869.355 1686.685 ;
        RECT 1870.445 1686.640 1870.735 1686.685 ;
        RECT 1869.065 1686.500 1870.735 1686.640 ;
        RECT 1869.065 1686.455 1869.355 1686.500 ;
        RECT 1870.445 1686.455 1870.735 1686.500 ;
        RECT 1858.470 1685.280 1858.790 1685.340 ;
        RECT 1869.065 1685.280 1869.355 1685.325 ;
        RECT 1858.470 1685.140 1869.355 1685.280 ;
        RECT 1858.470 1685.080 1858.790 1685.140 ;
        RECT 1869.065 1685.095 1869.355 1685.140 ;
        RECT 1870.445 1685.095 1870.735 1685.325 ;
        RECT 2038.790 1685.280 2039.110 1685.340 ;
        RECT 1890.760 1685.140 2039.110 1685.280 ;
        RECT 1870.520 1684.940 1870.660 1685.095 ;
        RECT 1890.760 1684.940 1890.900 1685.140 ;
        RECT 2038.790 1685.080 2039.110 1685.140 ;
        RECT 1870.520 1684.800 1890.900 1684.940 ;
        RECT 2039.250 18.600 2039.570 18.660 ;
        RECT 2087.105 18.600 2087.395 18.645 ;
        RECT 2039.250 18.460 2087.395 18.600 ;
        RECT 2039.250 18.400 2039.570 18.460 ;
        RECT 2087.105 18.415 2087.395 18.460 ;
        RECT 2087.105 16.560 2087.395 16.605 ;
        RECT 2625.290 16.560 2625.610 16.620 ;
        RECT 2087.105 16.420 2625.610 16.560 ;
        RECT 2087.105 16.375 2087.395 16.420 ;
        RECT 2625.290 16.360 2625.610 16.420 ;
      LAYER via ;
        RECT 1858.500 1685.080 1858.760 1685.340 ;
        RECT 2038.820 1685.080 2039.080 1685.340 ;
        RECT 2039.280 18.400 2039.540 18.660 ;
        RECT 2625.320 16.360 2625.580 16.620 ;
      LAYER met2 ;
        RECT 1858.490 1700.000 1858.770 1704.000 ;
        RECT 1858.560 1685.370 1858.700 1700.000 ;
        RECT 1858.500 1685.050 1858.760 1685.370 ;
        RECT 2038.820 1685.050 2039.080 1685.370 ;
        RECT 2038.880 18.770 2039.020 1685.050 ;
        RECT 2038.880 18.690 2039.480 18.770 ;
        RECT 2038.880 18.630 2039.540 18.690 ;
        RECT 2039.280 18.370 2039.540 18.630 ;
        RECT 2625.320 16.330 2625.580 16.650 ;
        RECT 2625.380 2.400 2625.520 16.330 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1863.530 1686.640 1863.850 1686.700 ;
        RECT 1868.590 1686.640 1868.910 1686.700 ;
        RECT 1863.530 1686.500 1868.910 1686.640 ;
        RECT 1863.530 1686.440 1863.850 1686.500 ;
        RECT 1868.590 1686.440 1868.910 1686.500 ;
        RECT 1868.590 51.920 1868.910 51.980 ;
        RECT 2642.770 51.920 2643.090 51.980 ;
        RECT 1868.590 51.780 2643.090 51.920 ;
        RECT 1868.590 51.720 1868.910 51.780 ;
        RECT 2642.770 51.720 2643.090 51.780 ;
      LAYER via ;
        RECT 1863.560 1686.440 1863.820 1686.700 ;
        RECT 1868.620 1686.440 1868.880 1686.700 ;
        RECT 1868.620 51.720 1868.880 51.980 ;
        RECT 2642.800 51.720 2643.060 51.980 ;
      LAYER met2 ;
        RECT 1863.550 1700.000 1863.830 1704.000 ;
        RECT 1863.620 1686.730 1863.760 1700.000 ;
        RECT 1863.560 1686.410 1863.820 1686.730 ;
        RECT 1868.620 1686.410 1868.880 1686.730 ;
        RECT 1868.680 52.010 1868.820 1686.410 ;
        RECT 1868.620 51.690 1868.880 52.010 ;
        RECT 2642.800 51.690 2643.060 52.010 ;
        RECT 2642.860 3.130 2643.000 51.690 ;
        RECT 2642.860 2.990 2643.460 3.130 ;
        RECT 2643.320 2.400 2643.460 2.990 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 0.300 ;
=======
      LAYER li1 ;
        RECT 1893.965 1684.785 1894.135 1685.975 ;
      LAYER mcon ;
        RECT 1893.965 1685.805 1894.135 1685.975 ;
      LAYER met1 ;
        RECT 1868.130 1685.960 1868.450 1686.020 ;
        RECT 1893.905 1685.960 1894.195 1686.005 ;
        RECT 1868.130 1685.820 1894.195 1685.960 ;
        RECT 1868.130 1685.760 1868.450 1685.820 ;
        RECT 1893.905 1685.775 1894.195 1685.820 ;
        RECT 1893.905 1684.940 1894.195 1684.985 ;
        RECT 2039.250 1684.940 2039.570 1685.000 ;
        RECT 1893.905 1684.800 2039.570 1684.940 ;
        RECT 1893.905 1684.755 1894.195 1684.800 ;
        RECT 2039.250 1684.740 2039.570 1684.800 ;
        RECT 2054.890 20.300 2055.210 20.360 ;
        RECT 2661.170 20.300 2661.490 20.360 ;
        RECT 2054.890 20.160 2661.490 20.300 ;
        RECT 2054.890 20.100 2055.210 20.160 ;
        RECT 2661.170 20.100 2661.490 20.160 ;
      LAYER via ;
        RECT 1868.160 1685.760 1868.420 1686.020 ;
        RECT 2039.280 1684.740 2039.540 1685.000 ;
        RECT 2054.920 20.100 2055.180 20.360 ;
        RECT 2661.200 20.100 2661.460 20.360 ;
      LAYER met2 ;
        RECT 1868.150 1700.000 1868.430 1704.000 ;
        RECT 1868.220 1686.050 1868.360 1700.000 ;
        RECT 1868.160 1685.730 1868.420 1686.050 ;
        RECT 2039.280 1684.710 2039.540 1685.030 ;
        RECT 2039.340 20.925 2039.480 1684.710 ;
        RECT 2039.270 20.555 2039.550 20.925 ;
        RECT 2054.910 20.555 2055.190 20.925 ;
        RECT 2054.980 20.390 2055.120 20.555 ;
        RECT 2054.920 20.070 2055.180 20.390 ;
        RECT 2661.200 20.070 2661.460 20.390 ;
        RECT 2661.260 2.400 2661.400 20.070 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
      LAYER via2 ;
        RECT 2039.270 20.600 2039.550 20.880 ;
        RECT 2054.910 20.600 2055.190 20.880 ;
      LAYER met3 ;
        RECT 2039.245 20.890 2039.575 20.905 ;
        RECT 2054.885 20.890 2055.215 20.905 ;
        RECT 2039.245 20.590 2055.215 20.890 ;
        RECT 2039.245 20.575 2039.575 20.590 ;
        RECT 2054.885 20.575 2055.215 20.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1874.110 1683.580 1874.430 1683.640 ;
        RECT 1876.410 1683.580 1876.730 1683.640 ;
        RECT 1874.110 1683.440 1876.730 1683.580 ;
        RECT 1874.110 1683.380 1874.430 1683.440 ;
        RECT 1876.410 1683.380 1876.730 1683.440 ;
        RECT 1876.410 17.240 1876.730 17.300 ;
        RECT 2678.650 17.240 2678.970 17.300 ;
        RECT 1876.410 17.100 2678.970 17.240 ;
        RECT 1876.410 17.040 1876.730 17.100 ;
        RECT 2678.650 17.040 2678.970 17.100 ;
      LAYER via ;
        RECT 1874.140 1683.380 1874.400 1683.640 ;
        RECT 1876.440 1683.380 1876.700 1683.640 ;
        RECT 1876.440 17.040 1876.700 17.300 ;
        RECT 2678.680 17.040 2678.940 17.300 ;
      LAYER met2 ;
        RECT 1873.210 1700.410 1873.490 1704.000 ;
        RECT 1873.210 1700.270 1874.340 1700.410 ;
        RECT 1873.210 1700.000 1873.490 1700.270 ;
        RECT 1874.200 1683.670 1874.340 1700.270 ;
        RECT 1874.140 1683.350 1874.400 1683.670 ;
        RECT 1876.440 1683.350 1876.700 1683.670 ;
        RECT 1876.500 17.330 1876.640 1683.350 ;
        RECT 1876.440 17.010 1876.700 17.330 ;
        RECT 2678.680 17.010 2678.940 17.330 ;
        RECT 2678.740 2.400 2678.880 17.010 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 0.300 ;
=======
      LAYER li1 ;
        RECT 1939.045 1685.465 1939.215 1690.735 ;
      LAYER mcon ;
        RECT 1939.045 1690.565 1939.215 1690.735 ;
      LAYER met1 ;
        RECT 1879.170 1690.720 1879.490 1690.780 ;
        RECT 1938.985 1690.720 1939.275 1690.765 ;
        RECT 1879.170 1690.580 1939.275 1690.720 ;
        RECT 1879.170 1690.520 1879.490 1690.580 ;
        RECT 1938.985 1690.535 1939.275 1690.580 ;
        RECT 1938.985 1685.620 1939.275 1685.665 ;
        RECT 2073.290 1685.620 2073.610 1685.680 ;
        RECT 1938.985 1685.480 2073.610 1685.620 ;
        RECT 1938.985 1685.435 1939.275 1685.480 ;
        RECT 2073.290 1685.420 2073.610 1685.480 ;
      LAYER via ;
        RECT 1879.200 1690.520 1879.460 1690.780 ;
        RECT 2073.320 1685.420 2073.580 1685.680 ;
      LAYER met2 ;
        RECT 1877.810 1700.410 1878.090 1704.000 ;
        RECT 1877.810 1700.270 1879.400 1700.410 ;
        RECT 1877.810 1700.000 1878.090 1700.270 ;
        RECT 1879.260 1690.810 1879.400 1700.270 ;
        RECT 1879.200 1690.490 1879.460 1690.810 ;
        RECT 2073.320 1685.390 2073.580 1685.710 ;
        RECT 2073.380 20.245 2073.520 1685.390 ;
        RECT 2073.310 19.875 2073.590 20.245 ;
        RECT 2696.610 19.875 2696.890 20.245 ;
        RECT 2696.680 2.400 2696.820 19.875 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
      LAYER via2 ;
        RECT 2073.310 19.920 2073.590 20.200 ;
        RECT 2696.610 19.920 2696.890 20.200 ;
      LAYER met3 ;
        RECT 2073.285 20.210 2073.615 20.225 ;
        RECT 2696.585 20.210 2696.915 20.225 ;
        RECT 2073.285 19.910 2696.915 20.210 ;
        RECT 2073.285 19.895 2073.615 19.910 ;
        RECT 2696.585 19.895 2696.915 19.910 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 0.300 ;
=======
      LAYER met1 ;
        RECT 1883.310 1608.920 1883.630 1609.180 ;
        RECT 1883.400 1608.160 1883.540 1608.920 ;
        RECT 1883.310 1607.900 1883.630 1608.160 ;
      LAYER via ;
        RECT 1883.340 1608.920 1883.600 1609.180 ;
        RECT 1883.340 1607.900 1883.600 1608.160 ;
      LAYER met2 ;
        RECT 1882.870 1700.410 1883.150 1704.000 ;
        RECT 1882.870 1700.270 1883.540 1700.410 ;
        RECT 1882.870 1700.000 1883.150 1700.270 ;
        RECT 1883.400 1609.210 1883.540 1700.270 ;
        RECT 1883.340 1608.890 1883.600 1609.210 ;
        RECT 1883.340 1607.870 1883.600 1608.190 ;
        RECT 1883.400 18.885 1883.540 1607.870 ;
        RECT 1883.330 18.515 1883.610 18.885 ;
        RECT 2714.550 18.515 2714.830 18.885 ;
        RECT 2714.620 2.400 2714.760 18.515 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
      LAYER via2 ;
        RECT 1883.330 18.560 1883.610 18.840 ;
        RECT 2714.550 18.560 2714.830 18.840 ;
      LAYER met3 ;
        RECT 1883.305 18.850 1883.635 18.865 ;
        RECT 2714.525 18.850 2714.855 18.865 ;
        RECT 1883.305 18.550 2714.855 18.850 ;
        RECT 1883.305 18.535 1883.635 18.550 ;
        RECT 2714.525 18.535 2714.855 18.550 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1897.570 1686.640 1897.890 1686.700 ;
        RECT 2121.590 1686.640 2121.910 1686.700 ;
        RECT 1897.570 1686.500 2121.910 1686.640 ;
        RECT 1897.570 1686.440 1897.890 1686.500 ;
        RECT 2121.590 1686.440 2121.910 1686.500 ;
        RECT 2121.590 20.640 2121.910 20.700 ;
        RECT 2732.470 20.640 2732.790 20.700 ;
        RECT 2121.590 20.500 2732.790 20.640 ;
        RECT 2121.590 20.440 2121.910 20.500 ;
        RECT 2732.470 20.440 2732.790 20.500 ;
      LAYER via ;
        RECT 1897.600 1686.440 1897.860 1686.700 ;
        RECT 2121.620 1686.440 2121.880 1686.700 ;
        RECT 2121.620 20.440 2121.880 20.700 ;
        RECT 2732.500 20.440 2732.760 20.700 ;
      LAYER met2 ;
        RECT 1887.470 1700.000 1887.750 1704.000 ;
        RECT 1887.540 1686.925 1887.680 1700.000 ;
        RECT 1887.470 1686.555 1887.750 1686.925 ;
        RECT 1897.590 1686.555 1897.870 1686.925 ;
        RECT 1897.600 1686.410 1897.860 1686.555 ;
        RECT 2121.620 1686.410 2121.880 1686.730 ;
        RECT 2121.680 20.730 2121.820 1686.410 ;
        RECT 2121.620 20.410 2121.880 20.730 ;
        RECT 2732.500 20.410 2732.760 20.730 ;
        RECT 2732.560 2.400 2732.700 20.410 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
      LAYER via2 ;
        RECT 1887.470 1686.600 1887.750 1686.880 ;
        RECT 1897.590 1686.600 1897.870 1686.880 ;
      LAYER met3 ;
        RECT 1887.445 1686.890 1887.775 1686.905 ;
        RECT 1897.565 1686.890 1897.895 1686.905 ;
        RECT 1887.445 1686.590 1897.895 1686.890 ;
        RECT 1887.445 1686.575 1887.775 1686.590 ;
        RECT 1897.565 1686.575 1897.895 1686.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1893.430 1700.920 1893.750 1700.980 ;
        RECT 1895.270 1700.920 1895.590 1700.980 ;
        RECT 1893.430 1700.780 1895.590 1700.920 ;
        RECT 1893.430 1700.720 1893.750 1700.780 ;
        RECT 1895.270 1700.720 1895.590 1700.780 ;
        RECT 1895.730 51.580 1896.050 51.640 ;
        RECT 2746.270 51.580 2746.590 51.640 ;
        RECT 1895.730 51.440 2746.590 51.580 ;
        RECT 1895.730 51.380 1896.050 51.440 ;
        RECT 2746.270 51.380 2746.590 51.440 ;
        RECT 2746.270 2.960 2746.590 3.020 ;
        RECT 2750.410 2.960 2750.730 3.020 ;
        RECT 2746.270 2.820 2750.730 2.960 ;
        RECT 2746.270 2.760 2746.590 2.820 ;
        RECT 2750.410 2.760 2750.730 2.820 ;
      LAYER via ;
        RECT 1893.460 1700.720 1893.720 1700.980 ;
        RECT 1895.300 1700.720 1895.560 1700.980 ;
        RECT 1895.760 51.380 1896.020 51.640 ;
        RECT 2746.300 51.380 2746.560 51.640 ;
        RECT 2746.300 2.760 2746.560 3.020 ;
        RECT 2750.440 2.760 2750.700 3.020 ;
      LAYER met2 ;
        RECT 1892.530 1701.090 1892.810 1704.000 ;
        RECT 1892.530 1701.010 1893.660 1701.090 ;
        RECT 1892.530 1700.950 1893.720 1701.010 ;
        RECT 1892.530 1700.000 1892.810 1700.950 ;
        RECT 1893.460 1700.690 1893.720 1700.950 ;
        RECT 1895.300 1700.690 1895.560 1701.010 ;
        RECT 1895.360 1686.130 1895.500 1700.690 ;
        RECT 1895.360 1685.990 1895.960 1686.130 ;
        RECT 1895.820 51.670 1895.960 1685.990 ;
        RECT 1895.760 51.350 1896.020 51.670 ;
        RECT 2746.300 51.350 2746.560 51.670 ;
        RECT 2746.360 3.050 2746.500 51.350 ;
        RECT 2746.300 2.730 2746.560 3.050 ;
        RECT 2750.440 2.730 2750.700 3.050 ;
        RECT 2750.500 2.400 2750.640 2.730 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 0.300 ;
=======
      LAYER met1 ;
        RECT 2087.090 1685.960 2087.410 1686.020 ;
        RECT 1899.040 1685.820 2087.410 1685.960 ;
        RECT 1897.110 1685.620 1897.430 1685.680 ;
        RECT 1899.040 1685.620 1899.180 1685.820 ;
        RECT 2087.090 1685.760 2087.410 1685.820 ;
        RECT 1897.110 1685.480 1899.180 1685.620 ;
        RECT 1897.110 1685.420 1897.430 1685.480 ;
        RECT 2767.890 18.940 2768.210 19.000 ;
        RECT 2090.400 18.800 2768.210 18.940 ;
        RECT 2088.010 18.600 2088.330 18.660 ;
        RECT 2090.400 18.600 2090.540 18.800 ;
        RECT 2767.890 18.740 2768.210 18.800 ;
        RECT 2088.010 18.460 2090.540 18.600 ;
        RECT 2088.010 18.400 2088.330 18.460 ;
      LAYER via ;
        RECT 1897.140 1685.420 1897.400 1685.680 ;
        RECT 2087.120 1685.760 2087.380 1686.020 ;
        RECT 2088.040 18.400 2088.300 18.660 ;
        RECT 2767.920 18.740 2768.180 19.000 ;
      LAYER met2 ;
        RECT 1897.130 1700.000 1897.410 1704.000 ;
        RECT 1897.200 1685.710 1897.340 1700.000 ;
        RECT 2087.120 1685.730 2087.380 1686.050 ;
        RECT 1897.140 1685.390 1897.400 1685.710 ;
        RECT 2087.180 18.090 2087.320 1685.730 ;
        RECT 2767.920 18.710 2768.180 19.030 ;
        RECT 2088.040 18.370 2088.300 18.690 ;
        RECT 2088.100 18.090 2088.240 18.370 ;
        RECT 2087.180 17.950 2088.240 18.090 ;
        RECT 2767.980 2.400 2768.120 18.710 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1374.090 1678.140 1374.410 1678.200 ;
        RECT 1375.470 1678.140 1375.790 1678.200 ;
        RECT 1374.090 1678.000 1375.790 1678.140 ;
        RECT 1374.090 1677.940 1374.410 1678.000 ;
        RECT 1375.470 1677.940 1375.790 1678.000 ;
        RECT 840.950 37.640 841.270 37.700 ;
        RECT 1374.090 37.640 1374.410 37.700 ;
        RECT 840.950 37.500 1374.410 37.640 ;
        RECT 840.950 37.440 841.270 37.500 ;
        RECT 1374.090 37.440 1374.410 37.500 ;
      LAYER via ;
        RECT 1374.120 1677.940 1374.380 1678.200 ;
        RECT 1375.500 1677.940 1375.760 1678.200 ;
        RECT 840.980 37.440 841.240 37.700 ;
        RECT 1374.120 37.440 1374.380 37.700 ;
      LAYER met2 ;
        RECT 1376.870 1700.410 1377.150 1704.000 ;
        RECT 1375.560 1700.270 1377.150 1700.410 ;
        RECT 1375.560 1678.230 1375.700 1700.270 ;
        RECT 1376.870 1700.000 1377.150 1700.270 ;
        RECT 1374.120 1677.910 1374.380 1678.230 ;
        RECT 1375.500 1677.910 1375.760 1678.230 ;
        RECT 1374.180 37.730 1374.320 1677.910 ;
        RECT 840.980 37.410 841.240 37.730 ;
        RECT 1374.120 37.410 1374.380 37.730 ;
        RECT 841.040 2.400 841.180 37.410 ;
        RECT 840.830 -4.800 841.390 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1898.030 1684.260 1898.350 1684.320 ;
        RECT 1902.170 1684.260 1902.490 1684.320 ;
        RECT 1898.030 1684.120 1902.490 1684.260 ;
        RECT 1898.030 1684.060 1898.350 1684.120 ;
        RECT 1902.170 1684.060 1902.490 1684.120 ;
        RECT 1898.030 1632.240 1898.350 1632.300 ;
        RECT 1904.010 1632.240 1904.330 1632.300 ;
        RECT 1898.030 1632.100 1904.330 1632.240 ;
        RECT 1898.030 1632.040 1898.350 1632.100 ;
        RECT 1904.010 1632.040 1904.330 1632.100 ;
      LAYER via ;
        RECT 1898.060 1684.060 1898.320 1684.320 ;
        RECT 1902.200 1684.060 1902.460 1684.320 ;
        RECT 1898.060 1632.040 1898.320 1632.300 ;
        RECT 1904.040 1632.040 1904.300 1632.300 ;
      LAYER met2 ;
        RECT 1902.190 1700.000 1902.470 1704.000 ;
        RECT 1902.260 1684.350 1902.400 1700.000 ;
        RECT 1898.060 1684.030 1898.320 1684.350 ;
        RECT 1902.200 1684.030 1902.460 1684.350 ;
        RECT 1898.120 1632.330 1898.260 1684.030 ;
        RECT 1898.060 1632.010 1898.320 1632.330 ;
        RECT 1904.040 1632.010 1904.300 1632.330 ;
        RECT 1904.100 18.205 1904.240 1632.010 ;
        RECT 1904.030 17.835 1904.310 18.205 ;
        RECT 2785.850 17.835 2786.130 18.205 ;
        RECT 2785.920 2.400 2786.060 17.835 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
      LAYER via2 ;
        RECT 1904.030 17.880 1904.310 18.160 ;
        RECT 2785.850 17.880 2786.130 18.160 ;
      LAYER met3 ;
        RECT 1904.005 18.170 1904.335 18.185 ;
        RECT 2785.825 18.170 2786.155 18.185 ;
        RECT 1904.005 17.870 2786.155 18.170 ;
        RECT 1904.005 17.855 1904.335 17.870 ;
        RECT 2785.825 17.855 2786.155 17.870 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 0.300 ;
=======
      LAYER met1 ;
        RECT 2142.290 19.620 2142.610 19.680 ;
        RECT 2803.770 19.620 2804.090 19.680 ;
        RECT 2142.290 19.480 2804.090 19.620 ;
        RECT 2142.290 19.420 2142.610 19.480 ;
        RECT 2803.770 19.420 2804.090 19.480 ;
      LAYER via ;
        RECT 2142.320 19.420 2142.580 19.680 ;
        RECT 2803.800 19.420 2804.060 19.680 ;
      LAYER met2 ;
        RECT 1906.790 1700.000 1907.070 1704.000 ;
        RECT 1906.860 1688.965 1907.000 1700.000 ;
        RECT 1906.790 1688.595 1907.070 1688.965 ;
        RECT 2142.310 1688.595 2142.590 1688.965 ;
        RECT 2142.380 19.710 2142.520 1688.595 ;
        RECT 2142.320 19.390 2142.580 19.710 ;
        RECT 2803.800 19.390 2804.060 19.710 ;
        RECT 2803.860 2.400 2804.000 19.390 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
      LAYER via2 ;
        RECT 1906.790 1688.640 1907.070 1688.920 ;
        RECT 2142.310 1688.640 2142.590 1688.920 ;
      LAYER met3 ;
        RECT 1906.765 1688.930 1907.095 1688.945 ;
        RECT 2142.285 1688.930 2142.615 1688.945 ;
        RECT 1906.765 1688.630 2142.615 1688.930 ;
        RECT 1906.765 1688.615 1907.095 1688.630 ;
        RECT 2142.285 1688.615 2142.615 1688.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 0.300 ;
=======
      LAYER met1 ;
        RECT 1911.830 1686.300 1912.150 1686.360 ;
        RECT 1916.890 1686.300 1917.210 1686.360 ;
        RECT 1911.830 1686.160 1917.210 1686.300 ;
        RECT 1911.830 1686.100 1912.150 1686.160 ;
        RECT 1916.890 1686.100 1917.210 1686.160 ;
      LAYER via ;
        RECT 1911.860 1686.100 1912.120 1686.360 ;
        RECT 1916.920 1686.100 1917.180 1686.360 ;
      LAYER met2 ;
        RECT 1911.850 1700.000 1912.130 1704.000 ;
        RECT 1911.920 1686.390 1912.060 1700.000 ;
        RECT 1911.860 1686.070 1912.120 1686.390 ;
        RECT 1916.920 1686.070 1917.180 1686.390 ;
        RECT 1916.980 44.725 1917.120 1686.070 ;
        RECT 1916.910 44.355 1917.190 44.725 ;
        RECT 2821.730 44.355 2822.010 44.725 ;
        RECT 2821.800 2.400 2821.940 44.355 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
      LAYER via2 ;
        RECT 1916.910 44.400 1917.190 44.680 ;
        RECT 2821.730 44.400 2822.010 44.680 ;
      LAYER met3 ;
        RECT 1916.885 44.690 1917.215 44.705 ;
        RECT 2821.705 44.690 2822.035 44.705 ;
        RECT 1916.885 44.390 2822.035 44.690 ;
        RECT 1916.885 44.375 1917.215 44.390 ;
        RECT 2821.705 44.375 2822.035 44.390 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 0.300 ;
=======
      LAYER li1 ;
        RECT 2183.765 17.765 2183.935 18.615 ;
      LAYER mcon ;
        RECT 2183.765 18.445 2183.935 18.615 ;
      LAYER met1 ;
        RECT 2183.705 18.600 2183.995 18.645 ;
        RECT 2839.190 18.600 2839.510 18.660 ;
        RECT 2183.705 18.460 2839.510 18.600 ;
        RECT 2183.705 18.415 2183.995 18.460 ;
        RECT 2839.190 18.400 2839.510 18.460 ;
        RECT 2149.190 17.920 2149.510 17.980 ;
        RECT 2183.705 17.920 2183.995 17.965 ;
        RECT 2149.190 17.780 2183.995 17.920 ;
        RECT 2149.190 17.720 2149.510 17.780 ;
        RECT 2183.705 17.735 2183.995 17.780 ;
      LAYER via ;
        RECT 2839.220 18.400 2839.480 18.660 ;
        RECT 2149.220 17.720 2149.480 17.980 ;
      LAYER met2 ;
        RECT 1916.450 1700.000 1916.730 1704.000 ;
        RECT 1916.520 1688.285 1916.660 1700.000 ;
        RECT 1916.450 1687.915 1916.730 1688.285 ;
        RECT 2149.210 1687.915 2149.490 1688.285 ;
        RECT 2149.280 18.010 2149.420 1687.915 ;
        RECT 2839.220 18.370 2839.480 18.690 ;
        RECT 2149.220 17.690 2149.480 18.010 ;
        RECT 2839.280 2.400 2839.420 18.370 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
      LAYER via2 ;
        RECT 1916.450 1687.960 1916.730 1688.240 ;
        RECT 2149.210 1687.960 2149.490 1688.240 ;
      LAYER met3 ;
        RECT 1916.425 1688.250 1916.755 1688.265 ;
        RECT 2149.185 1688.250 2149.515 1688.265 ;
        RECT 1916.425 1687.950 2149.515 1688.250 ;
        RECT 1916.425 1687.935 1916.755 1687.950 ;
        RECT 2149.185 1687.935 2149.515 1687.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1920.110 1632.240 1920.430 1632.300 ;
        RECT 1924.710 1632.240 1925.030 1632.300 ;
        RECT 1920.110 1632.100 1925.030 1632.240 ;
        RECT 1920.110 1632.040 1920.430 1632.100 ;
        RECT 1924.710 1632.040 1925.030 1632.100 ;
      LAYER via ;
        RECT 1920.140 1632.040 1920.400 1632.300 ;
        RECT 1924.740 1632.040 1925.000 1632.300 ;
      LAYER met2 ;
        RECT 1921.510 1700.410 1921.790 1704.000 ;
        RECT 1920.200 1700.270 1921.790 1700.410 ;
        RECT 1920.200 1632.330 1920.340 1700.270 ;
        RECT 1921.510 1700.000 1921.790 1700.270 ;
        RECT 1920.140 1632.010 1920.400 1632.330 ;
        RECT 1924.740 1632.010 1925.000 1632.330 ;
        RECT 1924.800 17.525 1924.940 1632.010 ;
        RECT 1924.730 17.155 1925.010 17.525 ;
        RECT 2857.150 17.155 2857.430 17.525 ;
        RECT 2857.220 2.400 2857.360 17.155 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
      LAYER via2 ;
        RECT 1924.730 17.200 1925.010 17.480 ;
        RECT 2857.150 17.200 2857.430 17.480 ;
      LAYER met3 ;
        RECT 1924.705 17.490 1925.035 17.505 ;
        RECT 2857.125 17.490 2857.455 17.505 ;
        RECT 1924.705 17.190 2857.455 17.490 ;
        RECT 1924.705 17.175 1925.035 17.190 ;
        RECT 2857.125 17.175 2857.455 17.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 0.300 ;
=======
      LAYER li1 ;
        RECT 2183.305 18.785 2184.395 18.955 ;
        RECT 2183.305 18.445 2183.475 18.785 ;
        RECT 2184.225 17.765 2184.395 18.785 ;
      LAYER met1 ;
        RECT 2180.010 18.600 2180.330 18.660 ;
        RECT 2183.245 18.600 2183.535 18.645 ;
        RECT 2180.010 18.460 2183.535 18.600 ;
        RECT 2180.010 18.400 2180.330 18.460 ;
        RECT 2183.245 18.415 2183.535 18.460 ;
        RECT 2184.165 17.920 2184.455 17.965 ;
        RECT 2875.070 17.920 2875.390 17.980 ;
        RECT 2184.165 17.780 2875.390 17.920 ;
        RECT 2184.165 17.735 2184.455 17.780 ;
        RECT 2875.070 17.720 2875.390 17.780 ;
      LAYER via ;
        RECT 2180.040 18.400 2180.300 18.660 ;
        RECT 2875.100 17.720 2875.360 17.980 ;
      LAYER met2 ;
        RECT 1926.110 1700.000 1926.390 1704.000 ;
        RECT 1926.180 1687.605 1926.320 1700.000 ;
        RECT 1926.110 1687.235 1926.390 1687.605 ;
        RECT 2176.810 1687.235 2177.090 1687.605 ;
        RECT 2176.880 26.250 2177.020 1687.235 ;
        RECT 2176.880 26.110 2180.240 26.250 ;
        RECT 2180.100 18.690 2180.240 26.110 ;
        RECT 2180.040 18.370 2180.300 18.690 ;
        RECT 2875.100 17.690 2875.360 18.010 ;
        RECT 2875.160 2.400 2875.300 17.690 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
      LAYER via2 ;
        RECT 1926.110 1687.280 1926.390 1687.560 ;
        RECT 2176.810 1687.280 2177.090 1687.560 ;
      LAYER met3 ;
        RECT 1926.085 1687.570 1926.415 1687.585 ;
        RECT 2176.785 1687.570 2177.115 1687.585 ;
        RECT 1926.085 1687.270 2177.115 1687.570 ;
        RECT 1926.085 1687.255 1926.415 1687.270 ;
        RECT 2176.785 1687.255 2177.115 1687.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1925.170 1685.620 1925.490 1685.680 ;
        RECT 1931.150 1685.620 1931.470 1685.680 ;
        RECT 1925.170 1685.480 1931.470 1685.620 ;
        RECT 1925.170 1685.420 1925.490 1685.480 ;
        RECT 1931.150 1685.420 1931.470 1685.480 ;
        RECT 1925.170 1631.900 1925.490 1631.960 ;
        RECT 1931.610 1631.900 1931.930 1631.960 ;
        RECT 1925.170 1631.760 1931.930 1631.900 ;
        RECT 1925.170 1631.700 1925.490 1631.760 ;
        RECT 1931.610 1631.700 1931.930 1631.760 ;
      LAYER via ;
        RECT 1925.200 1685.420 1925.460 1685.680 ;
        RECT 1931.180 1685.420 1931.440 1685.680 ;
        RECT 1925.200 1631.700 1925.460 1631.960 ;
        RECT 1931.640 1631.700 1931.900 1631.960 ;
      LAYER met2 ;
        RECT 1931.170 1700.000 1931.450 1704.000 ;
        RECT 1931.240 1685.710 1931.380 1700.000 ;
        RECT 1925.200 1685.390 1925.460 1685.710 ;
        RECT 1931.180 1685.390 1931.440 1685.710 ;
        RECT 1925.260 1631.990 1925.400 1685.390 ;
        RECT 1925.200 1631.670 1925.460 1631.990 ;
        RECT 1931.640 1631.670 1931.900 1631.990 ;
        RECT 1931.700 16.845 1931.840 1631.670 ;
        RECT 1931.630 16.475 1931.910 16.845 ;
        RECT 2893.030 16.475 2893.310 16.845 ;
        RECT 2893.100 2.400 2893.240 16.475 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 1931.630 16.520 1931.910 16.800 ;
        RECT 2893.030 16.520 2893.310 16.800 ;
      LAYER met3 ;
        RECT 1931.605 16.810 1931.935 16.825 ;
        RECT 2893.005 16.810 2893.335 16.825 ;
        RECT 1931.605 16.510 2893.335 16.810 ;
        RECT 1931.605 16.495 1931.935 16.510 ;
        RECT 2893.005 16.495 2893.335 16.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 0.300 ;
=======
      LAYER met1 ;
        RECT 2218.190 18.260 2218.510 18.320 ;
        RECT 2910.950 18.260 2911.270 18.320 ;
        RECT 2218.190 18.120 2911.270 18.260 ;
        RECT 2218.190 18.060 2218.510 18.120 ;
        RECT 2910.950 18.060 2911.270 18.120 ;
      LAYER via ;
        RECT 2218.220 18.060 2218.480 18.320 ;
        RECT 2910.980 18.060 2911.240 18.320 ;
      LAYER met2 ;
        RECT 1935.770 1700.000 1936.050 1704.000 ;
        RECT 1935.840 1686.925 1935.980 1700.000 ;
        RECT 1935.770 1686.555 1936.050 1686.925 ;
        RECT 2218.210 1686.555 2218.490 1686.925 ;
        RECT 2218.280 18.350 2218.420 1686.555 ;
        RECT 2218.220 18.030 2218.480 18.350 ;
        RECT 2910.980 18.030 2911.240 18.350 ;
        RECT 2911.040 2.400 2911.180 18.030 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 1935.770 1686.600 1936.050 1686.880 ;
        RECT 2218.210 1686.600 2218.490 1686.880 ;
      LAYER met3 ;
        RECT 1935.745 1686.890 1936.075 1686.905 ;
        RECT 2218.185 1686.890 2218.515 1686.905 ;
        RECT 1935.745 1686.590 2218.515 1686.890 ;
        RECT 1935.745 1686.575 1936.075 1686.590 ;
        RECT 2218.185 1686.575 2218.515 1686.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 0.300 ;
=======
      LAYER met1 ;
        RECT 858.890 37.300 859.210 37.360 ;
        RECT 1381.910 37.300 1382.230 37.360 ;
        RECT 858.890 37.160 1382.230 37.300 ;
        RECT 858.890 37.100 859.210 37.160 ;
        RECT 1381.910 37.100 1382.230 37.160 ;
      LAYER via ;
        RECT 858.920 37.100 859.180 37.360 ;
        RECT 1381.940 37.100 1382.200 37.360 ;
      LAYER met2 ;
        RECT 1381.470 1700.410 1381.750 1704.000 ;
        RECT 1381.470 1700.270 1382.140 1700.410 ;
        RECT 1381.470 1700.000 1381.750 1700.270 ;
        RECT 1382.000 37.390 1382.140 1700.270 ;
        RECT 858.920 37.070 859.180 37.390 ;
        RECT 1381.940 37.070 1382.200 37.390 ;
        RECT 858.980 2.400 859.120 37.070 ;
        RECT 858.770 -4.800 859.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 0.300 ;
=======
      LAYER li1 ;
        RECT 1383.365 593.045 1383.535 627.895 ;
        RECT 1382.905 469.285 1383.075 496.995 ;
        RECT 1383.365 372.725 1383.535 420.835 ;
        RECT 1382.905 179.605 1383.075 227.715 ;
      LAYER mcon ;
        RECT 1383.365 627.725 1383.535 627.895 ;
        RECT 1382.905 496.825 1383.075 496.995 ;
        RECT 1383.365 420.665 1383.535 420.835 ;
        RECT 1382.905 227.545 1383.075 227.715 ;
      LAYER met1 ;
        RECT 1382.830 1678.480 1383.150 1678.540 ;
        RECT 1386.050 1678.480 1386.370 1678.540 ;
        RECT 1382.830 1678.340 1386.370 1678.480 ;
        RECT 1382.830 1678.280 1383.150 1678.340 ;
        RECT 1386.050 1678.280 1386.370 1678.340 ;
        RECT 1382.830 1607.900 1383.150 1608.160 ;
        RECT 1382.920 1607.420 1383.060 1607.900 ;
        RECT 1383.290 1607.420 1383.610 1607.480 ;
        RECT 1382.920 1607.280 1383.610 1607.420 ;
        RECT 1383.290 1607.220 1383.610 1607.280 ;
        RECT 1383.290 1593.620 1383.610 1593.880 ;
        RECT 1383.380 1593.200 1383.520 1593.620 ;
        RECT 1383.290 1592.940 1383.610 1593.200 ;
        RECT 1383.290 1159.300 1383.610 1159.360 ;
        RECT 1384.210 1159.300 1384.530 1159.360 ;
        RECT 1383.290 1159.160 1384.530 1159.300 ;
        RECT 1383.290 1159.100 1383.610 1159.160 ;
        RECT 1384.210 1159.100 1384.530 1159.160 ;
        RECT 1383.290 966.180 1383.610 966.240 ;
        RECT 1384.210 966.180 1384.530 966.240 ;
        RECT 1383.290 966.040 1384.530 966.180 ;
        RECT 1383.290 965.980 1383.610 966.040 ;
        RECT 1384.210 965.980 1384.530 966.040 ;
        RECT 1383.290 627.880 1383.610 627.940 ;
        RECT 1383.095 627.740 1383.610 627.880 ;
        RECT 1383.290 627.680 1383.610 627.740 ;
        RECT 1383.290 593.200 1383.610 593.260 ;
        RECT 1383.095 593.060 1383.610 593.200 ;
        RECT 1383.290 593.000 1383.610 593.060 ;
        RECT 1382.845 496.980 1383.135 497.025 ;
        RECT 1383.290 496.980 1383.610 497.040 ;
        RECT 1382.845 496.840 1383.610 496.980 ;
        RECT 1382.845 496.795 1383.135 496.840 ;
        RECT 1383.290 496.780 1383.610 496.840 ;
        RECT 1382.830 469.440 1383.150 469.500 ;
        RECT 1382.635 469.300 1383.150 469.440 ;
        RECT 1382.830 469.240 1383.150 469.300 ;
        RECT 1382.830 427.960 1383.150 428.020 ;
        RECT 1383.290 427.960 1383.610 428.020 ;
        RECT 1382.830 427.820 1383.610 427.960 ;
        RECT 1382.830 427.760 1383.150 427.820 ;
        RECT 1383.290 427.760 1383.610 427.820 ;
        RECT 1383.290 420.820 1383.610 420.880 ;
        RECT 1383.095 420.680 1383.610 420.820 ;
        RECT 1383.290 420.620 1383.610 420.680 ;
        RECT 1383.290 372.880 1383.610 372.940 ;
        RECT 1383.095 372.740 1383.610 372.880 ;
        RECT 1383.290 372.680 1383.610 372.740 ;
        RECT 1382.845 227.700 1383.135 227.745 ;
        RECT 1383.750 227.700 1384.070 227.760 ;
        RECT 1382.845 227.560 1384.070 227.700 ;
        RECT 1382.845 227.515 1383.135 227.560 ;
        RECT 1383.750 227.500 1384.070 227.560 ;
        RECT 1382.830 179.760 1383.150 179.820 ;
        RECT 1382.635 179.620 1383.150 179.760 ;
        RECT 1382.830 179.560 1383.150 179.620 ;
        RECT 876.830 36.960 877.150 37.020 ;
        RECT 1383.290 36.960 1383.610 37.020 ;
        RECT 876.830 36.820 1383.610 36.960 ;
        RECT 876.830 36.760 877.150 36.820 ;
        RECT 1383.290 36.760 1383.610 36.820 ;
      LAYER via ;
        RECT 1382.860 1678.280 1383.120 1678.540 ;
        RECT 1386.080 1678.280 1386.340 1678.540 ;
        RECT 1382.860 1607.900 1383.120 1608.160 ;
        RECT 1383.320 1607.220 1383.580 1607.480 ;
        RECT 1383.320 1593.620 1383.580 1593.880 ;
        RECT 1383.320 1592.940 1383.580 1593.200 ;
        RECT 1383.320 1159.100 1383.580 1159.360 ;
        RECT 1384.240 1159.100 1384.500 1159.360 ;
        RECT 1383.320 965.980 1383.580 966.240 ;
        RECT 1384.240 965.980 1384.500 966.240 ;
        RECT 1383.320 627.680 1383.580 627.940 ;
        RECT 1383.320 593.000 1383.580 593.260 ;
        RECT 1383.320 496.780 1383.580 497.040 ;
        RECT 1382.860 469.240 1383.120 469.500 ;
        RECT 1382.860 427.760 1383.120 428.020 ;
        RECT 1383.320 427.760 1383.580 428.020 ;
        RECT 1383.320 420.620 1383.580 420.880 ;
        RECT 1383.320 372.680 1383.580 372.940 ;
        RECT 1383.780 227.500 1384.040 227.760 ;
        RECT 1382.860 179.560 1383.120 179.820 ;
        RECT 876.860 36.760 877.120 37.020 ;
        RECT 1383.320 36.760 1383.580 37.020 ;
      LAYER met2 ;
        RECT 1386.530 1700.410 1386.810 1704.000 ;
        RECT 1386.140 1700.270 1386.810 1700.410 ;
        RECT 1386.140 1678.570 1386.280 1700.270 ;
        RECT 1386.530 1700.000 1386.810 1700.270 ;
        RECT 1382.860 1678.250 1383.120 1678.570 ;
        RECT 1386.080 1678.250 1386.340 1678.570 ;
        RECT 1382.920 1608.190 1383.060 1678.250 ;
        RECT 1382.860 1607.870 1383.120 1608.190 ;
        RECT 1383.320 1607.190 1383.580 1607.510 ;
        RECT 1383.380 1593.910 1383.520 1607.190 ;
        RECT 1383.320 1593.590 1383.580 1593.910 ;
        RECT 1383.320 1592.910 1383.580 1593.230 ;
        RECT 1383.380 1463.090 1383.520 1592.910 ;
        RECT 1382.920 1462.950 1383.520 1463.090 ;
        RECT 1382.920 1462.410 1383.060 1462.950 ;
        RECT 1382.920 1462.270 1383.520 1462.410 ;
        RECT 1383.380 1366.530 1383.520 1462.270 ;
        RECT 1382.920 1366.390 1383.520 1366.530 ;
        RECT 1382.920 1365.850 1383.060 1366.390 ;
        RECT 1382.920 1365.710 1383.520 1365.850 ;
        RECT 1383.380 1269.970 1383.520 1365.710 ;
        RECT 1382.920 1269.830 1383.520 1269.970 ;
        RECT 1382.920 1269.290 1383.060 1269.830 ;
        RECT 1382.920 1269.150 1383.520 1269.290 ;
        RECT 1383.380 1207.525 1383.520 1269.150 ;
        RECT 1383.310 1207.155 1383.590 1207.525 ;
        RECT 1384.230 1207.155 1384.510 1207.525 ;
        RECT 1384.300 1159.390 1384.440 1207.155 ;
        RECT 1383.320 1159.070 1383.580 1159.390 ;
        RECT 1384.240 1159.070 1384.500 1159.390 ;
        RECT 1383.380 1014.405 1383.520 1159.070 ;
        RECT 1383.310 1014.035 1383.590 1014.405 ;
        RECT 1384.230 1014.035 1384.510 1014.405 ;
        RECT 1384.300 966.270 1384.440 1014.035 ;
        RECT 1383.320 965.950 1383.580 966.270 ;
        RECT 1384.240 965.950 1384.500 966.270 ;
        RECT 1383.380 883.730 1383.520 965.950 ;
        RECT 1382.920 883.590 1383.520 883.730 ;
        RECT 1382.920 883.050 1383.060 883.590 ;
        RECT 1382.920 882.910 1383.520 883.050 ;
        RECT 1383.380 787.170 1383.520 882.910 ;
        RECT 1382.920 787.030 1383.520 787.170 ;
        RECT 1382.920 785.810 1383.060 787.030 ;
        RECT 1382.920 785.670 1383.520 785.810 ;
        RECT 1383.380 627.970 1383.520 785.670 ;
        RECT 1383.320 627.650 1383.580 627.970 ;
        RECT 1383.320 592.970 1383.580 593.290 ;
        RECT 1383.380 497.070 1383.520 592.970 ;
        RECT 1383.320 496.750 1383.580 497.070 ;
        RECT 1382.860 469.210 1383.120 469.530 ;
        RECT 1382.920 428.050 1383.060 469.210 ;
        RECT 1382.860 427.730 1383.120 428.050 ;
        RECT 1383.320 427.730 1383.580 428.050 ;
        RECT 1383.380 420.910 1383.520 427.730 ;
        RECT 1383.320 420.590 1383.580 420.910 ;
        RECT 1383.320 372.650 1383.580 372.970 ;
        RECT 1383.380 235.125 1383.520 372.650 ;
        RECT 1383.310 234.755 1383.590 235.125 ;
        RECT 1383.770 234.075 1384.050 234.445 ;
        RECT 1383.840 227.790 1383.980 234.075 ;
        RECT 1383.780 227.470 1384.040 227.790 ;
        RECT 1382.860 179.530 1383.120 179.850 ;
        RECT 1382.920 144.570 1383.060 179.530 ;
        RECT 1382.920 144.430 1383.520 144.570 ;
        RECT 1383.380 37.050 1383.520 144.430 ;
        RECT 876.860 36.730 877.120 37.050 ;
        RECT 1383.320 36.730 1383.580 37.050 ;
        RECT 876.920 2.400 877.060 36.730 ;
        RECT 876.710 -4.800 877.270 2.400 ;
      LAYER via2 ;
        RECT 1383.310 1207.200 1383.590 1207.480 ;
        RECT 1384.230 1207.200 1384.510 1207.480 ;
        RECT 1383.310 1014.080 1383.590 1014.360 ;
        RECT 1384.230 1014.080 1384.510 1014.360 ;
        RECT 1383.310 234.800 1383.590 235.080 ;
        RECT 1383.770 234.120 1384.050 234.400 ;
      LAYER met3 ;
        RECT 1383.285 1207.490 1383.615 1207.505 ;
        RECT 1384.205 1207.490 1384.535 1207.505 ;
        RECT 1383.285 1207.190 1384.535 1207.490 ;
        RECT 1383.285 1207.175 1383.615 1207.190 ;
        RECT 1384.205 1207.175 1384.535 1207.190 ;
        RECT 1383.285 1014.370 1383.615 1014.385 ;
        RECT 1384.205 1014.370 1384.535 1014.385 ;
        RECT 1383.285 1014.070 1384.535 1014.370 ;
        RECT 1383.285 1014.055 1383.615 1014.070 ;
        RECT 1384.205 1014.055 1384.535 1014.070 ;
        RECT 1383.285 235.090 1383.615 235.105 ;
        RECT 1383.070 234.775 1383.615 235.090 ;
        RECT 1383.070 234.410 1383.370 234.775 ;
        RECT 1383.745 234.410 1384.075 234.425 ;
        RECT 1383.070 234.110 1384.075 234.410 ;
        RECT 1383.745 234.095 1384.075 234.110 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 0.300 ;
=======
      LAYER met1 ;
        RECT 1388.350 1678.140 1388.670 1678.200 ;
        RECT 1390.190 1678.140 1390.510 1678.200 ;
        RECT 1388.350 1678.000 1390.510 1678.140 ;
        RECT 1388.350 1677.940 1388.670 1678.000 ;
        RECT 1390.190 1677.940 1390.510 1678.000 ;
        RECT 894.770 36.620 895.090 36.680 ;
        RECT 1388.350 36.620 1388.670 36.680 ;
        RECT 894.770 36.480 1388.670 36.620 ;
        RECT 894.770 36.420 895.090 36.480 ;
        RECT 1388.350 36.420 1388.670 36.480 ;
      LAYER via ;
        RECT 1388.380 1677.940 1388.640 1678.200 ;
        RECT 1390.220 1677.940 1390.480 1678.200 ;
        RECT 894.800 36.420 895.060 36.680 ;
        RECT 1388.380 36.420 1388.640 36.680 ;
      LAYER met2 ;
        RECT 1391.130 1700.410 1391.410 1704.000 ;
        RECT 1390.280 1700.270 1391.410 1700.410 ;
        RECT 1390.280 1678.230 1390.420 1700.270 ;
        RECT 1391.130 1700.000 1391.410 1700.270 ;
        RECT 1388.380 1677.910 1388.640 1678.230 ;
        RECT 1390.220 1677.910 1390.480 1678.230 ;
        RECT 1388.440 36.710 1388.580 1677.910 ;
        RECT 894.800 36.390 895.060 36.710 ;
        RECT 1388.380 36.390 1388.640 36.710 ;
        RECT 894.860 2.400 895.000 36.390 ;
        RECT 894.650 -4.800 895.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 0.300 ;
=======
      LAYER met1 ;
        RECT 912.710 36.280 913.030 36.340 ;
        RECT 1395.250 36.280 1395.570 36.340 ;
        RECT 912.710 36.140 1395.570 36.280 ;
        RECT 912.710 36.080 913.030 36.140 ;
        RECT 1395.250 36.080 1395.570 36.140 ;
      LAYER via ;
        RECT 912.740 36.080 913.000 36.340 ;
        RECT 1395.280 36.080 1395.540 36.340 ;
      LAYER met2 ;
        RECT 1396.190 1700.410 1396.470 1704.000 ;
        RECT 1395.340 1700.270 1396.470 1700.410 ;
        RECT 1395.340 36.370 1395.480 1700.270 ;
        RECT 1396.190 1700.000 1396.470 1700.270 ;
        RECT 912.740 36.050 913.000 36.370 ;
        RECT 1395.280 36.050 1395.540 36.370 ;
        RECT 912.800 2.400 912.940 36.050 ;
        RECT 912.590 -4.800 913.150 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 0.300 ;
=======
      LAYER met1 ;
        RECT 930.190 35.940 930.510 36.000 ;
        RECT 1401.690 35.940 1402.010 36.000 ;
        RECT 930.190 35.800 1402.010 35.940 ;
        RECT 930.190 35.740 930.510 35.800 ;
        RECT 1401.690 35.740 1402.010 35.800 ;
      LAYER via ;
        RECT 930.220 35.740 930.480 36.000 ;
        RECT 1401.720 35.740 1401.980 36.000 ;
      LAYER met2 ;
        RECT 1400.790 1700.410 1401.070 1704.000 ;
        RECT 1400.790 1700.270 1401.920 1700.410 ;
        RECT 1400.790 1700.000 1401.070 1700.270 ;
        RECT 1401.780 36.030 1401.920 1700.270 ;
        RECT 930.220 35.710 930.480 36.030 ;
        RECT 1401.720 35.710 1401.980 36.030 ;
        RECT 930.280 2.400 930.420 35.710 ;
        RECT 930.070 -4.800 930.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1402.150 1678.140 1402.470 1678.200 ;
        RECT 1404.450 1678.140 1404.770 1678.200 ;
        RECT 1402.150 1678.000 1404.770 1678.140 ;
        RECT 1402.150 1677.940 1402.470 1678.000 ;
        RECT 1404.450 1677.940 1404.770 1678.000 ;
        RECT 948.130 35.600 948.450 35.660 ;
        RECT 1402.150 35.600 1402.470 35.660 ;
        RECT 948.130 35.460 1402.470 35.600 ;
        RECT 948.130 35.400 948.450 35.460 ;
        RECT 1402.150 35.400 1402.470 35.460 ;
      LAYER via ;
        RECT 1402.180 1677.940 1402.440 1678.200 ;
        RECT 1404.480 1677.940 1404.740 1678.200 ;
        RECT 948.160 35.400 948.420 35.660 ;
        RECT 1402.180 35.400 1402.440 35.660 ;
      LAYER met2 ;
        RECT 1405.850 1700.410 1406.130 1704.000 ;
        RECT 1404.540 1700.270 1406.130 1700.410 ;
        RECT 1404.540 1678.230 1404.680 1700.270 ;
        RECT 1405.850 1700.000 1406.130 1700.270 ;
        RECT 1402.180 1677.910 1402.440 1678.230 ;
        RECT 1404.480 1677.910 1404.740 1678.230 ;
        RECT 1402.240 35.690 1402.380 1677.910 ;
        RECT 948.160 35.370 948.420 35.690 ;
        RECT 1402.180 35.370 1402.440 35.690 ;
        RECT 948.220 2.400 948.360 35.370 ;
        RECT 948.010 -4.800 948.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 0.300 ;
=======
      LAYER met1 ;
        RECT 966.070 35.260 966.390 35.320 ;
        RECT 1409.510 35.260 1409.830 35.320 ;
        RECT 966.070 35.120 1409.830 35.260 ;
        RECT 966.070 35.060 966.390 35.120 ;
        RECT 1409.510 35.060 1409.830 35.120 ;
      LAYER via ;
        RECT 966.100 35.060 966.360 35.320 ;
        RECT 1409.540 35.060 1409.800 35.320 ;
      LAYER met2 ;
        RECT 1410.450 1700.410 1410.730 1704.000 ;
        RECT 1409.600 1700.270 1410.730 1700.410 ;
        RECT 1409.600 35.350 1409.740 1700.270 ;
        RECT 1410.450 1700.000 1410.730 1700.270 ;
        RECT 966.100 35.030 966.360 35.350 ;
        RECT 1409.540 35.030 1409.800 35.350 ;
        RECT 966.160 2.400 966.300 35.030 ;
        RECT 965.950 -4.800 966.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 0.300 ;
=======
      LAYER met1 ;
        RECT 984.010 34.920 984.330 34.980 ;
        RECT 1415.490 34.920 1415.810 34.980 ;
        RECT 984.010 34.780 1415.810 34.920 ;
        RECT 984.010 34.720 984.330 34.780 ;
        RECT 1415.490 34.720 1415.810 34.780 ;
      LAYER via ;
        RECT 984.040 34.720 984.300 34.980 ;
        RECT 1415.520 34.720 1415.780 34.980 ;
      LAYER met2 ;
        RECT 1415.510 1700.000 1415.790 1704.000 ;
        RECT 1415.580 35.010 1415.720 1700.000 ;
        RECT 984.040 34.690 984.300 35.010 ;
        RECT 1415.520 34.690 1415.780 35.010 ;
        RECT 984.100 2.400 984.240 34.690 ;
        RECT 983.890 -4.800 984.450 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 0.300 ;
=======
      LAYER met1 ;
        RECT 662.930 39.000 663.250 39.060 ;
        RECT 1326.250 39.000 1326.570 39.060 ;
        RECT 662.930 38.860 1326.570 39.000 ;
        RECT 662.930 38.800 663.250 38.860 ;
        RECT 1326.250 38.800 1326.570 38.860 ;
      LAYER via ;
        RECT 662.960 38.800 663.220 39.060 ;
        RECT 1326.280 38.800 1326.540 39.060 ;
      LAYER met2 ;
        RECT 1328.570 1700.410 1328.850 1704.000 ;
        RECT 1327.720 1700.270 1328.850 1700.410 ;
        RECT 1327.720 1677.970 1327.860 1700.270 ;
        RECT 1328.570 1700.000 1328.850 1700.270 ;
        RECT 1326.340 1677.830 1327.860 1677.970 ;
        RECT 1326.340 39.090 1326.480 1677.830 ;
        RECT 662.960 38.770 663.220 39.090 ;
        RECT 1326.280 38.770 1326.540 39.090 ;
        RECT 663.020 2.400 663.160 38.770 ;
        RECT 662.810 -4.800 663.370 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 0.300 ;
=======
      LAYER li1 ;
        RECT 1416.025 1442.025 1416.195 1449.675 ;
        RECT 1416.485 1200.625 1416.655 1207.595 ;
        RECT 1416.485 1074.825 1416.655 1097.095 ;
        RECT 1416.025 855.525 1416.195 903.975 ;
        RECT 1416.485 688.245 1416.655 717.655 ;
        RECT 1416.025 425.085 1416.195 517.395 ;
        RECT 1416.025 324.445 1416.195 414.035 ;
        RECT 1416.025 228.225 1416.195 275.995 ;
        RECT 1416.025 179.605 1416.195 227.715 ;
      LAYER mcon ;
        RECT 1416.025 1449.505 1416.195 1449.675 ;
        RECT 1416.485 1207.425 1416.655 1207.595 ;
        RECT 1416.485 1096.925 1416.655 1097.095 ;
        RECT 1416.025 903.805 1416.195 903.975 ;
        RECT 1416.485 717.485 1416.655 717.655 ;
        RECT 1416.025 517.225 1416.195 517.395 ;
        RECT 1416.025 413.865 1416.195 414.035 ;
        RECT 1416.025 275.825 1416.195 275.995 ;
        RECT 1416.025 227.545 1416.195 227.715 ;
      LAYER met1 ;
        RECT 1416.410 1635.640 1416.730 1635.700 ;
        RECT 1419.630 1635.640 1419.950 1635.700 ;
        RECT 1416.410 1635.500 1419.950 1635.640 ;
        RECT 1416.410 1635.440 1416.730 1635.500 ;
        RECT 1419.630 1635.440 1419.950 1635.500 ;
        RECT 1415.965 1449.660 1416.255 1449.705 ;
        RECT 1416.410 1449.660 1416.730 1449.720 ;
        RECT 1415.965 1449.520 1416.730 1449.660 ;
        RECT 1415.965 1449.475 1416.255 1449.520 ;
        RECT 1416.410 1449.460 1416.730 1449.520 ;
        RECT 1415.950 1442.180 1416.270 1442.240 ;
        RECT 1415.755 1442.040 1416.270 1442.180 ;
        RECT 1415.950 1441.980 1416.270 1442.040 ;
        RECT 1416.870 1297.680 1417.190 1297.740 ;
        RECT 1416.040 1297.540 1417.190 1297.680 ;
        RECT 1416.040 1297.400 1416.180 1297.540 ;
        RECT 1416.870 1297.480 1417.190 1297.540 ;
        RECT 1415.950 1297.140 1416.270 1297.400 ;
        RECT 1416.870 1249.200 1417.190 1249.460 ;
        RECT 1416.410 1249.060 1416.730 1249.120 ;
        RECT 1416.960 1249.060 1417.100 1249.200 ;
        RECT 1416.410 1248.920 1417.100 1249.060 ;
        RECT 1416.410 1248.860 1416.730 1248.920 ;
        RECT 1416.410 1207.580 1416.730 1207.640 ;
        RECT 1416.215 1207.440 1416.730 1207.580 ;
        RECT 1416.410 1207.380 1416.730 1207.440 ;
        RECT 1416.410 1200.780 1416.730 1200.840 ;
        RECT 1416.215 1200.640 1416.730 1200.780 ;
        RECT 1416.410 1200.580 1416.730 1200.640 ;
        RECT 1416.410 1152.300 1416.730 1152.560 ;
        RECT 1416.500 1151.880 1416.640 1152.300 ;
        RECT 1416.410 1151.620 1416.730 1151.880 ;
        RECT 1416.410 1145.360 1416.730 1145.420 ;
        RECT 1417.330 1145.360 1417.650 1145.420 ;
        RECT 1416.410 1145.220 1417.650 1145.360 ;
        RECT 1416.410 1145.160 1416.730 1145.220 ;
        RECT 1417.330 1145.160 1417.650 1145.220 ;
        RECT 1416.410 1097.080 1416.730 1097.140 ;
        RECT 1416.215 1096.940 1416.730 1097.080 ;
        RECT 1416.410 1096.880 1416.730 1096.940 ;
        RECT 1416.425 1074.980 1416.715 1075.025 ;
        RECT 1416.870 1074.980 1417.190 1075.040 ;
        RECT 1416.425 1074.840 1417.190 1074.980 ;
        RECT 1416.425 1074.795 1416.715 1074.840 ;
        RECT 1416.870 1074.780 1417.190 1074.840 ;
        RECT 1416.870 1048.800 1417.190 1048.860 ;
        RECT 1417.790 1048.800 1418.110 1048.860 ;
        RECT 1416.870 1048.660 1418.110 1048.800 ;
        RECT 1416.870 1048.600 1417.190 1048.660 ;
        RECT 1417.790 1048.600 1418.110 1048.660 ;
        RECT 1415.950 917.900 1416.270 917.960 ;
        RECT 1416.870 917.900 1417.190 917.960 ;
        RECT 1415.950 917.760 1417.190 917.900 ;
        RECT 1415.950 917.700 1416.270 917.760 ;
        RECT 1416.870 917.700 1417.190 917.760 ;
        RECT 1415.950 903.960 1416.270 904.020 ;
        RECT 1415.755 903.820 1416.270 903.960 ;
        RECT 1415.950 903.760 1416.270 903.820 ;
        RECT 1415.965 855.680 1416.255 855.725 ;
        RECT 1416.870 855.680 1417.190 855.740 ;
        RECT 1415.965 855.540 1417.190 855.680 ;
        RECT 1415.965 855.495 1416.255 855.540 ;
        RECT 1416.870 855.480 1417.190 855.540 ;
        RECT 1415.950 814.200 1416.270 814.260 ;
        RECT 1416.870 814.200 1417.190 814.260 ;
        RECT 1415.950 814.060 1417.190 814.200 ;
        RECT 1415.950 814.000 1416.270 814.060 ;
        RECT 1416.870 814.000 1417.190 814.060 ;
        RECT 1415.950 724.440 1416.270 724.500 ;
        RECT 1416.870 724.440 1417.190 724.500 ;
        RECT 1415.950 724.300 1417.190 724.440 ;
        RECT 1415.950 724.240 1416.270 724.300 ;
        RECT 1416.870 724.240 1417.190 724.300 ;
        RECT 1416.425 717.640 1416.715 717.685 ;
        RECT 1416.870 717.640 1417.190 717.700 ;
        RECT 1416.425 717.500 1417.190 717.640 ;
        RECT 1416.425 717.455 1416.715 717.500 ;
        RECT 1416.870 717.440 1417.190 717.500 ;
        RECT 1416.410 688.400 1416.730 688.460 ;
        RECT 1416.215 688.260 1416.730 688.400 ;
        RECT 1416.410 688.200 1416.730 688.260 ;
        RECT 1416.410 525.340 1416.730 525.600 ;
        RECT 1416.500 524.920 1416.640 525.340 ;
        RECT 1416.410 524.660 1416.730 524.920 ;
        RECT 1415.965 517.380 1416.255 517.425 ;
        RECT 1416.410 517.380 1416.730 517.440 ;
        RECT 1415.965 517.240 1416.730 517.380 ;
        RECT 1415.965 517.195 1416.255 517.240 ;
        RECT 1416.410 517.180 1416.730 517.240 ;
        RECT 1415.950 425.240 1416.270 425.300 ;
        RECT 1415.755 425.100 1416.270 425.240 ;
        RECT 1415.950 425.040 1416.270 425.100 ;
        RECT 1415.950 414.020 1416.270 414.080 ;
        RECT 1415.755 413.880 1416.270 414.020 ;
        RECT 1415.950 413.820 1416.270 413.880 ;
        RECT 1415.965 324.600 1416.255 324.645 ;
        RECT 1416.410 324.600 1416.730 324.660 ;
        RECT 1415.965 324.460 1416.730 324.600 ;
        RECT 1415.965 324.415 1416.255 324.460 ;
        RECT 1416.410 324.400 1416.730 324.460 ;
        RECT 1415.965 275.980 1416.255 276.025 ;
        RECT 1416.870 275.980 1417.190 276.040 ;
        RECT 1415.965 275.840 1417.190 275.980 ;
        RECT 1415.965 275.795 1416.255 275.840 ;
        RECT 1416.870 275.780 1417.190 275.840 ;
        RECT 1415.950 228.380 1416.270 228.440 ;
        RECT 1415.755 228.240 1416.270 228.380 ;
        RECT 1415.950 228.180 1416.270 228.240 ;
        RECT 1415.950 227.700 1416.270 227.760 ;
        RECT 1415.755 227.560 1416.270 227.700 ;
        RECT 1415.950 227.500 1416.270 227.560 ;
        RECT 1415.950 179.760 1416.270 179.820 ;
        RECT 1415.755 179.620 1416.270 179.760 ;
        RECT 1415.950 179.560 1416.270 179.620 ;
        RECT 1416.410 137.740 1416.730 138.000 ;
        RECT 1416.500 137.320 1416.640 137.740 ;
        RECT 1416.410 137.060 1416.730 137.320 ;
        RECT 1007.010 49.540 1007.330 49.600 ;
        RECT 1416.410 49.540 1416.730 49.600 ;
        RECT 1007.010 49.400 1416.730 49.540 ;
        RECT 1007.010 49.340 1007.330 49.400 ;
        RECT 1416.410 49.340 1416.730 49.400 ;
        RECT 1001.950 2.960 1002.270 3.020 ;
        RECT 1007.010 2.960 1007.330 3.020 ;
        RECT 1001.950 2.820 1007.330 2.960 ;
        RECT 1001.950 2.760 1002.270 2.820 ;
        RECT 1007.010 2.760 1007.330 2.820 ;
      LAYER via ;
        RECT 1416.440 1635.440 1416.700 1635.700 ;
        RECT 1419.660 1635.440 1419.920 1635.700 ;
        RECT 1416.440 1449.460 1416.700 1449.720 ;
        RECT 1415.980 1441.980 1416.240 1442.240 ;
        RECT 1416.900 1297.480 1417.160 1297.740 ;
        RECT 1415.980 1297.140 1416.240 1297.400 ;
        RECT 1416.900 1249.200 1417.160 1249.460 ;
        RECT 1416.440 1248.860 1416.700 1249.120 ;
        RECT 1416.440 1207.380 1416.700 1207.640 ;
        RECT 1416.440 1200.580 1416.700 1200.840 ;
        RECT 1416.440 1152.300 1416.700 1152.560 ;
        RECT 1416.440 1151.620 1416.700 1151.880 ;
        RECT 1416.440 1145.160 1416.700 1145.420 ;
        RECT 1417.360 1145.160 1417.620 1145.420 ;
        RECT 1416.440 1096.880 1416.700 1097.140 ;
        RECT 1416.900 1074.780 1417.160 1075.040 ;
        RECT 1416.900 1048.600 1417.160 1048.860 ;
        RECT 1417.820 1048.600 1418.080 1048.860 ;
        RECT 1415.980 917.700 1416.240 917.960 ;
        RECT 1416.900 917.700 1417.160 917.960 ;
        RECT 1415.980 903.760 1416.240 904.020 ;
        RECT 1416.900 855.480 1417.160 855.740 ;
        RECT 1415.980 814.000 1416.240 814.260 ;
        RECT 1416.900 814.000 1417.160 814.260 ;
        RECT 1415.980 724.240 1416.240 724.500 ;
        RECT 1416.900 724.240 1417.160 724.500 ;
        RECT 1416.900 717.440 1417.160 717.700 ;
        RECT 1416.440 688.200 1416.700 688.460 ;
        RECT 1416.440 525.340 1416.700 525.600 ;
        RECT 1416.440 524.660 1416.700 524.920 ;
        RECT 1416.440 517.180 1416.700 517.440 ;
        RECT 1415.980 425.040 1416.240 425.300 ;
        RECT 1415.980 413.820 1416.240 414.080 ;
        RECT 1416.440 324.400 1416.700 324.660 ;
        RECT 1416.900 275.780 1417.160 276.040 ;
        RECT 1415.980 228.180 1416.240 228.440 ;
        RECT 1415.980 227.500 1416.240 227.760 ;
        RECT 1415.980 179.560 1416.240 179.820 ;
        RECT 1416.440 137.740 1416.700 138.000 ;
        RECT 1416.440 137.060 1416.700 137.320 ;
        RECT 1007.040 49.340 1007.300 49.600 ;
        RECT 1416.440 49.340 1416.700 49.600 ;
        RECT 1001.980 2.760 1002.240 3.020 ;
        RECT 1007.040 2.760 1007.300 3.020 ;
      LAYER met2 ;
        RECT 1420.110 1700.410 1420.390 1704.000 ;
        RECT 1419.720 1700.270 1420.390 1700.410 ;
        RECT 1419.720 1635.730 1419.860 1700.270 ;
        RECT 1420.110 1700.000 1420.390 1700.270 ;
        RECT 1416.440 1635.410 1416.700 1635.730 ;
        RECT 1419.660 1635.410 1419.920 1635.730 ;
        RECT 1416.500 1449.750 1416.640 1635.410 ;
        RECT 1416.440 1449.430 1416.700 1449.750 ;
        RECT 1415.980 1441.950 1416.240 1442.270 ;
        RECT 1416.040 1400.530 1416.180 1441.950 ;
        RECT 1416.040 1400.390 1417.560 1400.530 ;
        RECT 1417.420 1398.490 1417.560 1400.390 ;
        RECT 1416.960 1398.350 1417.560 1398.490 ;
        RECT 1416.960 1297.770 1417.100 1398.350 ;
        RECT 1416.040 1297.430 1416.180 1297.585 ;
        RECT 1416.900 1297.450 1417.160 1297.770 ;
        RECT 1415.980 1297.170 1416.240 1297.430 ;
        RECT 1415.980 1297.110 1417.100 1297.170 ;
        RECT 1416.040 1297.030 1417.100 1297.110 ;
        RECT 1416.960 1249.490 1417.100 1297.030 ;
        RECT 1416.900 1249.170 1417.160 1249.490 ;
        RECT 1416.440 1248.830 1416.700 1249.150 ;
        RECT 1416.500 1207.670 1416.640 1248.830 ;
        RECT 1416.440 1207.350 1416.700 1207.670 ;
        RECT 1416.440 1200.725 1416.700 1200.870 ;
        RECT 1416.430 1200.355 1416.710 1200.725 ;
        RECT 1416.430 1199.675 1416.710 1200.045 ;
        RECT 1416.500 1152.590 1416.640 1199.675 ;
        RECT 1416.440 1152.270 1416.700 1152.590 ;
        RECT 1416.440 1151.590 1416.700 1151.910 ;
        RECT 1416.500 1145.450 1416.640 1151.590 ;
        RECT 1416.440 1145.130 1416.700 1145.450 ;
        RECT 1417.360 1145.130 1417.620 1145.450 ;
        RECT 1417.420 1097.365 1417.560 1145.130 ;
        RECT 1416.430 1096.995 1416.710 1097.365 ;
        RECT 1417.350 1096.995 1417.630 1097.365 ;
        RECT 1416.440 1096.850 1416.700 1096.995 ;
        RECT 1416.900 1074.750 1417.160 1075.070 ;
        RECT 1416.960 1048.890 1417.100 1074.750 ;
        RECT 1416.900 1048.570 1417.160 1048.890 ;
        RECT 1417.820 1048.570 1418.080 1048.890 ;
        RECT 1417.880 1000.805 1418.020 1048.570 ;
        RECT 1416.430 1000.435 1416.710 1000.805 ;
        RECT 1417.810 1000.435 1418.090 1000.805 ;
        RECT 1416.500 942.210 1416.640 1000.435 ;
        RECT 1416.500 942.070 1417.100 942.210 ;
        RECT 1416.960 917.990 1417.100 942.070 ;
        RECT 1415.980 917.670 1416.240 917.990 ;
        RECT 1416.900 917.670 1417.160 917.990 ;
        RECT 1416.040 904.050 1416.180 917.670 ;
        RECT 1415.980 903.730 1416.240 904.050 ;
        RECT 1416.900 855.450 1417.160 855.770 ;
        RECT 1416.960 834.770 1417.100 855.450 ;
        RECT 1416.040 834.630 1417.100 834.770 ;
        RECT 1416.040 814.290 1416.180 834.630 ;
        RECT 1415.980 813.970 1416.240 814.290 ;
        RECT 1416.900 813.970 1417.160 814.290 ;
        RECT 1416.960 724.725 1417.100 813.970 ;
        RECT 1415.970 724.355 1416.250 724.725 ;
        RECT 1416.890 724.355 1417.170 724.725 ;
        RECT 1415.980 724.210 1416.240 724.355 ;
        RECT 1416.900 724.210 1417.160 724.355 ;
        RECT 1416.960 717.730 1417.100 724.210 ;
        RECT 1416.900 717.410 1417.160 717.730 ;
        RECT 1416.440 688.170 1416.700 688.490 ;
        RECT 1416.500 573.765 1416.640 688.170 ;
        RECT 1416.430 573.395 1416.710 573.765 ;
        RECT 1415.970 572.970 1416.250 573.085 ;
        RECT 1415.970 572.830 1416.640 572.970 ;
        RECT 1415.970 572.715 1416.250 572.830 ;
        RECT 1416.500 525.630 1416.640 572.830 ;
        RECT 1416.440 525.310 1416.700 525.630 ;
        RECT 1416.440 524.630 1416.700 524.950 ;
        RECT 1416.500 517.470 1416.640 524.630 ;
        RECT 1416.440 517.150 1416.700 517.470 ;
        RECT 1415.980 425.010 1416.240 425.330 ;
        RECT 1416.040 414.110 1416.180 425.010 ;
        RECT 1415.980 413.790 1416.240 414.110 ;
        RECT 1416.440 324.370 1416.700 324.690 ;
        RECT 1416.500 282.610 1416.640 324.370 ;
        RECT 1416.500 282.470 1417.100 282.610 ;
        RECT 1416.960 276.070 1417.100 282.470 ;
        RECT 1416.900 275.750 1417.160 276.070 ;
        RECT 1415.980 228.150 1416.240 228.470 ;
        RECT 1416.040 227.790 1416.180 228.150 ;
        RECT 1415.980 227.470 1416.240 227.790 ;
        RECT 1415.980 179.530 1416.240 179.850 ;
        RECT 1416.040 157.490 1416.180 179.530 ;
        RECT 1416.040 157.350 1416.640 157.490 ;
        RECT 1416.500 138.030 1416.640 157.350 ;
        RECT 1416.440 137.710 1416.700 138.030 ;
        RECT 1416.440 137.030 1416.700 137.350 ;
        RECT 1416.500 49.630 1416.640 137.030 ;
        RECT 1007.040 49.310 1007.300 49.630 ;
        RECT 1416.440 49.310 1416.700 49.630 ;
        RECT 1007.100 3.050 1007.240 49.310 ;
        RECT 1001.980 2.730 1002.240 3.050 ;
        RECT 1007.040 2.730 1007.300 3.050 ;
        RECT 1002.040 2.400 1002.180 2.730 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
      LAYER via2 ;
        RECT 1416.430 1200.400 1416.710 1200.680 ;
        RECT 1416.430 1199.720 1416.710 1200.000 ;
        RECT 1416.430 1097.040 1416.710 1097.320 ;
        RECT 1417.350 1097.040 1417.630 1097.320 ;
        RECT 1416.430 1000.480 1416.710 1000.760 ;
        RECT 1417.810 1000.480 1418.090 1000.760 ;
        RECT 1415.970 724.400 1416.250 724.680 ;
        RECT 1416.890 724.400 1417.170 724.680 ;
        RECT 1416.430 573.440 1416.710 573.720 ;
        RECT 1415.970 572.760 1416.250 573.040 ;
      LAYER met3 ;
        RECT 1416.405 1200.690 1416.735 1200.705 ;
        RECT 1416.190 1200.375 1416.735 1200.690 ;
        RECT 1416.190 1200.025 1416.490 1200.375 ;
        RECT 1416.190 1199.710 1416.735 1200.025 ;
        RECT 1416.405 1199.695 1416.735 1199.710 ;
        RECT 1416.405 1097.330 1416.735 1097.345 ;
        RECT 1417.325 1097.330 1417.655 1097.345 ;
        RECT 1416.405 1097.030 1417.655 1097.330 ;
        RECT 1416.405 1097.015 1416.735 1097.030 ;
        RECT 1417.325 1097.015 1417.655 1097.030 ;
        RECT 1416.405 1000.770 1416.735 1000.785 ;
        RECT 1417.785 1000.770 1418.115 1000.785 ;
        RECT 1416.405 1000.470 1418.115 1000.770 ;
        RECT 1416.405 1000.455 1416.735 1000.470 ;
        RECT 1417.785 1000.455 1418.115 1000.470 ;
        RECT 1415.945 724.690 1416.275 724.705 ;
        RECT 1416.865 724.690 1417.195 724.705 ;
        RECT 1415.945 724.390 1417.195 724.690 ;
        RECT 1415.945 724.375 1416.275 724.390 ;
        RECT 1416.865 724.375 1417.195 724.390 ;
        RECT 1416.405 573.730 1416.735 573.745 ;
        RECT 1416.190 573.415 1416.735 573.730 ;
        RECT 1416.190 573.065 1416.490 573.415 ;
        RECT 1415.945 572.750 1416.490 573.065 ;
        RECT 1415.945 572.735 1416.275 572.750 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 0.300 ;
=======
      LAYER li1 ;
        RECT 1423.385 1635.485 1423.555 1683.595 ;
        RECT 1423.385 1442.025 1423.555 1490.475 ;
        RECT 1423.845 1352.605 1424.015 1400.715 ;
        RECT 1423.385 814.385 1423.555 862.495 ;
        RECT 1422.925 427.805 1423.095 475.915 ;
        RECT 1423.385 49.045 1423.555 113.815 ;
      LAYER mcon ;
        RECT 1423.385 1683.425 1423.555 1683.595 ;
        RECT 1423.385 1490.305 1423.555 1490.475 ;
        RECT 1423.845 1400.545 1424.015 1400.715 ;
        RECT 1423.385 862.325 1423.555 862.495 ;
        RECT 1422.925 475.745 1423.095 475.915 ;
        RECT 1423.385 113.645 1423.555 113.815 ;
      LAYER met1 ;
        RECT 1423.325 1683.580 1423.615 1683.625 ;
        RECT 1424.230 1683.580 1424.550 1683.640 ;
        RECT 1423.325 1683.440 1424.550 1683.580 ;
        RECT 1423.325 1683.395 1423.615 1683.440 ;
        RECT 1424.230 1683.380 1424.550 1683.440 ;
        RECT 1423.310 1635.640 1423.630 1635.700 ;
        RECT 1423.115 1635.500 1423.630 1635.640 ;
        RECT 1423.310 1635.440 1423.630 1635.500 ;
        RECT 1423.310 1545.880 1423.630 1545.940 ;
        RECT 1423.770 1545.880 1424.090 1545.940 ;
        RECT 1423.310 1545.740 1424.090 1545.880 ;
        RECT 1423.310 1545.680 1423.630 1545.740 ;
        RECT 1423.770 1545.680 1424.090 1545.740 ;
        RECT 1423.325 1490.460 1423.615 1490.505 ;
        RECT 1423.770 1490.460 1424.090 1490.520 ;
        RECT 1423.325 1490.320 1424.090 1490.460 ;
        RECT 1423.325 1490.275 1423.615 1490.320 ;
        RECT 1423.770 1490.260 1424.090 1490.320 ;
        RECT 1423.310 1442.180 1423.630 1442.240 ;
        RECT 1423.115 1442.040 1423.630 1442.180 ;
        RECT 1423.310 1441.980 1423.630 1442.040 ;
        RECT 1423.770 1400.700 1424.090 1400.760 ;
        RECT 1423.575 1400.560 1424.090 1400.700 ;
        RECT 1423.770 1400.500 1424.090 1400.560 ;
        RECT 1423.770 1352.760 1424.090 1352.820 ;
        RECT 1423.575 1352.620 1424.090 1352.760 ;
        RECT 1423.770 1352.560 1424.090 1352.620 ;
        RECT 1423.310 1303.940 1423.630 1304.200 ;
        RECT 1423.400 1303.800 1423.540 1303.940 ;
        RECT 1423.770 1303.800 1424.090 1303.860 ;
        RECT 1423.400 1303.660 1424.090 1303.800 ;
        RECT 1423.770 1303.600 1424.090 1303.660 ;
        RECT 1423.770 1159.640 1424.090 1159.700 ;
        RECT 1423.400 1159.500 1424.090 1159.640 ;
        RECT 1423.400 1159.360 1423.540 1159.500 ;
        RECT 1423.770 1159.440 1424.090 1159.500 ;
        RECT 1423.310 1159.100 1423.630 1159.360 ;
        RECT 1423.770 966.520 1424.090 966.580 ;
        RECT 1423.400 966.380 1424.090 966.520 ;
        RECT 1423.400 966.240 1423.540 966.380 ;
        RECT 1423.770 966.320 1424.090 966.380 ;
        RECT 1423.310 965.980 1423.630 966.240 ;
        RECT 1423.325 862.480 1423.615 862.525 ;
        RECT 1423.770 862.480 1424.090 862.540 ;
        RECT 1423.325 862.340 1424.090 862.480 ;
        RECT 1423.325 862.295 1423.615 862.340 ;
        RECT 1423.770 862.280 1424.090 862.340 ;
        RECT 1423.310 814.540 1423.630 814.600 ;
        RECT 1423.115 814.400 1423.630 814.540 ;
        RECT 1423.310 814.340 1423.630 814.400 ;
        RECT 1423.310 787.140 1423.630 787.400 ;
        RECT 1423.400 786.720 1423.540 787.140 ;
        RECT 1423.310 786.460 1423.630 786.720 ;
        RECT 1423.310 724.440 1423.630 724.500 ;
        RECT 1424.230 724.440 1424.550 724.500 ;
        RECT 1423.310 724.300 1424.550 724.440 ;
        RECT 1423.310 724.240 1423.630 724.300 ;
        RECT 1424.230 724.240 1424.550 724.300 ;
        RECT 1423.310 627.880 1423.630 627.940 ;
        RECT 1423.770 627.880 1424.090 627.940 ;
        RECT 1423.310 627.740 1424.090 627.880 ;
        RECT 1423.310 627.680 1423.630 627.740 ;
        RECT 1423.770 627.680 1424.090 627.740 ;
        RECT 1422.865 475.900 1423.155 475.945 ;
        RECT 1423.310 475.900 1423.630 475.960 ;
        RECT 1422.865 475.760 1423.630 475.900 ;
        RECT 1422.865 475.715 1423.155 475.760 ;
        RECT 1423.310 475.700 1423.630 475.760 ;
        RECT 1422.850 427.960 1423.170 428.020 ;
        RECT 1422.655 427.820 1423.170 427.960 ;
        RECT 1422.850 427.760 1423.170 427.820 ;
        RECT 1423.770 255.580 1424.090 255.640 ;
        RECT 1423.400 255.440 1424.090 255.580 ;
        RECT 1423.400 255.300 1423.540 255.440 ;
        RECT 1423.770 255.380 1424.090 255.440 ;
        RECT 1423.310 255.040 1423.630 255.300 ;
        RECT 1422.850 186.560 1423.170 186.620 ;
        RECT 1423.770 186.560 1424.090 186.620 ;
        RECT 1422.850 186.420 1424.090 186.560 ;
        RECT 1422.850 186.360 1423.170 186.420 ;
        RECT 1423.770 186.360 1424.090 186.420 ;
        RECT 1423.325 113.800 1423.615 113.845 ;
        RECT 1424.230 113.800 1424.550 113.860 ;
        RECT 1423.325 113.660 1424.550 113.800 ;
        RECT 1423.325 113.615 1423.615 113.660 ;
        RECT 1424.230 113.600 1424.550 113.660 ;
        RECT 1020.810 49.200 1021.130 49.260 ;
        RECT 1423.325 49.200 1423.615 49.245 ;
        RECT 1020.810 49.060 1423.615 49.200 ;
        RECT 1020.810 49.000 1021.130 49.060 ;
        RECT 1423.325 49.015 1423.615 49.060 ;
      LAYER via ;
        RECT 1424.260 1683.380 1424.520 1683.640 ;
        RECT 1423.340 1635.440 1423.600 1635.700 ;
        RECT 1423.340 1545.680 1423.600 1545.940 ;
        RECT 1423.800 1545.680 1424.060 1545.940 ;
        RECT 1423.800 1490.260 1424.060 1490.520 ;
        RECT 1423.340 1441.980 1423.600 1442.240 ;
        RECT 1423.800 1400.500 1424.060 1400.760 ;
        RECT 1423.800 1352.560 1424.060 1352.820 ;
        RECT 1423.340 1303.940 1423.600 1304.200 ;
        RECT 1423.800 1303.600 1424.060 1303.860 ;
        RECT 1423.800 1159.440 1424.060 1159.700 ;
        RECT 1423.340 1159.100 1423.600 1159.360 ;
        RECT 1423.800 966.320 1424.060 966.580 ;
        RECT 1423.340 965.980 1423.600 966.240 ;
        RECT 1423.800 862.280 1424.060 862.540 ;
        RECT 1423.340 814.340 1423.600 814.600 ;
        RECT 1423.340 787.140 1423.600 787.400 ;
        RECT 1423.340 786.460 1423.600 786.720 ;
        RECT 1423.340 724.240 1423.600 724.500 ;
        RECT 1424.260 724.240 1424.520 724.500 ;
        RECT 1423.340 627.680 1423.600 627.940 ;
        RECT 1423.800 627.680 1424.060 627.940 ;
        RECT 1423.340 475.700 1423.600 475.960 ;
        RECT 1422.880 427.760 1423.140 428.020 ;
        RECT 1423.800 255.380 1424.060 255.640 ;
        RECT 1423.340 255.040 1423.600 255.300 ;
        RECT 1422.880 186.360 1423.140 186.620 ;
        RECT 1423.800 186.360 1424.060 186.620 ;
        RECT 1424.260 113.600 1424.520 113.860 ;
        RECT 1020.840 49.000 1021.100 49.260 ;
      LAYER met2 ;
        RECT 1425.170 1700.410 1425.450 1704.000 ;
        RECT 1424.780 1700.270 1425.450 1700.410 ;
        RECT 1424.780 1686.640 1424.920 1700.270 ;
        RECT 1425.170 1700.000 1425.450 1700.270 ;
        RECT 1424.320 1686.500 1424.920 1686.640 ;
        RECT 1424.320 1683.670 1424.460 1686.500 ;
        RECT 1424.260 1683.350 1424.520 1683.670 ;
        RECT 1423.340 1635.410 1423.600 1635.730 ;
        RECT 1423.400 1545.970 1423.540 1635.410 ;
        RECT 1423.340 1545.650 1423.600 1545.970 ;
        RECT 1423.800 1545.650 1424.060 1545.970 ;
        RECT 1423.860 1490.550 1424.000 1545.650 ;
        RECT 1423.800 1490.230 1424.060 1490.550 ;
        RECT 1423.340 1441.950 1423.600 1442.270 ;
        RECT 1423.400 1425.010 1423.540 1441.950 ;
        RECT 1423.400 1424.870 1424.000 1425.010 ;
        RECT 1423.860 1400.790 1424.000 1424.870 ;
        RECT 1423.800 1400.470 1424.060 1400.790 ;
        RECT 1423.800 1352.530 1424.060 1352.850 ;
        RECT 1423.860 1316.890 1424.000 1352.530 ;
        RECT 1423.400 1316.750 1424.000 1316.890 ;
        RECT 1423.400 1304.230 1423.540 1316.750 ;
        RECT 1423.340 1303.910 1423.600 1304.230 ;
        RECT 1423.800 1303.570 1424.060 1303.890 ;
        RECT 1423.860 1159.730 1424.000 1303.570 ;
        RECT 1423.800 1159.410 1424.060 1159.730 ;
        RECT 1423.340 1159.070 1423.600 1159.390 ;
        RECT 1423.400 1136.010 1423.540 1159.070 ;
        RECT 1423.400 1135.870 1424.460 1136.010 ;
        RECT 1424.320 1124.450 1424.460 1135.870 ;
        RECT 1423.860 1124.310 1424.460 1124.450 ;
        RECT 1423.860 966.610 1424.000 1124.310 ;
        RECT 1423.800 966.290 1424.060 966.610 ;
        RECT 1423.340 965.950 1423.600 966.270 ;
        RECT 1423.400 917.900 1423.540 965.950 ;
        RECT 1423.400 917.760 1424.000 917.900 ;
        RECT 1423.860 862.570 1424.000 917.760 ;
        RECT 1423.800 862.250 1424.060 862.570 ;
        RECT 1423.340 814.310 1423.600 814.630 ;
        RECT 1423.400 787.430 1423.540 814.310 ;
        RECT 1423.340 787.110 1423.600 787.430 ;
        RECT 1423.340 786.430 1423.600 786.750 ;
        RECT 1423.400 724.530 1423.540 786.430 ;
        RECT 1423.340 724.210 1423.600 724.530 ;
        RECT 1424.260 724.210 1424.520 724.530 ;
        RECT 1424.320 699.450 1424.460 724.210 ;
        RECT 1423.860 699.310 1424.460 699.450 ;
        RECT 1423.860 651.850 1424.000 699.310 ;
        RECT 1423.400 651.710 1424.000 651.850 ;
        RECT 1423.400 627.970 1423.540 651.710 ;
        RECT 1423.340 627.650 1423.600 627.970 ;
        RECT 1423.800 627.650 1424.060 627.970 ;
        RECT 1423.860 531.320 1424.000 627.650 ;
        RECT 1423.860 531.180 1424.460 531.320 ;
        RECT 1424.320 483.325 1424.460 531.180 ;
        RECT 1423.330 482.955 1423.610 483.325 ;
        RECT 1424.250 482.955 1424.530 483.325 ;
        RECT 1423.400 475.990 1423.540 482.955 ;
        RECT 1423.340 475.670 1423.600 475.990 ;
        RECT 1422.880 427.730 1423.140 428.050 ;
        RECT 1422.940 404.330 1423.080 427.730 ;
        RECT 1422.940 404.190 1424.000 404.330 ;
        RECT 1423.860 255.670 1424.000 404.190 ;
        RECT 1423.800 255.350 1424.060 255.670 ;
        RECT 1423.340 255.010 1423.600 255.330 ;
        RECT 1423.400 234.330 1423.540 255.010 ;
        RECT 1422.940 234.190 1423.540 234.330 ;
        RECT 1422.940 186.650 1423.080 234.190 ;
        RECT 1422.880 186.330 1423.140 186.650 ;
        RECT 1423.800 186.330 1424.060 186.650 ;
        RECT 1423.860 186.050 1424.000 186.330 ;
        RECT 1423.860 185.910 1424.460 186.050 ;
        RECT 1424.320 113.890 1424.460 185.910 ;
        RECT 1424.260 113.570 1424.520 113.890 ;
        RECT 1020.840 48.970 1021.100 49.290 ;
        RECT 1020.900 3.130 1021.040 48.970 ;
        RECT 1019.520 2.990 1021.040 3.130 ;
        RECT 1019.520 2.400 1019.660 2.990 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
      LAYER via2 ;
        RECT 1423.330 483.000 1423.610 483.280 ;
        RECT 1424.250 483.000 1424.530 483.280 ;
      LAYER met3 ;
        RECT 1423.305 483.290 1423.635 483.305 ;
        RECT 1424.225 483.290 1424.555 483.305 ;
        RECT 1423.305 482.990 1424.555 483.290 ;
        RECT 1423.305 482.975 1423.635 482.990 ;
        RECT 1424.225 482.975 1424.555 482.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1037.370 43.760 1037.690 43.820 ;
        RECT 1429.750 43.760 1430.070 43.820 ;
        RECT 1037.370 43.620 1430.070 43.760 ;
        RECT 1037.370 43.560 1037.690 43.620 ;
        RECT 1429.750 43.560 1430.070 43.620 ;
      LAYER via ;
        RECT 1037.400 43.560 1037.660 43.820 ;
        RECT 1429.780 43.560 1430.040 43.820 ;
      LAYER met2 ;
        RECT 1429.770 1700.000 1430.050 1704.000 ;
        RECT 1429.840 43.850 1429.980 1700.000 ;
        RECT 1037.400 43.530 1037.660 43.850 ;
        RECT 1429.780 43.530 1430.040 43.850 ;
        RECT 1037.460 2.400 1037.600 43.530 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1430.210 1678.140 1430.530 1678.200 ;
        RECT 1433.430 1678.140 1433.750 1678.200 ;
        RECT 1430.210 1678.000 1433.750 1678.140 ;
        RECT 1430.210 1677.940 1430.530 1678.000 ;
        RECT 1433.430 1677.940 1433.750 1678.000 ;
        RECT 1055.310 43.420 1055.630 43.480 ;
        RECT 1430.210 43.420 1430.530 43.480 ;
        RECT 1055.310 43.280 1430.530 43.420 ;
        RECT 1055.310 43.220 1055.630 43.280 ;
        RECT 1430.210 43.220 1430.530 43.280 ;
      LAYER via ;
        RECT 1430.240 1677.940 1430.500 1678.200 ;
        RECT 1433.460 1677.940 1433.720 1678.200 ;
        RECT 1055.340 43.220 1055.600 43.480 ;
        RECT 1430.240 43.220 1430.500 43.480 ;
      LAYER met2 ;
        RECT 1434.830 1700.410 1435.110 1704.000 ;
        RECT 1433.520 1700.270 1435.110 1700.410 ;
        RECT 1433.520 1678.230 1433.660 1700.270 ;
        RECT 1434.830 1700.000 1435.110 1700.270 ;
        RECT 1430.240 1677.910 1430.500 1678.230 ;
        RECT 1433.460 1677.910 1433.720 1678.230 ;
        RECT 1430.300 43.510 1430.440 1677.910 ;
        RECT 1055.340 43.190 1055.600 43.510 ;
        RECT 1430.240 43.190 1430.500 43.510 ;
        RECT 1055.400 2.400 1055.540 43.190 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1436.650 1692.420 1436.970 1692.480 ;
        RECT 1439.410 1692.420 1439.730 1692.480 ;
        RECT 1436.650 1692.280 1439.730 1692.420 ;
        RECT 1436.650 1692.220 1436.970 1692.280 ;
        RECT 1439.410 1692.220 1439.730 1692.280 ;
        RECT 1073.250 43.080 1073.570 43.140 ;
        RECT 1436.650 43.080 1436.970 43.140 ;
        RECT 1073.250 42.940 1436.970 43.080 ;
        RECT 1073.250 42.880 1073.570 42.940 ;
        RECT 1436.650 42.880 1436.970 42.940 ;
      LAYER via ;
        RECT 1436.680 1692.220 1436.940 1692.480 ;
        RECT 1439.440 1692.220 1439.700 1692.480 ;
        RECT 1073.280 42.880 1073.540 43.140 ;
        RECT 1436.680 42.880 1436.940 43.140 ;
      LAYER met2 ;
        RECT 1439.430 1700.000 1439.710 1704.000 ;
        RECT 1439.500 1692.510 1439.640 1700.000 ;
        RECT 1436.680 1692.190 1436.940 1692.510 ;
        RECT 1439.440 1692.190 1439.700 1692.510 ;
        RECT 1436.740 43.170 1436.880 1692.190 ;
        RECT 1073.280 42.850 1073.540 43.170 ;
        RECT 1436.680 42.850 1436.940 43.170 ;
        RECT 1073.340 2.400 1073.480 42.850 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1090.730 42.740 1091.050 42.800 ;
        RECT 1443.550 42.740 1443.870 42.800 ;
        RECT 1090.730 42.600 1443.870 42.740 ;
        RECT 1090.730 42.540 1091.050 42.600 ;
        RECT 1443.550 42.540 1443.870 42.600 ;
      LAYER via ;
        RECT 1090.760 42.540 1091.020 42.800 ;
        RECT 1443.580 42.540 1443.840 42.800 ;
      LAYER met2 ;
        RECT 1444.490 1700.410 1444.770 1704.000 ;
        RECT 1443.640 1700.270 1444.770 1700.410 ;
        RECT 1443.640 42.830 1443.780 1700.270 ;
        RECT 1444.490 1700.000 1444.770 1700.270 ;
        RECT 1090.760 42.510 1091.020 42.830 ;
        RECT 1443.580 42.510 1443.840 42.830 ;
        RECT 1090.820 2.400 1090.960 42.510 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 0.300 ;
=======
      LAYER li1 ;
        RECT 1450.065 1607.605 1450.235 1635.315 ;
        RECT 1450.065 1400.885 1450.235 1562.895 ;
        RECT 1450.065 1158.805 1450.235 1200.115 ;
        RECT 1450.065 1062.585 1450.235 1128.375 ;
        RECT 1450.525 869.805 1450.695 917.575 ;
        RECT 1450.065 662.405 1450.235 676.855 ;
        RECT 1450.065 403.665 1450.235 434.435 ;
        RECT 1450.065 96.645 1450.235 144.755 ;
        RECT 1450.065 42.245 1450.235 48.195 ;
      LAYER mcon ;
        RECT 1450.065 1635.145 1450.235 1635.315 ;
        RECT 1450.065 1562.725 1450.235 1562.895 ;
        RECT 1450.065 1199.945 1450.235 1200.115 ;
        RECT 1450.065 1128.205 1450.235 1128.375 ;
        RECT 1450.525 917.405 1450.695 917.575 ;
        RECT 1450.065 676.685 1450.235 676.855 ;
        RECT 1450.065 434.265 1450.235 434.435 ;
        RECT 1450.065 144.585 1450.235 144.755 ;
        RECT 1450.065 48.025 1450.235 48.195 ;
      LAYER met1 ;
        RECT 1449.070 1656.380 1449.390 1656.440 ;
        RECT 1449.990 1656.380 1450.310 1656.440 ;
        RECT 1449.070 1656.240 1450.310 1656.380 ;
        RECT 1449.070 1656.180 1449.390 1656.240 ;
        RECT 1449.990 1656.180 1450.310 1656.240 ;
        RECT 1449.990 1635.300 1450.310 1635.360 ;
        RECT 1449.795 1635.160 1450.310 1635.300 ;
        RECT 1449.990 1635.100 1450.310 1635.160 ;
        RECT 1450.005 1607.760 1450.295 1607.805 ;
        RECT 1451.830 1607.760 1452.150 1607.820 ;
        RECT 1450.005 1607.620 1452.150 1607.760 ;
        RECT 1450.005 1607.575 1450.295 1607.620 ;
        RECT 1451.830 1607.560 1452.150 1607.620 ;
        RECT 1450.005 1562.880 1450.295 1562.925 ;
        RECT 1451.830 1562.880 1452.150 1562.940 ;
        RECT 1450.005 1562.740 1452.150 1562.880 ;
        RECT 1450.005 1562.695 1450.295 1562.740 ;
        RECT 1451.830 1562.680 1452.150 1562.740 ;
        RECT 1449.990 1401.040 1450.310 1401.100 ;
        RECT 1449.795 1400.900 1450.310 1401.040 ;
        RECT 1449.990 1400.840 1450.310 1400.900 ;
        RECT 1449.070 1297.340 1449.390 1297.400 ;
        RECT 1449.990 1297.340 1450.310 1297.400 ;
        RECT 1449.070 1297.200 1450.310 1297.340 ;
        RECT 1449.070 1297.140 1449.390 1297.200 ;
        RECT 1449.990 1297.140 1450.310 1297.200 ;
        RECT 1449.990 1249.060 1450.310 1249.120 ;
        RECT 1450.450 1249.060 1450.770 1249.120 ;
        RECT 1449.990 1248.920 1450.770 1249.060 ;
        RECT 1449.990 1248.860 1450.310 1248.920 ;
        RECT 1450.450 1248.860 1450.770 1248.920 ;
        RECT 1449.990 1200.100 1450.310 1200.160 ;
        RECT 1449.795 1199.960 1450.310 1200.100 ;
        RECT 1449.990 1199.900 1450.310 1199.960 ;
        RECT 1449.990 1158.960 1450.310 1159.020 ;
        RECT 1449.795 1158.820 1450.310 1158.960 ;
        RECT 1449.990 1158.760 1450.310 1158.820 ;
        RECT 1449.990 1128.360 1450.310 1128.420 ;
        RECT 1449.795 1128.220 1450.310 1128.360 ;
        RECT 1449.990 1128.160 1450.310 1128.220 ;
        RECT 1450.005 1062.740 1450.295 1062.785 ;
        RECT 1450.450 1062.740 1450.770 1062.800 ;
        RECT 1450.005 1062.600 1450.770 1062.740 ;
        RECT 1450.005 1062.555 1450.295 1062.600 ;
        RECT 1450.450 1062.540 1450.770 1062.600 ;
        RECT 1449.070 1014.460 1449.390 1014.520 ;
        RECT 1449.990 1014.460 1450.310 1014.520 ;
        RECT 1449.070 1014.320 1450.310 1014.460 ;
        RECT 1449.070 1014.260 1449.390 1014.320 ;
        RECT 1449.990 1014.260 1450.310 1014.320 ;
        RECT 1449.070 917.900 1449.390 917.960 ;
        RECT 1449.990 917.900 1450.310 917.960 ;
        RECT 1449.070 917.760 1450.310 917.900 ;
        RECT 1449.070 917.700 1449.390 917.760 ;
        RECT 1449.990 917.700 1450.310 917.760 ;
        RECT 1450.450 917.560 1450.770 917.620 ;
        RECT 1450.255 917.420 1450.770 917.560 ;
        RECT 1450.450 917.360 1450.770 917.420 ;
        RECT 1450.450 869.960 1450.770 870.020 ;
        RECT 1450.255 869.820 1450.770 869.960 ;
        RECT 1450.450 869.760 1450.770 869.820 ;
        RECT 1449.070 772.720 1449.390 772.780 ;
        RECT 1450.450 772.720 1450.770 772.780 ;
        RECT 1449.070 772.580 1450.770 772.720 ;
        RECT 1449.070 772.520 1449.390 772.580 ;
        RECT 1450.450 772.520 1450.770 772.580 ;
        RECT 1449.990 676.840 1450.310 676.900 ;
        RECT 1449.795 676.700 1450.310 676.840 ;
        RECT 1449.990 676.640 1450.310 676.700 ;
        RECT 1449.990 662.560 1450.310 662.620 ;
        RECT 1449.795 662.420 1450.310 662.560 ;
        RECT 1449.990 662.360 1450.310 662.420 ;
        RECT 1449.990 651.140 1450.310 651.400 ;
        RECT 1450.080 650.720 1450.220 651.140 ;
        RECT 1449.990 650.460 1450.310 650.720 ;
        RECT 1449.990 593.680 1450.310 593.940 ;
        RECT 1450.080 593.260 1450.220 593.680 ;
        RECT 1449.990 593.000 1450.310 593.260 ;
        RECT 1449.990 531.320 1450.310 531.380 ;
        RECT 1450.450 531.320 1450.770 531.380 ;
        RECT 1449.990 531.180 1450.770 531.320 ;
        RECT 1449.990 531.120 1450.310 531.180 ;
        RECT 1450.450 531.120 1450.770 531.180 ;
        RECT 1449.070 524.180 1449.390 524.240 ;
        RECT 1450.450 524.180 1450.770 524.240 ;
        RECT 1449.070 524.040 1450.770 524.180 ;
        RECT 1449.070 523.980 1449.390 524.040 ;
        RECT 1450.450 523.980 1450.770 524.040 ;
        RECT 1449.990 434.420 1450.310 434.480 ;
        RECT 1449.795 434.280 1450.310 434.420 ;
        RECT 1449.990 434.220 1450.310 434.280 ;
        RECT 1450.005 403.820 1450.295 403.865 ;
        RECT 1450.450 403.820 1450.770 403.880 ;
        RECT 1450.005 403.680 1450.770 403.820 ;
        RECT 1450.005 403.635 1450.295 403.680 ;
        RECT 1450.450 403.620 1450.770 403.680 ;
        RECT 1449.070 310.660 1449.390 310.720 ;
        RECT 1449.990 310.660 1450.310 310.720 ;
        RECT 1449.070 310.520 1450.310 310.660 ;
        RECT 1449.070 310.460 1449.390 310.520 ;
        RECT 1449.990 310.460 1450.310 310.520 ;
        RECT 1449.070 295.020 1449.390 295.080 ;
        RECT 1449.990 295.020 1450.310 295.080 ;
        RECT 1449.070 294.880 1450.310 295.020 ;
        RECT 1449.070 294.820 1449.390 294.880 ;
        RECT 1449.990 294.820 1450.310 294.880 ;
        RECT 1449.070 241.640 1449.390 241.700 ;
        RECT 1449.990 241.640 1450.310 241.700 ;
        RECT 1449.070 241.500 1450.310 241.640 ;
        RECT 1449.070 241.440 1449.390 241.500 ;
        RECT 1449.990 241.440 1450.310 241.500 ;
        RECT 1449.990 144.740 1450.310 144.800 ;
        RECT 1449.795 144.600 1450.310 144.740 ;
        RECT 1449.990 144.540 1450.310 144.600 ;
        RECT 1450.005 96.800 1450.295 96.845 ;
        RECT 1450.450 96.800 1450.770 96.860 ;
        RECT 1450.005 96.660 1450.770 96.800 ;
        RECT 1450.005 96.615 1450.295 96.660 ;
        RECT 1450.450 96.600 1450.770 96.660 ;
        RECT 1450.450 62.460 1450.770 62.520 ;
        RECT 1450.080 62.320 1450.770 62.460 ;
        RECT 1450.080 62.180 1450.220 62.320 ;
        RECT 1450.450 62.260 1450.770 62.320 ;
        RECT 1449.990 61.920 1450.310 62.180 ;
        RECT 1449.990 48.180 1450.310 48.240 ;
        RECT 1449.795 48.040 1450.310 48.180 ;
        RECT 1449.990 47.980 1450.310 48.040 ;
        RECT 1108.670 42.400 1108.990 42.460 ;
        RECT 1450.005 42.400 1450.295 42.445 ;
        RECT 1108.670 42.260 1450.295 42.400 ;
        RECT 1108.670 42.200 1108.990 42.260 ;
        RECT 1450.005 42.215 1450.295 42.260 ;
      LAYER via ;
        RECT 1449.100 1656.180 1449.360 1656.440 ;
        RECT 1450.020 1656.180 1450.280 1656.440 ;
        RECT 1450.020 1635.100 1450.280 1635.360 ;
        RECT 1451.860 1607.560 1452.120 1607.820 ;
        RECT 1451.860 1562.680 1452.120 1562.940 ;
        RECT 1450.020 1400.840 1450.280 1401.100 ;
        RECT 1449.100 1297.140 1449.360 1297.400 ;
        RECT 1450.020 1297.140 1450.280 1297.400 ;
        RECT 1450.020 1248.860 1450.280 1249.120 ;
        RECT 1450.480 1248.860 1450.740 1249.120 ;
        RECT 1450.020 1199.900 1450.280 1200.160 ;
        RECT 1450.020 1158.760 1450.280 1159.020 ;
        RECT 1450.020 1128.160 1450.280 1128.420 ;
        RECT 1450.480 1062.540 1450.740 1062.800 ;
        RECT 1449.100 1014.260 1449.360 1014.520 ;
        RECT 1450.020 1014.260 1450.280 1014.520 ;
        RECT 1449.100 917.700 1449.360 917.960 ;
        RECT 1450.020 917.700 1450.280 917.960 ;
        RECT 1450.480 917.360 1450.740 917.620 ;
        RECT 1450.480 869.760 1450.740 870.020 ;
        RECT 1449.100 772.520 1449.360 772.780 ;
        RECT 1450.480 772.520 1450.740 772.780 ;
        RECT 1450.020 676.640 1450.280 676.900 ;
        RECT 1450.020 662.360 1450.280 662.620 ;
        RECT 1450.020 651.140 1450.280 651.400 ;
        RECT 1450.020 650.460 1450.280 650.720 ;
        RECT 1450.020 593.680 1450.280 593.940 ;
        RECT 1450.020 593.000 1450.280 593.260 ;
        RECT 1450.020 531.120 1450.280 531.380 ;
        RECT 1450.480 531.120 1450.740 531.380 ;
        RECT 1449.100 523.980 1449.360 524.240 ;
        RECT 1450.480 523.980 1450.740 524.240 ;
        RECT 1450.020 434.220 1450.280 434.480 ;
        RECT 1450.480 403.620 1450.740 403.880 ;
        RECT 1449.100 310.460 1449.360 310.720 ;
        RECT 1450.020 310.460 1450.280 310.720 ;
        RECT 1449.100 294.820 1449.360 295.080 ;
        RECT 1450.020 294.820 1450.280 295.080 ;
        RECT 1449.100 241.440 1449.360 241.700 ;
        RECT 1450.020 241.440 1450.280 241.700 ;
        RECT 1450.020 144.540 1450.280 144.800 ;
        RECT 1450.480 96.600 1450.740 96.860 ;
        RECT 1450.480 62.260 1450.740 62.520 ;
        RECT 1450.020 61.920 1450.280 62.180 ;
        RECT 1450.020 47.980 1450.280 48.240 ;
        RECT 1108.700 42.200 1108.960 42.460 ;
      LAYER met2 ;
        RECT 1449.090 1700.000 1449.370 1704.000 ;
        RECT 1449.160 1656.470 1449.300 1700.000 ;
        RECT 1449.100 1656.150 1449.360 1656.470 ;
        RECT 1450.020 1656.150 1450.280 1656.470 ;
        RECT 1450.080 1635.390 1450.220 1656.150 ;
        RECT 1450.020 1635.070 1450.280 1635.390 ;
        RECT 1451.860 1607.530 1452.120 1607.850 ;
        RECT 1451.920 1562.970 1452.060 1607.530 ;
        RECT 1451.860 1562.650 1452.120 1562.970 ;
        RECT 1450.020 1400.810 1450.280 1401.130 ;
        RECT 1450.080 1393.845 1450.220 1400.810 ;
        RECT 1450.010 1393.475 1450.290 1393.845 ;
        RECT 1449.090 1345.195 1449.370 1345.565 ;
        RECT 1449.160 1297.430 1449.300 1345.195 ;
        RECT 1449.100 1297.110 1449.360 1297.430 ;
        RECT 1450.020 1297.285 1450.280 1297.430 ;
        RECT 1450.010 1296.915 1450.290 1297.285 ;
        RECT 1450.470 1296.235 1450.750 1296.605 ;
        RECT 1450.540 1249.150 1450.680 1296.235 ;
        RECT 1450.020 1248.830 1450.280 1249.150 ;
        RECT 1450.480 1248.830 1450.740 1249.150 ;
        RECT 1450.080 1200.190 1450.220 1248.830 ;
        RECT 1450.020 1199.870 1450.280 1200.190 ;
        RECT 1450.020 1158.730 1450.280 1159.050 ;
        RECT 1450.080 1128.450 1450.220 1158.730 ;
        RECT 1450.020 1128.130 1450.280 1128.450 ;
        RECT 1450.480 1062.685 1450.740 1062.830 ;
        RECT 1449.090 1062.315 1449.370 1062.685 ;
        RECT 1450.470 1062.315 1450.750 1062.685 ;
        RECT 1449.160 1014.550 1449.300 1062.315 ;
        RECT 1449.100 1014.230 1449.360 1014.550 ;
        RECT 1450.020 1014.405 1450.280 1014.550 ;
        RECT 1450.010 1014.035 1450.290 1014.405 ;
        RECT 1449.090 965.755 1449.370 966.125 ;
        RECT 1449.160 917.990 1449.300 965.755 ;
        RECT 1450.080 917.990 1450.220 918.145 ;
        RECT 1449.100 917.670 1449.360 917.990 ;
        RECT 1450.020 917.730 1450.280 917.990 ;
        RECT 1450.020 917.670 1450.680 917.730 ;
        RECT 1450.080 917.650 1450.680 917.670 ;
        RECT 1450.080 917.590 1450.740 917.650 ;
        RECT 1450.480 917.330 1450.740 917.590 ;
        RECT 1450.480 869.730 1450.740 870.050 ;
        RECT 1450.540 869.565 1450.680 869.730 ;
        RECT 1449.090 869.195 1449.370 869.565 ;
        RECT 1450.470 869.195 1450.750 869.565 ;
        RECT 1449.160 821.285 1449.300 869.195 ;
        RECT 1449.090 820.915 1449.370 821.285 ;
        RECT 1450.010 820.915 1450.290 821.285 ;
        RECT 1450.080 772.890 1450.220 820.915 ;
        RECT 1450.080 772.810 1450.680 772.890 ;
        RECT 1449.100 772.490 1449.360 772.810 ;
        RECT 1450.080 772.750 1450.740 772.810 ;
        RECT 1450.480 772.490 1450.740 772.750 ;
        RECT 1449.160 724.725 1449.300 772.490 ;
        RECT 1450.540 772.335 1450.680 772.490 ;
        RECT 1449.090 724.355 1449.370 724.725 ;
        RECT 1450.010 724.355 1450.290 724.725 ;
        RECT 1450.080 676.930 1450.220 724.355 ;
        RECT 1450.020 676.610 1450.280 676.930 ;
        RECT 1450.020 662.330 1450.280 662.650 ;
        RECT 1450.080 651.430 1450.220 662.330 ;
        RECT 1450.020 651.110 1450.280 651.430 ;
        RECT 1450.020 650.430 1450.280 650.750 ;
        RECT 1450.080 593.970 1450.220 650.430 ;
        RECT 1450.020 593.650 1450.280 593.970 ;
        RECT 1450.020 592.970 1450.280 593.290 ;
        RECT 1450.080 531.410 1450.220 592.970 ;
        RECT 1450.020 531.090 1450.280 531.410 ;
        RECT 1450.480 531.090 1450.740 531.410 ;
        RECT 1450.540 524.270 1450.680 531.090 ;
        RECT 1449.100 523.950 1449.360 524.270 ;
        RECT 1450.480 523.950 1450.740 524.270 ;
        RECT 1449.160 435.045 1449.300 523.950 ;
        RECT 1449.090 434.675 1449.370 435.045 ;
        RECT 1450.010 434.675 1450.290 435.045 ;
        RECT 1450.080 434.510 1450.220 434.675 ;
        RECT 1450.020 434.190 1450.280 434.510 ;
        RECT 1450.480 403.590 1450.740 403.910 ;
        RECT 1450.540 358.885 1450.680 403.590 ;
        RECT 1449.090 358.515 1449.370 358.885 ;
        RECT 1450.470 358.515 1450.750 358.885 ;
        RECT 1449.160 310.750 1449.300 358.515 ;
        RECT 1449.100 310.430 1449.360 310.750 ;
        RECT 1450.020 310.430 1450.280 310.750 ;
        RECT 1450.080 295.110 1450.220 310.430 ;
        RECT 1449.100 294.790 1449.360 295.110 ;
        RECT 1450.020 294.790 1450.280 295.110 ;
        RECT 1449.160 241.730 1449.300 294.790 ;
        RECT 1449.100 241.410 1449.360 241.730 ;
        RECT 1450.020 241.410 1450.280 241.730 ;
        RECT 1450.080 217.330 1450.220 241.410 ;
        RECT 1450.080 217.190 1450.680 217.330 ;
        RECT 1450.540 145.250 1450.680 217.190 ;
        RECT 1450.080 145.110 1450.680 145.250 ;
        RECT 1450.080 144.830 1450.220 145.110 ;
        RECT 1450.020 144.510 1450.280 144.830 ;
        RECT 1450.480 96.570 1450.740 96.890 ;
        RECT 1450.540 62.550 1450.680 96.570 ;
        RECT 1450.480 62.230 1450.740 62.550 ;
        RECT 1450.020 61.890 1450.280 62.210 ;
        RECT 1450.080 48.270 1450.220 61.890 ;
        RECT 1450.020 47.950 1450.280 48.270 ;
        RECT 1108.700 42.170 1108.960 42.490 ;
        RECT 1108.760 2.400 1108.900 42.170 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
      LAYER via2 ;
        RECT 1450.010 1393.520 1450.290 1393.800 ;
        RECT 1449.090 1345.240 1449.370 1345.520 ;
        RECT 1450.010 1296.960 1450.290 1297.240 ;
        RECT 1450.470 1296.280 1450.750 1296.560 ;
        RECT 1449.090 1062.360 1449.370 1062.640 ;
        RECT 1450.470 1062.360 1450.750 1062.640 ;
        RECT 1450.010 1014.080 1450.290 1014.360 ;
        RECT 1449.090 965.800 1449.370 966.080 ;
        RECT 1449.090 869.240 1449.370 869.520 ;
        RECT 1450.470 869.240 1450.750 869.520 ;
        RECT 1449.090 820.960 1449.370 821.240 ;
        RECT 1450.010 820.960 1450.290 821.240 ;
        RECT 1449.090 724.400 1449.370 724.680 ;
        RECT 1450.010 724.400 1450.290 724.680 ;
        RECT 1449.090 434.720 1449.370 435.000 ;
        RECT 1450.010 434.720 1450.290 435.000 ;
        RECT 1449.090 358.560 1449.370 358.840 ;
        RECT 1450.470 358.560 1450.750 358.840 ;
      LAYER met3 ;
        RECT 1449.985 1393.810 1450.315 1393.825 ;
        RECT 1451.110 1393.810 1451.490 1393.820 ;
        RECT 1449.985 1393.510 1451.490 1393.810 ;
        RECT 1449.985 1393.495 1450.315 1393.510 ;
        RECT 1451.110 1393.500 1451.490 1393.510 ;
        RECT 1451.110 1345.900 1451.490 1346.220 ;
        RECT 1449.065 1345.530 1449.395 1345.545 ;
        RECT 1451.150 1345.530 1451.450 1345.900 ;
        RECT 1449.065 1345.230 1451.450 1345.530 ;
        RECT 1449.065 1345.215 1449.395 1345.230 ;
        RECT 1449.985 1297.250 1450.315 1297.265 ;
        RECT 1449.985 1296.935 1450.530 1297.250 ;
        RECT 1450.230 1296.585 1450.530 1296.935 ;
        RECT 1450.230 1296.270 1450.775 1296.585 ;
        RECT 1450.445 1296.255 1450.775 1296.270 ;
        RECT 1449.065 1062.650 1449.395 1062.665 ;
        RECT 1450.445 1062.650 1450.775 1062.665 ;
        RECT 1449.065 1062.350 1450.775 1062.650 ;
        RECT 1449.065 1062.335 1449.395 1062.350 ;
        RECT 1450.445 1062.335 1450.775 1062.350 ;
        RECT 1449.985 1014.380 1450.315 1014.385 ;
        RECT 1449.985 1014.370 1450.570 1014.380 ;
        RECT 1449.760 1014.070 1450.570 1014.370 ;
        RECT 1449.985 1014.060 1450.570 1014.070 ;
        RECT 1449.985 1014.055 1450.315 1014.060 ;
        RECT 1450.190 967.450 1450.570 967.460 ;
        RECT 1450.190 967.150 1451.450 967.450 ;
        RECT 1450.190 967.140 1450.570 967.150 ;
        RECT 1449.065 966.090 1449.395 966.105 ;
        RECT 1451.150 966.090 1451.450 967.150 ;
        RECT 1449.065 965.790 1451.450 966.090 ;
        RECT 1449.065 965.775 1449.395 965.790 ;
        RECT 1449.065 869.530 1449.395 869.545 ;
        RECT 1450.445 869.530 1450.775 869.545 ;
        RECT 1449.065 869.230 1450.775 869.530 ;
        RECT 1449.065 869.215 1449.395 869.230 ;
        RECT 1450.445 869.215 1450.775 869.230 ;
        RECT 1449.065 821.250 1449.395 821.265 ;
        RECT 1449.985 821.250 1450.315 821.265 ;
        RECT 1449.065 820.950 1450.315 821.250 ;
        RECT 1449.065 820.935 1449.395 820.950 ;
        RECT 1449.985 820.935 1450.315 820.950 ;
        RECT 1449.065 724.690 1449.395 724.705 ;
        RECT 1449.985 724.690 1450.315 724.705 ;
        RECT 1449.065 724.390 1450.315 724.690 ;
        RECT 1449.065 724.375 1449.395 724.390 ;
        RECT 1449.985 724.375 1450.315 724.390 ;
        RECT 1449.065 435.010 1449.395 435.025 ;
        RECT 1449.985 435.010 1450.315 435.025 ;
        RECT 1449.065 434.710 1450.315 435.010 ;
        RECT 1449.065 434.695 1449.395 434.710 ;
        RECT 1449.985 434.695 1450.315 434.710 ;
        RECT 1449.065 358.850 1449.395 358.865 ;
        RECT 1450.445 358.850 1450.775 358.865 ;
        RECT 1449.065 358.550 1450.775 358.850 ;
        RECT 1449.065 358.535 1449.395 358.550 ;
        RECT 1450.445 358.535 1450.775 358.550 ;
      LAYER via3 ;
        RECT 1451.140 1393.500 1451.460 1393.820 ;
        RECT 1451.140 1345.900 1451.460 1346.220 ;
        RECT 1450.220 1014.060 1450.540 1014.380 ;
        RECT 1450.220 967.140 1450.540 967.460 ;
      LAYER met4 ;
        RECT 1451.135 1393.495 1451.465 1393.825 ;
        RECT 1451.150 1346.225 1451.450 1393.495 ;
        RECT 1451.135 1345.895 1451.465 1346.225 ;
        RECT 1450.215 1014.055 1450.545 1014.385 ;
        RECT 1450.230 967.465 1450.530 1014.055 ;
        RECT 1450.215 967.135 1450.545 967.465 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 0.300 ;
=======
      LAYER li1 ;
        RECT 1452.365 1545.045 1452.535 1635.315 ;
        RECT 1451.905 965.005 1452.075 1007.335 ;
        RECT 1451.905 917.745 1452.075 931.855 ;
        RECT 1451.905 379.525 1452.075 434.435 ;
        RECT 1451.905 41.905 1452.075 48.195 ;
      LAYER mcon ;
        RECT 1452.365 1635.145 1452.535 1635.315 ;
        RECT 1451.905 1007.165 1452.075 1007.335 ;
        RECT 1451.905 931.685 1452.075 931.855 ;
        RECT 1451.905 434.265 1452.075 434.435 ;
        RECT 1451.905 48.025 1452.075 48.195 ;
      LAYER met1 ;
        RECT 1451.830 1635.300 1452.150 1635.360 ;
        RECT 1452.305 1635.300 1452.595 1635.345 ;
        RECT 1451.830 1635.160 1452.595 1635.300 ;
        RECT 1451.830 1635.100 1452.150 1635.160 ;
        RECT 1452.305 1635.115 1452.595 1635.160 ;
        RECT 1452.305 1545.200 1452.595 1545.245 ;
        RECT 1452.750 1545.200 1453.070 1545.260 ;
        RECT 1452.305 1545.060 1453.070 1545.200 ;
        RECT 1452.305 1545.015 1452.595 1545.060 ;
        RECT 1452.750 1545.000 1453.070 1545.060 ;
        RECT 1452.750 1490.260 1453.070 1490.520 ;
        RECT 1452.840 1489.840 1452.980 1490.260 ;
        RECT 1452.750 1489.580 1453.070 1489.840 ;
        RECT 1451.830 1393.900 1452.150 1393.960 ;
        RECT 1452.750 1393.900 1453.070 1393.960 ;
        RECT 1451.830 1393.760 1453.070 1393.900 ;
        RECT 1451.830 1393.700 1452.150 1393.760 ;
        RECT 1452.750 1393.700 1453.070 1393.760 ;
        RECT 1451.830 1345.620 1452.150 1345.680 ;
        RECT 1453.210 1345.620 1453.530 1345.680 ;
        RECT 1451.830 1345.480 1453.530 1345.620 ;
        RECT 1451.830 1345.420 1452.150 1345.480 ;
        RECT 1453.210 1345.420 1453.530 1345.480 ;
        RECT 1451.830 1297.340 1452.150 1297.400 ;
        RECT 1452.750 1297.340 1453.070 1297.400 ;
        RECT 1451.830 1297.200 1453.070 1297.340 ;
        RECT 1451.830 1297.140 1452.150 1297.200 ;
        RECT 1452.750 1297.140 1453.070 1297.200 ;
        RECT 1451.830 1269.600 1452.150 1269.860 ;
        RECT 1451.920 1269.460 1452.060 1269.600 ;
        RECT 1452.290 1269.460 1452.610 1269.520 ;
        RECT 1451.920 1269.320 1452.610 1269.460 ;
        RECT 1452.290 1269.260 1452.610 1269.320 ;
        RECT 1451.830 1152.500 1452.150 1152.560 ;
        RECT 1452.750 1152.500 1453.070 1152.560 ;
        RECT 1451.830 1152.360 1453.070 1152.500 ;
        RECT 1451.830 1152.300 1452.150 1152.360 ;
        RECT 1452.750 1152.300 1453.070 1152.360 ;
        RECT 1451.830 1007.320 1452.150 1007.380 ;
        RECT 1451.635 1007.180 1452.150 1007.320 ;
        RECT 1451.830 1007.120 1452.150 1007.180 ;
        RECT 1451.830 965.160 1452.150 965.220 ;
        RECT 1451.635 965.020 1452.150 965.160 ;
        RECT 1451.830 964.960 1452.150 965.020 ;
        RECT 1451.830 931.840 1452.150 931.900 ;
        RECT 1451.635 931.700 1452.150 931.840 ;
        RECT 1451.830 931.640 1452.150 931.700 ;
        RECT 1451.830 917.900 1452.150 917.960 ;
        RECT 1451.635 917.760 1452.150 917.900 ;
        RECT 1451.830 917.700 1452.150 917.760 ;
        RECT 1451.830 910.760 1452.150 910.820 ;
        RECT 1453.210 910.760 1453.530 910.820 ;
        RECT 1451.830 910.620 1453.530 910.760 ;
        RECT 1451.830 910.560 1452.150 910.620 ;
        RECT 1453.210 910.560 1453.530 910.620 ;
        RECT 1452.290 820.800 1452.610 821.060 ;
        RECT 1452.380 820.380 1452.520 820.800 ;
        RECT 1452.290 820.120 1452.610 820.380 ;
        RECT 1452.290 765.920 1452.610 765.980 ;
        RECT 1453.210 765.920 1453.530 765.980 ;
        RECT 1452.290 765.780 1453.530 765.920 ;
        RECT 1452.290 765.720 1452.610 765.780 ;
        RECT 1453.210 765.720 1453.530 765.780 ;
        RECT 1451.830 593.340 1452.150 593.600 ;
        RECT 1451.920 593.200 1452.060 593.340 ;
        RECT 1452.290 593.200 1452.610 593.260 ;
        RECT 1451.920 593.060 1452.610 593.200 ;
        RECT 1452.290 593.000 1452.610 593.060 ;
        RECT 1452.290 449.040 1452.610 449.100 ;
        RECT 1451.920 448.900 1452.610 449.040 ;
        RECT 1451.920 448.420 1452.060 448.900 ;
        RECT 1452.290 448.840 1452.610 448.900 ;
        RECT 1451.830 448.160 1452.150 448.420 ;
        RECT 1451.830 434.420 1452.150 434.480 ;
        RECT 1451.635 434.280 1452.150 434.420 ;
        RECT 1451.830 434.220 1452.150 434.280 ;
        RECT 1451.845 379.680 1452.135 379.725 ;
        RECT 1452.290 379.680 1452.610 379.740 ;
        RECT 1451.845 379.540 1452.610 379.680 ;
        RECT 1451.845 379.495 1452.135 379.540 ;
        RECT 1452.290 379.480 1452.610 379.540 ;
        RECT 1451.830 303.520 1452.150 303.580 ;
        RECT 1453.210 303.520 1453.530 303.580 ;
        RECT 1451.830 303.380 1453.530 303.520 ;
        RECT 1451.830 303.320 1452.150 303.380 ;
        RECT 1453.210 303.320 1453.530 303.380 ;
        RECT 1451.830 214.100 1452.150 214.160 ;
        RECT 1452.290 214.100 1452.610 214.160 ;
        RECT 1451.830 213.960 1452.610 214.100 ;
        RECT 1451.830 213.900 1452.150 213.960 ;
        RECT 1452.290 213.900 1452.610 213.960 ;
        RECT 1451.830 193.360 1452.150 193.420 ;
        RECT 1452.290 193.360 1452.610 193.420 ;
        RECT 1451.830 193.220 1452.610 193.360 ;
        RECT 1451.830 193.160 1452.150 193.220 ;
        RECT 1452.290 193.160 1452.610 193.220 ;
        RECT 1452.290 96.800 1452.610 96.860 ;
        RECT 1452.750 96.800 1453.070 96.860 ;
        RECT 1452.290 96.660 1453.070 96.800 ;
        RECT 1452.290 96.600 1452.610 96.660 ;
        RECT 1452.750 96.600 1453.070 96.660 ;
        RECT 1451.830 48.180 1452.150 48.240 ;
        RECT 1451.635 48.040 1452.150 48.180 ;
        RECT 1451.830 47.980 1452.150 48.040 ;
        RECT 1126.610 42.060 1126.930 42.120 ;
        RECT 1451.845 42.060 1452.135 42.105 ;
        RECT 1126.610 41.920 1452.135 42.060 ;
        RECT 1126.610 41.860 1126.930 41.920 ;
        RECT 1451.845 41.875 1452.135 41.920 ;
      LAYER via ;
        RECT 1451.860 1635.100 1452.120 1635.360 ;
        RECT 1452.780 1545.000 1453.040 1545.260 ;
        RECT 1452.780 1490.260 1453.040 1490.520 ;
        RECT 1452.780 1489.580 1453.040 1489.840 ;
        RECT 1451.860 1393.700 1452.120 1393.960 ;
        RECT 1452.780 1393.700 1453.040 1393.960 ;
        RECT 1451.860 1345.420 1452.120 1345.680 ;
        RECT 1453.240 1345.420 1453.500 1345.680 ;
        RECT 1451.860 1297.140 1452.120 1297.400 ;
        RECT 1452.780 1297.140 1453.040 1297.400 ;
        RECT 1451.860 1269.600 1452.120 1269.860 ;
        RECT 1452.320 1269.260 1452.580 1269.520 ;
        RECT 1451.860 1152.300 1452.120 1152.560 ;
        RECT 1452.780 1152.300 1453.040 1152.560 ;
        RECT 1451.860 1007.120 1452.120 1007.380 ;
        RECT 1451.860 964.960 1452.120 965.220 ;
        RECT 1451.860 931.640 1452.120 931.900 ;
        RECT 1451.860 917.700 1452.120 917.960 ;
        RECT 1451.860 910.560 1452.120 910.820 ;
        RECT 1453.240 910.560 1453.500 910.820 ;
        RECT 1452.320 820.800 1452.580 821.060 ;
        RECT 1452.320 820.120 1452.580 820.380 ;
        RECT 1452.320 765.720 1452.580 765.980 ;
        RECT 1453.240 765.720 1453.500 765.980 ;
        RECT 1451.860 593.340 1452.120 593.600 ;
        RECT 1452.320 593.000 1452.580 593.260 ;
        RECT 1452.320 448.840 1452.580 449.100 ;
        RECT 1451.860 448.160 1452.120 448.420 ;
        RECT 1451.860 434.220 1452.120 434.480 ;
        RECT 1452.320 379.480 1452.580 379.740 ;
        RECT 1451.860 303.320 1452.120 303.580 ;
        RECT 1453.240 303.320 1453.500 303.580 ;
        RECT 1451.860 213.900 1452.120 214.160 ;
        RECT 1452.320 213.900 1452.580 214.160 ;
        RECT 1451.860 193.160 1452.120 193.420 ;
        RECT 1452.320 193.160 1452.580 193.420 ;
        RECT 1452.320 96.600 1452.580 96.860 ;
        RECT 1452.780 96.600 1453.040 96.860 ;
        RECT 1451.860 47.980 1452.120 48.240 ;
        RECT 1126.640 41.860 1126.900 42.120 ;
      LAYER met2 ;
        RECT 1453.690 1700.410 1453.970 1704.000 ;
        RECT 1453.300 1700.270 1453.970 1700.410 ;
        RECT 1453.300 1656.210 1453.440 1700.270 ;
        RECT 1453.690 1700.000 1453.970 1700.270 ;
        RECT 1451.920 1656.070 1453.440 1656.210 ;
        RECT 1451.920 1635.390 1452.060 1656.070 ;
        RECT 1451.860 1635.070 1452.120 1635.390 ;
        RECT 1452.780 1544.970 1453.040 1545.290 ;
        RECT 1452.840 1490.550 1452.980 1544.970 ;
        RECT 1452.780 1490.230 1453.040 1490.550 ;
        RECT 1452.780 1489.550 1453.040 1489.870 ;
        RECT 1452.840 1393.990 1452.980 1489.550 ;
        RECT 1451.860 1393.845 1452.120 1393.990 ;
        RECT 1451.850 1393.475 1452.130 1393.845 ;
        RECT 1452.780 1393.670 1453.040 1393.990 ;
        RECT 1453.230 1393.475 1453.510 1393.845 ;
        RECT 1453.300 1345.710 1453.440 1393.475 ;
        RECT 1451.860 1345.565 1452.120 1345.710 ;
        RECT 1451.850 1345.195 1452.130 1345.565 ;
        RECT 1452.770 1345.195 1453.050 1345.565 ;
        RECT 1453.240 1345.390 1453.500 1345.710 ;
        RECT 1452.840 1297.430 1452.980 1345.195 ;
        RECT 1451.860 1297.110 1452.120 1297.430 ;
        RECT 1452.780 1297.110 1453.040 1297.430 ;
        RECT 1451.920 1269.890 1452.060 1297.110 ;
        RECT 1451.860 1269.570 1452.120 1269.890 ;
        RECT 1452.320 1269.230 1452.580 1269.550 ;
        RECT 1452.380 1231.890 1452.520 1269.230 ;
        RECT 1452.380 1231.750 1452.980 1231.890 ;
        RECT 1452.840 1152.590 1452.980 1231.750 ;
        RECT 1451.860 1152.270 1452.120 1152.590 ;
        RECT 1452.780 1152.270 1453.040 1152.590 ;
        RECT 1451.920 1110.965 1452.060 1152.270 ;
        RECT 1451.850 1110.595 1452.130 1110.965 ;
        RECT 1453.230 1110.595 1453.510 1110.965 ;
        RECT 1453.300 1049.650 1453.440 1110.595 ;
        RECT 1452.840 1049.510 1453.440 1049.650 ;
        RECT 1452.840 1049.085 1452.980 1049.510 ;
        RECT 1451.850 1048.715 1452.130 1049.085 ;
        RECT 1452.770 1048.715 1453.050 1049.085 ;
        RECT 1451.920 1007.410 1452.060 1048.715 ;
        RECT 1451.860 1007.090 1452.120 1007.410 ;
        RECT 1451.860 964.930 1452.120 965.250 ;
        RECT 1451.920 931.930 1452.060 964.930 ;
        RECT 1451.860 931.610 1452.120 931.930 ;
        RECT 1451.860 917.670 1452.120 917.990 ;
        RECT 1451.920 910.850 1452.060 917.670 ;
        RECT 1451.860 910.530 1452.120 910.850 ;
        RECT 1453.240 910.530 1453.500 910.850 ;
        RECT 1453.300 862.765 1453.440 910.530 ;
        RECT 1452.310 862.395 1452.590 862.765 ;
        RECT 1453.230 862.395 1453.510 862.765 ;
        RECT 1452.380 821.090 1452.520 862.395 ;
        RECT 1452.320 820.770 1452.580 821.090 ;
        RECT 1452.320 820.090 1452.580 820.410 ;
        RECT 1452.380 766.010 1452.520 820.090 ;
        RECT 1452.320 765.690 1452.580 766.010 ;
        RECT 1453.240 765.690 1453.500 766.010 ;
        RECT 1453.300 717.925 1453.440 765.690 ;
        RECT 1451.850 717.555 1452.130 717.925 ;
        RECT 1453.230 717.555 1453.510 717.925 ;
        RECT 1451.920 593.630 1452.060 717.555 ;
        RECT 1451.860 593.310 1452.120 593.630 ;
        RECT 1452.320 592.970 1452.580 593.290 ;
        RECT 1452.380 548.490 1452.520 592.970 ;
        RECT 1452.380 548.350 1453.440 548.490 ;
        RECT 1453.300 494.090 1453.440 548.350 ;
        RECT 1452.840 493.950 1453.440 494.090 ;
        RECT 1452.840 483.210 1452.980 493.950 ;
        RECT 1452.380 483.070 1452.980 483.210 ;
        RECT 1452.380 449.130 1452.520 483.070 ;
        RECT 1452.320 448.810 1452.580 449.130 ;
        RECT 1451.860 448.130 1452.120 448.450 ;
        RECT 1451.920 434.510 1452.060 448.130 ;
        RECT 1451.860 434.190 1452.120 434.510 ;
        RECT 1452.320 379.450 1452.580 379.770 ;
        RECT 1452.380 311.170 1452.520 379.450 ;
        RECT 1451.920 311.030 1452.520 311.170 ;
        RECT 1451.920 303.610 1452.060 311.030 ;
        RECT 1451.860 303.290 1452.120 303.610 ;
        RECT 1453.240 303.290 1453.500 303.610 ;
        RECT 1453.300 255.525 1453.440 303.290 ;
        RECT 1452.310 255.155 1452.590 255.525 ;
        RECT 1453.230 255.155 1453.510 255.525 ;
        RECT 1452.380 214.190 1452.520 255.155 ;
        RECT 1451.860 213.870 1452.120 214.190 ;
        RECT 1452.320 213.870 1452.580 214.190 ;
        RECT 1451.920 193.450 1452.060 213.870 ;
        RECT 1451.860 193.130 1452.120 193.450 ;
        RECT 1452.320 193.130 1452.580 193.450 ;
        RECT 1452.380 145.365 1452.520 193.130 ;
        RECT 1452.310 144.995 1452.590 145.365 ;
        RECT 1452.770 143.635 1453.050 144.005 ;
        RECT 1452.840 96.890 1452.980 143.635 ;
        RECT 1452.320 96.570 1452.580 96.890 ;
        RECT 1452.780 96.570 1453.040 96.890 ;
        RECT 1452.380 62.970 1452.520 96.570 ;
        RECT 1452.380 62.830 1452.980 62.970 ;
        RECT 1452.840 48.690 1452.980 62.830 ;
        RECT 1451.920 48.550 1452.980 48.690 ;
        RECT 1451.920 48.270 1452.060 48.550 ;
        RECT 1451.860 47.950 1452.120 48.270 ;
        RECT 1126.640 41.830 1126.900 42.150 ;
        RECT 1126.700 2.400 1126.840 41.830 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
      LAYER via2 ;
        RECT 1451.850 1393.520 1452.130 1393.800 ;
        RECT 1453.230 1393.520 1453.510 1393.800 ;
        RECT 1451.850 1345.240 1452.130 1345.520 ;
        RECT 1452.770 1345.240 1453.050 1345.520 ;
        RECT 1451.850 1110.640 1452.130 1110.920 ;
        RECT 1453.230 1110.640 1453.510 1110.920 ;
        RECT 1451.850 1048.760 1452.130 1049.040 ;
        RECT 1452.770 1048.760 1453.050 1049.040 ;
        RECT 1452.310 862.440 1452.590 862.720 ;
        RECT 1453.230 862.440 1453.510 862.720 ;
        RECT 1451.850 717.600 1452.130 717.880 ;
        RECT 1453.230 717.600 1453.510 717.880 ;
        RECT 1452.310 255.200 1452.590 255.480 ;
        RECT 1453.230 255.200 1453.510 255.480 ;
        RECT 1452.310 145.040 1452.590 145.320 ;
        RECT 1452.770 143.680 1453.050 143.960 ;
      LAYER met3 ;
        RECT 1451.825 1393.810 1452.155 1393.825 ;
        RECT 1453.205 1393.810 1453.535 1393.825 ;
        RECT 1451.825 1393.510 1453.535 1393.810 ;
        RECT 1451.825 1393.495 1452.155 1393.510 ;
        RECT 1453.205 1393.495 1453.535 1393.510 ;
        RECT 1451.825 1345.530 1452.155 1345.545 ;
        RECT 1452.745 1345.530 1453.075 1345.545 ;
        RECT 1451.825 1345.230 1453.075 1345.530 ;
        RECT 1451.825 1345.215 1452.155 1345.230 ;
        RECT 1452.745 1345.215 1453.075 1345.230 ;
        RECT 1451.825 1110.930 1452.155 1110.945 ;
        RECT 1453.205 1110.930 1453.535 1110.945 ;
        RECT 1451.825 1110.630 1453.535 1110.930 ;
        RECT 1451.825 1110.615 1452.155 1110.630 ;
        RECT 1453.205 1110.615 1453.535 1110.630 ;
        RECT 1451.825 1049.050 1452.155 1049.065 ;
        RECT 1452.745 1049.050 1453.075 1049.065 ;
        RECT 1451.825 1048.750 1453.075 1049.050 ;
        RECT 1451.825 1048.735 1452.155 1048.750 ;
        RECT 1452.745 1048.735 1453.075 1048.750 ;
        RECT 1452.285 862.730 1452.615 862.745 ;
        RECT 1453.205 862.730 1453.535 862.745 ;
        RECT 1452.285 862.430 1453.535 862.730 ;
        RECT 1452.285 862.415 1452.615 862.430 ;
        RECT 1453.205 862.415 1453.535 862.430 ;
        RECT 1451.825 717.890 1452.155 717.905 ;
        RECT 1453.205 717.890 1453.535 717.905 ;
        RECT 1451.825 717.590 1453.535 717.890 ;
        RECT 1451.825 717.575 1452.155 717.590 ;
        RECT 1453.205 717.575 1453.535 717.590 ;
        RECT 1452.285 255.490 1452.615 255.505 ;
        RECT 1453.205 255.490 1453.535 255.505 ;
        RECT 1452.285 255.190 1453.535 255.490 ;
        RECT 1452.285 255.175 1452.615 255.190 ;
        RECT 1453.205 255.175 1453.535 255.190 ;
        RECT 1452.285 145.330 1452.615 145.345 ;
        RECT 1451.150 145.030 1452.615 145.330 ;
        RECT 1451.150 143.970 1451.450 145.030 ;
        RECT 1452.285 145.015 1452.615 145.030 ;
        RECT 1452.745 143.970 1453.075 143.985 ;
        RECT 1451.150 143.670 1453.075 143.970 ;
        RECT 1452.745 143.655 1453.075 143.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1144.550 41.720 1144.870 41.780 ;
        RECT 1457.810 41.720 1458.130 41.780 ;
        RECT 1144.550 41.580 1458.130 41.720 ;
        RECT 1144.550 41.520 1144.870 41.580 ;
        RECT 1457.810 41.520 1458.130 41.580 ;
      LAYER via ;
        RECT 1144.580 41.520 1144.840 41.780 ;
        RECT 1457.840 41.520 1458.100 41.780 ;
      LAYER met2 ;
        RECT 1458.750 1700.410 1459.030 1704.000 ;
        RECT 1457.900 1700.270 1459.030 1700.410 ;
        RECT 1457.900 41.810 1458.040 1700.270 ;
        RECT 1458.750 1700.000 1459.030 1700.270 ;
        RECT 1144.580 41.490 1144.840 41.810 ;
        RECT 1457.840 41.490 1458.100 41.810 ;
        RECT 1144.640 2.400 1144.780 41.490 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1162.490 24.380 1162.810 24.440 ;
        RECT 1463.790 24.380 1464.110 24.440 ;
        RECT 1162.490 24.240 1464.110 24.380 ;
        RECT 1162.490 24.180 1162.810 24.240 ;
        RECT 1463.790 24.180 1464.110 24.240 ;
      LAYER via ;
        RECT 1162.520 24.180 1162.780 24.440 ;
        RECT 1463.820 24.180 1464.080 24.440 ;
      LAYER met2 ;
        RECT 1463.350 1700.410 1463.630 1704.000 ;
        RECT 1463.350 1700.270 1464.020 1700.410 ;
        RECT 1463.350 1700.000 1463.630 1700.270 ;
        RECT 1463.880 24.470 1464.020 1700.270 ;
        RECT 1162.520 24.150 1162.780 24.470 ;
        RECT 1463.820 24.150 1464.080 24.470 ;
        RECT 1162.580 2.400 1162.720 24.150 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 0.300 ;
=======
      LAYER met1 ;
        RECT 680.410 46.480 680.730 46.540 ;
        RECT 1332.690 46.480 1333.010 46.540 ;
        RECT 680.410 46.340 1333.010 46.480 ;
        RECT 680.410 46.280 680.730 46.340 ;
        RECT 1332.690 46.280 1333.010 46.340 ;
      LAYER via ;
        RECT 680.440 46.280 680.700 46.540 ;
        RECT 1332.720 46.280 1332.980 46.540 ;
      LAYER met2 ;
        RECT 1333.630 1700.410 1333.910 1704.000 ;
        RECT 1332.780 1700.270 1333.910 1700.410 ;
        RECT 1332.780 46.570 1332.920 1700.270 ;
        RECT 1333.630 1700.000 1333.910 1700.270 ;
        RECT 680.440 46.250 680.700 46.570 ;
        RECT 1332.720 46.250 1332.980 46.570 ;
        RECT 680.500 2.400 680.640 46.250 ;
        RECT 680.290 -4.800 680.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 0.300 ;
=======
      LAYER li1 ;
        RECT 1465.245 386.325 1465.415 410.635 ;
      LAYER mcon ;
        RECT 1465.245 410.465 1465.415 410.635 ;
      LAYER met1 ;
        RECT 1464.710 1607.900 1465.030 1608.160 ;
        RECT 1464.800 1607.480 1464.940 1607.900 ;
        RECT 1464.710 1607.220 1465.030 1607.480 ;
        RECT 1464.710 1497.060 1465.030 1497.320 ;
        RECT 1464.800 1496.920 1464.940 1497.060 ;
        RECT 1465.630 1496.920 1465.950 1496.980 ;
        RECT 1464.800 1496.780 1465.950 1496.920 ;
        RECT 1465.630 1496.720 1465.950 1496.780 ;
        RECT 1465.170 1111.020 1465.490 1111.080 ;
        RECT 1466.090 1111.020 1466.410 1111.080 ;
        RECT 1465.170 1110.880 1466.410 1111.020 ;
        RECT 1465.170 1110.820 1465.490 1110.880 ;
        RECT 1466.090 1110.820 1466.410 1110.880 ;
        RECT 1465.170 869.620 1465.490 869.680 ;
        RECT 1465.630 869.620 1465.950 869.680 ;
        RECT 1465.170 869.480 1465.950 869.620 ;
        RECT 1465.170 869.420 1465.490 869.480 ;
        RECT 1465.630 869.420 1465.950 869.480 ;
        RECT 1465.185 410.620 1465.475 410.665 ;
        RECT 1465.630 410.620 1465.950 410.680 ;
        RECT 1465.185 410.480 1465.950 410.620 ;
        RECT 1465.185 410.435 1465.475 410.480 ;
        RECT 1465.630 410.420 1465.950 410.480 ;
        RECT 1465.170 386.480 1465.490 386.540 ;
        RECT 1464.975 386.340 1465.490 386.480 ;
        RECT 1465.170 386.280 1465.490 386.340 ;
        RECT 1179.970 17.240 1180.290 17.300 ;
        RECT 1465.170 17.240 1465.490 17.300 ;
        RECT 1179.970 17.100 1465.490 17.240 ;
        RECT 1179.970 17.040 1180.290 17.100 ;
        RECT 1465.170 17.040 1465.490 17.100 ;
      LAYER via ;
        RECT 1464.740 1607.900 1465.000 1608.160 ;
        RECT 1464.740 1607.220 1465.000 1607.480 ;
        RECT 1464.740 1497.060 1465.000 1497.320 ;
        RECT 1465.660 1496.720 1465.920 1496.980 ;
        RECT 1465.200 1110.820 1465.460 1111.080 ;
        RECT 1466.120 1110.820 1466.380 1111.080 ;
        RECT 1465.200 869.420 1465.460 869.680 ;
        RECT 1465.660 869.420 1465.920 869.680 ;
        RECT 1465.660 410.420 1465.920 410.680 ;
        RECT 1465.200 386.280 1465.460 386.540 ;
        RECT 1180.000 17.040 1180.260 17.300 ;
        RECT 1465.200 17.040 1465.460 17.300 ;
      LAYER met2 ;
        RECT 1468.410 1700.410 1468.690 1704.000 ;
        RECT 1467.560 1700.270 1468.690 1700.410 ;
        RECT 1467.560 1677.290 1467.700 1700.270 ;
        RECT 1468.410 1700.000 1468.690 1700.270 ;
        RECT 1464.800 1677.150 1467.700 1677.290 ;
        RECT 1464.800 1608.190 1464.940 1677.150 ;
        RECT 1464.740 1607.870 1465.000 1608.190 ;
        RECT 1464.740 1607.190 1465.000 1607.510 ;
        RECT 1464.800 1497.350 1464.940 1607.190 ;
        RECT 1464.740 1497.030 1465.000 1497.350 ;
        RECT 1465.660 1496.690 1465.920 1497.010 ;
        RECT 1465.720 1366.530 1465.860 1496.690 ;
        RECT 1464.800 1366.390 1465.860 1366.530 ;
        RECT 1464.800 1365.850 1464.940 1366.390 ;
        RECT 1464.800 1365.710 1465.400 1365.850 ;
        RECT 1465.260 1297.170 1465.400 1365.710 ;
        RECT 1465.260 1297.030 1465.860 1297.170 ;
        RECT 1465.720 1207.410 1465.860 1297.030 ;
        RECT 1465.720 1207.270 1466.320 1207.410 ;
        RECT 1466.180 1200.725 1466.320 1207.270 ;
        RECT 1465.190 1200.355 1465.470 1200.725 ;
        RECT 1466.110 1200.355 1466.390 1200.725 ;
        RECT 1465.260 1157.770 1465.400 1200.355 ;
        RECT 1465.260 1157.630 1466.320 1157.770 ;
        RECT 1466.180 1111.110 1466.320 1157.630 ;
        RECT 1465.200 1110.790 1465.460 1111.110 ;
        RECT 1466.120 1110.790 1466.380 1111.110 ;
        RECT 1465.260 1014.290 1465.400 1110.790 ;
        RECT 1465.260 1014.150 1465.860 1014.290 ;
        RECT 1465.720 869.710 1465.860 1014.150 ;
        RECT 1465.200 869.390 1465.460 869.710 ;
        RECT 1465.660 869.390 1465.920 869.710 ;
        RECT 1465.260 786.490 1465.400 869.390 ;
        RECT 1464.800 786.350 1465.400 786.490 ;
        RECT 1464.800 785.130 1464.940 786.350 ;
        RECT 1464.800 784.990 1465.400 785.130 ;
        RECT 1465.260 594.050 1465.400 784.990 ;
        RECT 1464.800 593.910 1465.400 594.050 ;
        RECT 1464.800 593.370 1464.940 593.910 ;
        RECT 1464.800 593.230 1465.400 593.370 ;
        RECT 1465.260 483.210 1465.400 593.230 ;
        RECT 1465.260 483.070 1465.860 483.210 ;
        RECT 1465.720 410.710 1465.860 483.070 ;
        RECT 1465.660 410.390 1465.920 410.710 ;
        RECT 1465.200 386.250 1465.460 386.570 ;
        RECT 1465.260 207.130 1465.400 386.250 ;
        RECT 1464.800 206.990 1465.400 207.130 ;
        RECT 1464.800 206.450 1464.940 206.990 ;
        RECT 1464.800 206.310 1465.400 206.450 ;
        RECT 1465.260 110.570 1465.400 206.310 ;
        RECT 1464.800 110.430 1465.400 110.570 ;
        RECT 1464.800 109.890 1464.940 110.430 ;
        RECT 1464.800 109.750 1465.400 109.890 ;
        RECT 1465.260 17.330 1465.400 109.750 ;
        RECT 1180.000 17.010 1180.260 17.330 ;
        RECT 1465.200 17.010 1465.460 17.330 ;
        RECT 1180.060 2.400 1180.200 17.010 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
      LAYER via2 ;
        RECT 1465.190 1200.400 1465.470 1200.680 ;
        RECT 1466.110 1200.400 1466.390 1200.680 ;
      LAYER met3 ;
        RECT 1465.165 1200.690 1465.495 1200.705 ;
        RECT 1466.085 1200.690 1466.415 1200.705 ;
        RECT 1465.165 1200.390 1466.415 1200.690 ;
        RECT 1465.165 1200.375 1465.495 1200.390 ;
        RECT 1466.085 1200.375 1466.415 1200.390 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1197.790 -4.800 1198.350 0.300 ;
=======
        RECT 1473.010 1700.410 1473.290 1704.000 ;
        RECT 1472.160 1700.270 1473.290 1700.410 ;
        RECT 1472.160 18.885 1472.300 1700.270 ;
        RECT 1473.010 1700.000 1473.290 1700.270 ;
        RECT 1197.930 18.515 1198.210 18.885 ;
        RECT 1472.090 18.515 1472.370 18.885 ;
        RECT 1198.000 2.400 1198.140 18.515 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
      LAYER via2 ;
        RECT 1197.930 18.560 1198.210 18.840 ;
        RECT 1472.090 18.560 1472.370 18.840 ;
      LAYER met3 ;
        RECT 1197.905 18.850 1198.235 18.865 ;
        RECT 1472.065 18.850 1472.395 18.865 ;
        RECT 1197.905 18.550 1472.395 18.850 ;
        RECT 1197.905 18.535 1198.235 18.550 ;
        RECT 1472.065 18.535 1472.395 18.550 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1476.670 39.000 1476.990 39.060 ;
        RECT 1478.050 39.000 1478.370 39.060 ;
        RECT 1476.670 38.860 1478.370 39.000 ;
        RECT 1476.670 38.800 1476.990 38.860 ;
        RECT 1478.050 38.800 1478.370 38.860 ;
      LAYER via ;
        RECT 1476.700 38.800 1476.960 39.060 ;
        RECT 1478.080 38.800 1478.340 39.060 ;
      LAYER met2 ;
        RECT 1478.070 1700.000 1478.350 1704.000 ;
        RECT 1478.140 39.090 1478.280 1700.000 ;
        RECT 1476.700 38.770 1476.960 39.090 ;
        RECT 1478.080 38.770 1478.340 39.090 ;
        RECT 1476.760 20.245 1476.900 38.770 ;
        RECT 1215.870 19.875 1216.150 20.245 ;
        RECT 1476.690 19.875 1476.970 20.245 ;
        RECT 1215.940 2.400 1216.080 19.875 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
      LAYER via2 ;
        RECT 1215.870 19.920 1216.150 20.200 ;
        RECT 1476.690 19.920 1476.970 20.200 ;
      LAYER met3 ;
        RECT 1215.845 20.210 1216.175 20.225 ;
        RECT 1476.665 20.210 1476.995 20.225 ;
        RECT 1215.845 19.910 1476.995 20.210 ;
        RECT 1215.845 19.895 1216.175 19.910 ;
        RECT 1476.665 19.895 1476.995 19.910 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 0.300 ;
=======
      LAYER li1 ;
        RECT 1438.105 1684.445 1438.275 1687.335 ;
      LAYER mcon ;
        RECT 1438.105 1687.165 1438.275 1687.335 ;
      LAYER met1 ;
        RECT 1259.550 1687.320 1259.870 1687.380 ;
        RECT 1438.045 1687.320 1438.335 1687.365 ;
        RECT 1259.550 1687.180 1438.335 1687.320 ;
        RECT 1259.550 1687.120 1259.870 1687.180 ;
        RECT 1438.045 1687.135 1438.335 1687.180 ;
        RECT 1438.045 1684.600 1438.335 1684.645 ;
        RECT 1438.045 1684.460 1472.760 1684.600 ;
        RECT 1438.045 1684.415 1438.335 1684.460 ;
        RECT 1472.620 1684.260 1472.760 1684.460 ;
        RECT 1482.650 1684.260 1482.970 1684.320 ;
        RECT 1472.620 1684.120 1482.970 1684.260 ;
        RECT 1482.650 1684.060 1482.970 1684.120 ;
        RECT 1233.790 20.300 1234.110 20.360 ;
        RECT 1259.550 20.300 1259.870 20.360 ;
        RECT 1233.790 20.160 1259.870 20.300 ;
        RECT 1233.790 20.100 1234.110 20.160 ;
        RECT 1259.550 20.100 1259.870 20.160 ;
      LAYER via ;
        RECT 1259.580 1687.120 1259.840 1687.380 ;
        RECT 1482.680 1684.060 1482.940 1684.320 ;
        RECT 1233.820 20.100 1234.080 20.360 ;
        RECT 1259.580 20.100 1259.840 20.360 ;
      LAYER met2 ;
        RECT 1482.670 1700.000 1482.950 1704.000 ;
        RECT 1259.580 1687.090 1259.840 1687.410 ;
        RECT 1259.640 20.390 1259.780 1687.090 ;
        RECT 1482.740 1684.350 1482.880 1700.000 ;
        RECT 1482.680 1684.030 1482.940 1684.350 ;
        RECT 1233.820 20.070 1234.080 20.390 ;
        RECT 1259.580 20.070 1259.840 20.390 ;
        RECT 1233.880 2.400 1234.020 20.070 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1259.090 1686.980 1259.410 1687.040 ;
        RECT 1486.330 1686.980 1486.650 1687.040 ;
        RECT 1259.090 1686.840 1486.650 1686.980 ;
        RECT 1259.090 1686.780 1259.410 1686.840 ;
        RECT 1486.330 1686.780 1486.650 1686.840 ;
        RECT 1251.730 20.640 1252.050 20.700 ;
        RECT 1259.090 20.640 1259.410 20.700 ;
        RECT 1251.730 20.500 1259.410 20.640 ;
        RECT 1251.730 20.440 1252.050 20.500 ;
        RECT 1259.090 20.440 1259.410 20.500 ;
      LAYER via ;
        RECT 1259.120 1686.780 1259.380 1687.040 ;
        RECT 1486.360 1686.780 1486.620 1687.040 ;
        RECT 1251.760 20.440 1252.020 20.700 ;
        RECT 1259.120 20.440 1259.380 20.700 ;
      LAYER met2 ;
        RECT 1487.730 1700.410 1488.010 1704.000 ;
        RECT 1486.420 1700.270 1488.010 1700.410 ;
        RECT 1486.420 1687.070 1486.560 1700.270 ;
        RECT 1487.730 1700.000 1488.010 1700.270 ;
        RECT 1259.120 1686.750 1259.380 1687.070 ;
        RECT 1486.360 1686.750 1486.620 1687.070 ;
        RECT 1259.180 20.730 1259.320 1686.750 ;
        RECT 1251.760 20.410 1252.020 20.730 ;
        RECT 1259.120 20.410 1259.380 20.730 ;
        RECT 1251.820 2.400 1251.960 20.410 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 0.300 ;
=======
      LAYER li1 ;
        RECT 1341.965 1642.965 1342.135 1689.035 ;
        RECT 1308.385 1580.065 1308.555 1594.175 ;
        RECT 1308.385 1145.885 1308.555 1193.655 ;
        RECT 1309.305 807.245 1309.475 821.355 ;
        RECT 1309.305 421.345 1309.475 469.115 ;
        RECT 1309.765 379.185 1309.935 420.835 ;
        RECT 1307.925 34.425 1308.095 82.875 ;
      LAYER mcon ;
        RECT 1341.965 1688.865 1342.135 1689.035 ;
        RECT 1308.385 1594.005 1308.555 1594.175 ;
        RECT 1308.385 1193.485 1308.555 1193.655 ;
        RECT 1309.305 821.185 1309.475 821.355 ;
        RECT 1309.305 468.945 1309.475 469.115 ;
        RECT 1309.765 420.665 1309.935 420.835 ;
        RECT 1307.925 82.705 1308.095 82.875 ;
      LAYER met1 ;
        RECT 1341.905 1689.020 1342.195 1689.065 ;
        RECT 1492.310 1689.020 1492.630 1689.080 ;
        RECT 1341.905 1688.880 1492.630 1689.020 ;
        RECT 1341.905 1688.835 1342.195 1688.880 ;
        RECT 1492.310 1688.820 1492.630 1688.880 ;
        RECT 1308.770 1643.120 1309.090 1643.180 ;
        RECT 1341.905 1643.120 1342.195 1643.165 ;
        RECT 1308.770 1642.980 1342.195 1643.120 ;
        RECT 1308.770 1642.920 1309.090 1642.980 ;
        RECT 1341.905 1642.935 1342.195 1642.980 ;
        RECT 1308.325 1594.160 1308.615 1594.205 ;
        RECT 1308.770 1594.160 1309.090 1594.220 ;
        RECT 1308.325 1594.020 1309.090 1594.160 ;
        RECT 1308.325 1593.975 1308.615 1594.020 ;
        RECT 1308.770 1593.960 1309.090 1594.020 ;
        RECT 1308.310 1580.220 1308.630 1580.280 ;
        RECT 1308.115 1580.080 1308.630 1580.220 ;
        RECT 1308.310 1580.020 1308.630 1580.080 ;
        RECT 1307.850 1490.460 1308.170 1490.520 ;
        RECT 1308.770 1490.460 1309.090 1490.520 ;
        RECT 1307.850 1490.320 1309.090 1490.460 ;
        RECT 1307.850 1490.260 1308.170 1490.320 ;
        RECT 1308.770 1490.260 1309.090 1490.320 ;
        RECT 1308.310 1249.060 1308.630 1249.120 ;
        RECT 1308.770 1249.060 1309.090 1249.120 ;
        RECT 1308.310 1248.920 1309.090 1249.060 ;
        RECT 1308.310 1248.860 1308.630 1248.920 ;
        RECT 1308.770 1248.860 1309.090 1248.920 ;
        RECT 1308.325 1193.640 1308.615 1193.685 ;
        RECT 1308.770 1193.640 1309.090 1193.700 ;
        RECT 1308.325 1193.500 1309.090 1193.640 ;
        RECT 1308.325 1193.455 1308.615 1193.500 ;
        RECT 1308.770 1193.440 1309.090 1193.500 ;
        RECT 1308.310 1146.040 1308.630 1146.100 ;
        RECT 1308.115 1145.900 1308.630 1146.040 ;
        RECT 1308.310 1145.840 1308.630 1145.900 ;
        RECT 1307.850 1145.360 1308.170 1145.420 ;
        RECT 1308.310 1145.360 1308.630 1145.420 ;
        RECT 1307.850 1145.220 1308.630 1145.360 ;
        RECT 1307.850 1145.160 1308.170 1145.220 ;
        RECT 1308.310 1145.160 1308.630 1145.220 ;
        RECT 1308.310 1072.940 1308.630 1073.000 ;
        RECT 1309.230 1072.940 1309.550 1073.000 ;
        RECT 1308.310 1072.800 1309.550 1072.940 ;
        RECT 1308.310 1072.740 1308.630 1072.800 ;
        RECT 1309.230 1072.740 1309.550 1072.800 ;
        RECT 1308.310 917.900 1308.630 917.960 ;
        RECT 1308.770 917.900 1309.090 917.960 ;
        RECT 1308.310 917.760 1309.090 917.900 ;
        RECT 1308.310 917.700 1308.630 917.760 ;
        RECT 1308.770 917.700 1309.090 917.760 ;
        RECT 1308.770 910.760 1309.090 910.820 ;
        RECT 1309.230 910.760 1309.550 910.820 ;
        RECT 1308.770 910.620 1309.550 910.760 ;
        RECT 1308.770 910.560 1309.090 910.620 ;
        RECT 1309.230 910.560 1309.550 910.620 ;
        RECT 1309.230 821.340 1309.550 821.400 ;
        RECT 1309.035 821.200 1309.550 821.340 ;
        RECT 1309.230 821.140 1309.550 821.200 ;
        RECT 1309.230 807.400 1309.550 807.460 ;
        RECT 1309.035 807.260 1309.550 807.400 ;
        RECT 1309.230 807.200 1309.550 807.260 ;
        RECT 1308.770 613.940 1309.090 614.000 ;
        RECT 1309.230 613.940 1309.550 614.000 ;
        RECT 1308.770 613.800 1309.550 613.940 ;
        RECT 1308.770 613.740 1309.090 613.800 ;
        RECT 1309.230 613.740 1309.550 613.800 ;
        RECT 1308.770 524.520 1309.090 524.580 ;
        RECT 1309.230 524.520 1309.550 524.580 ;
        RECT 1308.770 524.380 1309.550 524.520 ;
        RECT 1308.770 524.320 1309.090 524.380 ;
        RECT 1309.230 524.320 1309.550 524.380 ;
        RECT 1308.770 517.380 1309.090 517.440 ;
        RECT 1309.230 517.380 1309.550 517.440 ;
        RECT 1308.770 517.240 1309.550 517.380 ;
        RECT 1308.770 517.180 1309.090 517.240 ;
        RECT 1309.230 517.180 1309.550 517.240 ;
        RECT 1309.230 469.100 1309.550 469.160 ;
        RECT 1309.035 468.960 1309.550 469.100 ;
        RECT 1309.230 468.900 1309.550 468.960 ;
        RECT 1309.245 421.500 1309.535 421.545 ;
        RECT 1309.690 421.500 1310.010 421.560 ;
        RECT 1309.245 421.360 1310.010 421.500 ;
        RECT 1309.245 421.315 1309.535 421.360 ;
        RECT 1309.690 421.300 1310.010 421.360 ;
        RECT 1309.690 420.820 1310.010 420.880 ;
        RECT 1309.495 420.680 1310.010 420.820 ;
        RECT 1309.690 420.620 1310.010 420.680 ;
        RECT 1309.690 379.340 1310.010 379.400 ;
        RECT 1309.495 379.200 1310.010 379.340 ;
        RECT 1309.690 379.140 1310.010 379.200 ;
        RECT 1308.770 324.600 1309.090 324.660 ;
        RECT 1309.690 324.600 1310.010 324.660 ;
        RECT 1308.770 324.460 1310.010 324.600 ;
        RECT 1308.770 324.400 1309.090 324.460 ;
        RECT 1309.690 324.400 1310.010 324.460 ;
        RECT 1308.310 282.780 1308.630 282.840 ;
        RECT 1308.770 282.780 1309.090 282.840 ;
        RECT 1308.310 282.640 1309.090 282.780 ;
        RECT 1308.310 282.580 1308.630 282.640 ;
        RECT 1308.770 282.580 1309.090 282.640 ;
        RECT 1308.310 179.420 1308.630 179.480 ;
        RECT 1309.230 179.420 1309.550 179.480 ;
        RECT 1308.310 179.280 1309.550 179.420 ;
        RECT 1308.310 179.220 1308.630 179.280 ;
        RECT 1309.230 179.220 1309.550 179.280 ;
        RECT 1307.865 82.860 1308.155 82.905 ;
        RECT 1308.310 82.860 1308.630 82.920 ;
        RECT 1307.865 82.720 1308.630 82.860 ;
        RECT 1307.865 82.675 1308.155 82.720 ;
        RECT 1308.310 82.660 1308.630 82.720 ;
        RECT 1307.850 34.580 1308.170 34.640 ;
        RECT 1307.655 34.440 1308.170 34.580 ;
        RECT 1307.850 34.380 1308.170 34.440 ;
        RECT 1269.210 19.620 1269.530 19.680 ;
        RECT 1307.850 19.620 1308.170 19.680 ;
        RECT 1269.210 19.480 1308.170 19.620 ;
        RECT 1269.210 19.420 1269.530 19.480 ;
        RECT 1307.850 19.420 1308.170 19.480 ;
      LAYER via ;
        RECT 1492.340 1688.820 1492.600 1689.080 ;
        RECT 1308.800 1642.920 1309.060 1643.180 ;
        RECT 1308.800 1593.960 1309.060 1594.220 ;
        RECT 1308.340 1580.020 1308.600 1580.280 ;
        RECT 1307.880 1490.260 1308.140 1490.520 ;
        RECT 1308.800 1490.260 1309.060 1490.520 ;
        RECT 1308.340 1248.860 1308.600 1249.120 ;
        RECT 1308.800 1248.860 1309.060 1249.120 ;
        RECT 1308.800 1193.440 1309.060 1193.700 ;
        RECT 1308.340 1145.840 1308.600 1146.100 ;
        RECT 1307.880 1145.160 1308.140 1145.420 ;
        RECT 1308.340 1145.160 1308.600 1145.420 ;
        RECT 1308.340 1072.740 1308.600 1073.000 ;
        RECT 1309.260 1072.740 1309.520 1073.000 ;
        RECT 1308.340 917.700 1308.600 917.960 ;
        RECT 1308.800 917.700 1309.060 917.960 ;
        RECT 1308.800 910.560 1309.060 910.820 ;
        RECT 1309.260 910.560 1309.520 910.820 ;
        RECT 1309.260 821.140 1309.520 821.400 ;
        RECT 1309.260 807.200 1309.520 807.460 ;
        RECT 1308.800 613.740 1309.060 614.000 ;
        RECT 1309.260 613.740 1309.520 614.000 ;
        RECT 1308.800 524.320 1309.060 524.580 ;
        RECT 1309.260 524.320 1309.520 524.580 ;
        RECT 1308.800 517.180 1309.060 517.440 ;
        RECT 1309.260 517.180 1309.520 517.440 ;
        RECT 1309.260 468.900 1309.520 469.160 ;
        RECT 1309.720 421.300 1309.980 421.560 ;
        RECT 1309.720 420.620 1309.980 420.880 ;
        RECT 1309.720 379.140 1309.980 379.400 ;
        RECT 1308.800 324.400 1309.060 324.660 ;
        RECT 1309.720 324.400 1309.980 324.660 ;
        RECT 1308.340 282.580 1308.600 282.840 ;
        RECT 1308.800 282.580 1309.060 282.840 ;
        RECT 1308.340 179.220 1308.600 179.480 ;
        RECT 1309.260 179.220 1309.520 179.480 ;
        RECT 1308.340 82.660 1308.600 82.920 ;
        RECT 1307.880 34.380 1308.140 34.640 ;
        RECT 1269.240 19.420 1269.500 19.680 ;
        RECT 1307.880 19.420 1308.140 19.680 ;
      LAYER met2 ;
        RECT 1492.330 1700.000 1492.610 1704.000 ;
        RECT 1492.400 1689.110 1492.540 1700.000 ;
        RECT 1492.340 1688.790 1492.600 1689.110 ;
        RECT 1308.800 1642.890 1309.060 1643.210 ;
        RECT 1308.860 1594.250 1309.000 1642.890 ;
        RECT 1308.800 1593.930 1309.060 1594.250 ;
        RECT 1308.340 1579.990 1308.600 1580.310 ;
        RECT 1308.400 1514.770 1308.540 1579.990 ;
        RECT 1308.400 1514.630 1309.460 1514.770 ;
        RECT 1309.320 1510.690 1309.460 1514.630 ;
        RECT 1308.860 1510.550 1309.460 1510.690 ;
        RECT 1308.860 1490.550 1309.000 1510.550 ;
        RECT 1307.880 1490.230 1308.140 1490.550 ;
        RECT 1308.800 1490.230 1309.060 1490.550 ;
        RECT 1307.940 1435.325 1308.080 1490.230 ;
        RECT 1307.870 1434.955 1308.150 1435.325 ;
        RECT 1309.250 1434.955 1309.530 1435.325 ;
        RECT 1309.320 1387.725 1309.460 1434.955 ;
        RECT 1309.250 1387.355 1309.530 1387.725 ;
        RECT 1309.250 1386.675 1309.530 1387.045 ;
        RECT 1309.320 1363.130 1309.460 1386.675 ;
        RECT 1308.860 1362.990 1309.460 1363.130 ;
        RECT 1308.860 1249.150 1309.000 1362.990 ;
        RECT 1308.340 1249.005 1308.600 1249.150 ;
        RECT 1308.330 1248.635 1308.610 1249.005 ;
        RECT 1308.800 1248.830 1309.060 1249.150 ;
        RECT 1309.250 1248.635 1309.530 1249.005 ;
        RECT 1309.320 1221.010 1309.460 1248.635 ;
        RECT 1308.860 1220.870 1309.460 1221.010 ;
        RECT 1308.860 1193.730 1309.000 1220.870 ;
        RECT 1308.800 1193.410 1309.060 1193.730 ;
        RECT 1308.340 1145.810 1308.600 1146.130 ;
        RECT 1308.400 1145.450 1308.540 1145.810 ;
        RECT 1307.880 1145.130 1308.140 1145.450 ;
        RECT 1308.340 1145.130 1308.600 1145.450 ;
        RECT 1307.940 1097.365 1308.080 1145.130 ;
        RECT 1307.870 1096.995 1308.150 1097.365 ;
        RECT 1309.250 1096.995 1309.530 1097.365 ;
        RECT 1309.320 1073.030 1309.460 1096.995 ;
        RECT 1308.340 1072.710 1308.600 1073.030 ;
        RECT 1309.260 1072.710 1309.520 1073.030 ;
        RECT 1308.400 917.990 1308.540 1072.710 ;
        RECT 1308.340 917.670 1308.600 917.990 ;
        RECT 1308.800 917.670 1309.060 917.990 ;
        RECT 1308.860 910.850 1309.000 917.670 ;
        RECT 1308.800 910.530 1309.060 910.850 ;
        RECT 1309.260 910.530 1309.520 910.850 ;
        RECT 1309.320 821.430 1309.460 910.530 ;
        RECT 1309.260 821.110 1309.520 821.430 ;
        RECT 1309.260 807.170 1309.520 807.490 ;
        RECT 1309.320 782.410 1309.460 807.170 ;
        RECT 1308.400 782.270 1309.460 782.410 ;
        RECT 1308.400 741.610 1308.540 782.270 ;
        RECT 1308.400 741.470 1309.000 741.610 ;
        RECT 1308.860 669.530 1309.000 741.470 ;
        RECT 1308.400 669.390 1309.000 669.530 ;
        RECT 1308.400 644.370 1308.540 669.390 ;
        RECT 1308.400 644.230 1309.000 644.370 ;
        RECT 1308.860 614.030 1309.000 644.230 ;
        RECT 1308.800 613.710 1309.060 614.030 ;
        RECT 1309.260 613.710 1309.520 614.030 ;
        RECT 1309.320 524.610 1309.460 613.710 ;
        RECT 1308.800 524.290 1309.060 524.610 ;
        RECT 1309.260 524.290 1309.520 524.610 ;
        RECT 1308.860 517.470 1309.000 524.290 ;
        RECT 1308.800 517.150 1309.060 517.470 ;
        RECT 1309.260 517.150 1309.520 517.470 ;
        RECT 1309.320 469.190 1309.460 517.150 ;
        RECT 1309.260 468.870 1309.520 469.190 ;
        RECT 1309.720 421.270 1309.980 421.590 ;
        RECT 1309.780 420.910 1309.920 421.270 ;
        RECT 1309.720 420.590 1309.980 420.910 ;
        RECT 1309.720 379.110 1309.980 379.430 ;
        RECT 1309.780 324.690 1309.920 379.110 ;
        RECT 1308.800 324.370 1309.060 324.690 ;
        RECT 1309.720 324.370 1309.980 324.690 ;
        RECT 1308.860 282.870 1309.000 324.370 ;
        RECT 1308.340 282.550 1308.600 282.870 ;
        RECT 1308.800 282.550 1309.060 282.870 ;
        RECT 1308.400 258.130 1308.540 282.550 ;
        RECT 1308.400 257.990 1309.000 258.130 ;
        RECT 1308.860 186.730 1309.000 257.990 ;
        RECT 1308.400 186.590 1309.000 186.730 ;
        RECT 1308.400 179.510 1308.540 186.590 ;
        RECT 1308.340 179.190 1308.600 179.510 ;
        RECT 1309.260 179.190 1309.520 179.510 ;
        RECT 1309.320 107.170 1309.460 179.190 ;
        RECT 1308.400 107.030 1309.460 107.170 ;
        RECT 1308.400 82.950 1308.540 107.030 ;
        RECT 1308.340 82.630 1308.600 82.950 ;
        RECT 1307.880 34.350 1308.140 34.670 ;
        RECT 1307.940 19.710 1308.080 34.350 ;
        RECT 1269.240 19.390 1269.500 19.710 ;
        RECT 1307.880 19.390 1308.140 19.710 ;
        RECT 1269.300 2.400 1269.440 19.390 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
      LAYER via2 ;
        RECT 1307.870 1435.000 1308.150 1435.280 ;
        RECT 1309.250 1435.000 1309.530 1435.280 ;
        RECT 1309.250 1387.400 1309.530 1387.680 ;
        RECT 1309.250 1386.720 1309.530 1387.000 ;
        RECT 1308.330 1248.680 1308.610 1248.960 ;
        RECT 1309.250 1248.680 1309.530 1248.960 ;
        RECT 1307.870 1097.040 1308.150 1097.320 ;
        RECT 1309.250 1097.040 1309.530 1097.320 ;
      LAYER met3 ;
        RECT 1307.845 1435.290 1308.175 1435.305 ;
        RECT 1309.225 1435.290 1309.555 1435.305 ;
        RECT 1307.845 1434.990 1309.555 1435.290 ;
        RECT 1307.845 1434.975 1308.175 1434.990 ;
        RECT 1309.225 1434.975 1309.555 1434.990 ;
        RECT 1309.225 1387.690 1309.555 1387.705 ;
        RECT 1308.550 1387.390 1309.555 1387.690 ;
        RECT 1308.550 1387.010 1308.850 1387.390 ;
        RECT 1309.225 1387.375 1309.555 1387.390 ;
        RECT 1309.225 1387.010 1309.555 1387.025 ;
        RECT 1308.550 1386.710 1309.555 1387.010 ;
        RECT 1309.225 1386.695 1309.555 1386.710 ;
        RECT 1308.305 1248.970 1308.635 1248.985 ;
        RECT 1309.225 1248.970 1309.555 1248.985 ;
        RECT 1308.305 1248.670 1309.555 1248.970 ;
        RECT 1308.305 1248.655 1308.635 1248.670 ;
        RECT 1309.225 1248.655 1309.555 1248.670 ;
        RECT 1307.845 1097.330 1308.175 1097.345 ;
        RECT 1309.225 1097.330 1309.555 1097.345 ;
        RECT 1307.845 1097.030 1309.555 1097.330 ;
        RECT 1307.845 1097.015 1308.175 1097.030 ;
        RECT 1309.225 1097.015 1309.555 1097.030 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1290.370 1687.660 1290.690 1687.720 ;
        RECT 1497.370 1687.660 1497.690 1687.720 ;
        RECT 1290.370 1687.520 1497.690 1687.660 ;
        RECT 1290.370 1687.460 1290.690 1687.520 ;
        RECT 1497.370 1687.460 1497.690 1687.520 ;
        RECT 1289.910 671.200 1290.230 671.460 ;
        RECT 1290.000 670.780 1290.140 671.200 ;
        RECT 1289.910 670.520 1290.230 670.780 ;
        RECT 1289.910 616.120 1290.230 616.380 ;
        RECT 1290.000 615.700 1290.140 616.120 ;
        RECT 1289.910 615.440 1290.230 615.700 ;
        RECT 1287.150 20.640 1287.470 20.700 ;
        RECT 1289.910 20.640 1290.230 20.700 ;
        RECT 1287.150 20.500 1290.230 20.640 ;
        RECT 1287.150 20.440 1287.470 20.500 ;
        RECT 1289.910 20.440 1290.230 20.500 ;
      LAYER via ;
        RECT 1290.400 1687.460 1290.660 1687.720 ;
        RECT 1497.400 1687.460 1497.660 1687.720 ;
        RECT 1289.940 671.200 1290.200 671.460 ;
        RECT 1289.940 670.520 1290.200 670.780 ;
        RECT 1289.940 616.120 1290.200 616.380 ;
        RECT 1289.940 615.440 1290.200 615.700 ;
        RECT 1287.180 20.440 1287.440 20.700 ;
        RECT 1289.940 20.440 1290.200 20.700 ;
      LAYER met2 ;
        RECT 1497.390 1700.000 1497.670 1704.000 ;
        RECT 1497.460 1687.750 1497.600 1700.000 ;
        RECT 1290.400 1687.430 1290.660 1687.750 ;
        RECT 1497.400 1687.430 1497.660 1687.750 ;
        RECT 1290.460 1685.450 1290.600 1687.430 ;
        RECT 1290.000 1685.310 1290.600 1685.450 ;
        RECT 1290.000 671.490 1290.140 1685.310 ;
        RECT 1289.940 671.170 1290.200 671.490 ;
        RECT 1289.940 670.490 1290.200 670.810 ;
        RECT 1290.000 616.410 1290.140 670.490 ;
        RECT 1289.940 616.090 1290.200 616.410 ;
        RECT 1289.940 615.410 1290.200 615.730 ;
        RECT 1290.000 20.730 1290.140 615.410 ;
        RECT 1287.180 20.410 1287.440 20.730 ;
        RECT 1289.940 20.410 1290.200 20.730 ;
        RECT 1287.240 2.400 1287.380 20.410 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1310.610 1689.020 1310.930 1689.080 ;
        RECT 1310.610 1688.880 1341.660 1689.020 ;
        RECT 1310.610 1688.820 1310.930 1688.880 ;
        RECT 1341.520 1688.680 1341.660 1688.880 ;
        RECT 1501.970 1688.680 1502.290 1688.740 ;
        RECT 1341.520 1688.540 1502.290 1688.680 ;
        RECT 1501.970 1688.480 1502.290 1688.540 ;
        RECT 1305.090 20.300 1305.410 20.360 ;
        RECT 1310.610 20.300 1310.930 20.360 ;
        RECT 1305.090 20.160 1310.930 20.300 ;
        RECT 1305.090 20.100 1305.410 20.160 ;
        RECT 1310.610 20.100 1310.930 20.160 ;
      LAYER via ;
        RECT 1310.640 1688.820 1310.900 1689.080 ;
        RECT 1502.000 1688.480 1502.260 1688.740 ;
        RECT 1305.120 20.100 1305.380 20.360 ;
        RECT 1310.640 20.100 1310.900 20.360 ;
      LAYER met2 ;
        RECT 1501.990 1700.000 1502.270 1704.000 ;
        RECT 1310.640 1688.790 1310.900 1689.110 ;
        RECT 1310.700 20.390 1310.840 1688.790 ;
        RECT 1502.060 1688.770 1502.200 1700.000 ;
        RECT 1502.000 1688.450 1502.260 1688.770 ;
        RECT 1305.120 20.070 1305.380 20.390 ;
        RECT 1310.640 20.070 1310.900 20.390 ;
        RECT 1305.180 2.400 1305.320 20.070 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 0.300 ;
=======
      LAYER li1 ;
        RECT 1390.265 1686.485 1390.435 1690.055 ;
      LAYER mcon ;
        RECT 1390.265 1689.885 1390.435 1690.055 ;
      LAYER met1 ;
        RECT 1390.205 1690.040 1390.495 1690.085 ;
        RECT 1507.030 1690.040 1507.350 1690.100 ;
        RECT 1390.205 1689.900 1507.350 1690.040 ;
        RECT 1390.205 1689.855 1390.495 1689.900 ;
        RECT 1507.030 1689.840 1507.350 1689.900 ;
        RECT 1348.790 1686.640 1349.110 1686.700 ;
        RECT 1390.205 1686.640 1390.495 1686.685 ;
        RECT 1348.790 1686.500 1390.495 1686.640 ;
        RECT 1348.790 1686.440 1349.110 1686.500 ;
        RECT 1390.205 1686.455 1390.495 1686.500 ;
        RECT 1323.030 15.200 1323.350 15.260 ;
        RECT 1348.790 15.200 1349.110 15.260 ;
        RECT 1323.030 15.060 1349.110 15.200 ;
        RECT 1323.030 15.000 1323.350 15.060 ;
        RECT 1348.790 15.000 1349.110 15.060 ;
      LAYER via ;
        RECT 1507.060 1689.840 1507.320 1690.100 ;
        RECT 1348.820 1686.440 1349.080 1686.700 ;
        RECT 1323.060 15.000 1323.320 15.260 ;
        RECT 1348.820 15.000 1349.080 15.260 ;
      LAYER met2 ;
        RECT 1507.050 1700.000 1507.330 1704.000 ;
        RECT 1507.120 1690.130 1507.260 1700.000 ;
        RECT 1507.060 1689.810 1507.320 1690.130 ;
        RECT 1348.820 1686.410 1349.080 1686.730 ;
        RECT 1348.880 15.290 1349.020 1686.410 ;
        RECT 1323.060 14.970 1323.320 15.290 ;
        RECT 1348.820 14.970 1349.080 15.290 ;
        RECT 1323.120 2.400 1323.260 14.970 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 0.300 ;
=======
      LAYER li1 ;
        RECT 1389.805 1686.145 1389.975 1689.715 ;
      LAYER mcon ;
        RECT 1389.805 1689.545 1389.975 1689.715 ;
      LAYER met1 ;
        RECT 1511.630 1690.380 1511.950 1690.440 ;
        RECT 1507.580 1690.240 1511.950 1690.380 ;
        RECT 1389.745 1689.700 1390.035 1689.745 ;
        RECT 1507.580 1689.700 1507.720 1690.240 ;
        RECT 1511.630 1690.180 1511.950 1690.240 ;
        RECT 1389.745 1689.560 1507.720 1689.700 ;
        RECT 1389.745 1689.515 1390.035 1689.560 ;
        RECT 1345.110 1686.300 1345.430 1686.360 ;
        RECT 1389.745 1686.300 1390.035 1686.345 ;
        RECT 1345.110 1686.160 1390.035 1686.300 ;
        RECT 1345.110 1686.100 1345.430 1686.160 ;
        RECT 1389.745 1686.115 1390.035 1686.160 ;
        RECT 1340.510 20.640 1340.830 20.700 ;
        RECT 1345.110 20.640 1345.430 20.700 ;
        RECT 1340.510 20.500 1345.430 20.640 ;
        RECT 1340.510 20.440 1340.830 20.500 ;
        RECT 1345.110 20.440 1345.430 20.500 ;
      LAYER via ;
        RECT 1511.660 1690.180 1511.920 1690.440 ;
        RECT 1345.140 1686.100 1345.400 1686.360 ;
        RECT 1340.540 20.440 1340.800 20.700 ;
        RECT 1345.140 20.440 1345.400 20.700 ;
      LAYER met2 ;
        RECT 1511.650 1700.000 1511.930 1704.000 ;
        RECT 1511.720 1690.470 1511.860 1700.000 ;
        RECT 1511.660 1690.150 1511.920 1690.470 ;
        RECT 1345.140 1686.070 1345.400 1686.390 ;
        RECT 1345.200 20.730 1345.340 1686.070 ;
        RECT 1340.540 20.410 1340.800 20.730 ;
        RECT 1345.140 20.410 1345.400 20.730 ;
        RECT 1340.600 2.400 1340.740 20.410 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 0.300 ;
=======
      LAYER met1 ;
        RECT 1333.150 1678.140 1333.470 1678.200 ;
        RECT 1337.290 1678.140 1337.610 1678.200 ;
        RECT 1333.150 1678.000 1337.610 1678.140 ;
        RECT 1333.150 1677.940 1333.470 1678.000 ;
        RECT 1337.290 1677.940 1337.610 1678.000 ;
        RECT 698.350 46.820 698.670 46.880 ;
        RECT 1333.150 46.820 1333.470 46.880 ;
        RECT 698.350 46.680 1333.470 46.820 ;
        RECT 698.350 46.620 698.670 46.680 ;
        RECT 1333.150 46.620 1333.470 46.680 ;
      LAYER via ;
        RECT 1333.180 1677.940 1333.440 1678.200 ;
        RECT 1337.320 1677.940 1337.580 1678.200 ;
        RECT 698.380 46.620 698.640 46.880 ;
        RECT 1333.180 46.620 1333.440 46.880 ;
      LAYER met2 ;
        RECT 1338.230 1700.410 1338.510 1704.000 ;
        RECT 1337.380 1700.270 1338.510 1700.410 ;
        RECT 1337.380 1678.230 1337.520 1700.270 ;
        RECT 1338.230 1700.000 1338.510 1700.270 ;
        RECT 1333.180 1677.910 1333.440 1678.230 ;
        RECT 1337.320 1677.910 1337.580 1678.230 ;
        RECT 1333.240 46.910 1333.380 1677.910 ;
        RECT 698.380 46.590 698.640 46.910 ;
        RECT 1333.180 46.590 1333.440 46.910 ;
        RECT 698.440 2.400 698.580 46.590 ;
        RECT 698.230 -4.800 698.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 0.300 ;
=======
      LAYER li1 ;
        RECT 1513.085 1594.005 1513.255 1642.115 ;
        RECT 1514.005 1497.445 1514.175 1511.215 ;
        RECT 1513.085 766.105 1513.255 790.075 ;
        RECT 1513.085 544.765 1513.255 596.955 ;
        RECT 1513.545 447.865 1513.715 524.195 ;
        RECT 1513.545 157.845 1513.715 234.515 ;
        RECT 1514.005 89.845 1514.175 137.955 ;
      LAYER mcon ;
        RECT 1513.085 1641.945 1513.255 1642.115 ;
        RECT 1514.005 1511.045 1514.175 1511.215 ;
        RECT 1513.085 789.905 1513.255 790.075 ;
        RECT 1513.085 596.785 1513.255 596.955 ;
        RECT 1513.545 524.025 1513.715 524.195 ;
        RECT 1513.545 234.345 1513.715 234.515 ;
        RECT 1514.005 137.785 1514.175 137.955 ;
      LAYER met1 ;
        RECT 1513.010 1666.580 1513.330 1666.640 ;
        RECT 1515.310 1666.580 1515.630 1666.640 ;
        RECT 1513.010 1666.440 1515.630 1666.580 ;
        RECT 1513.010 1666.380 1513.330 1666.440 ;
        RECT 1515.310 1666.380 1515.630 1666.440 ;
        RECT 1513.010 1642.100 1513.330 1642.160 ;
        RECT 1512.815 1641.960 1513.330 1642.100 ;
        RECT 1513.010 1641.900 1513.330 1641.960 ;
        RECT 1513.025 1594.160 1513.315 1594.205 ;
        RECT 1513.930 1594.160 1514.250 1594.220 ;
        RECT 1513.025 1594.020 1514.250 1594.160 ;
        RECT 1513.025 1593.975 1513.315 1594.020 ;
        RECT 1513.930 1593.960 1514.250 1594.020 ;
        RECT 1513.930 1569.680 1514.250 1569.740 ;
        RECT 1514.850 1569.680 1515.170 1569.740 ;
        RECT 1513.930 1569.540 1515.170 1569.680 ;
        RECT 1513.930 1569.480 1514.250 1569.540 ;
        RECT 1514.850 1569.480 1515.170 1569.540 ;
        RECT 1513.930 1511.200 1514.250 1511.260 ;
        RECT 1513.735 1511.060 1514.250 1511.200 ;
        RECT 1513.930 1511.000 1514.250 1511.060 ;
        RECT 1513.930 1497.600 1514.250 1497.660 ;
        RECT 1513.735 1497.460 1514.250 1497.600 ;
        RECT 1513.930 1497.400 1514.250 1497.460 ;
        RECT 1513.010 1435.380 1513.330 1435.440 ;
        RECT 1513.930 1435.380 1514.250 1435.440 ;
        RECT 1513.010 1435.240 1514.250 1435.380 ;
        RECT 1513.010 1435.180 1513.330 1435.240 ;
        RECT 1513.930 1435.180 1514.250 1435.240 ;
        RECT 1513.010 1393.900 1513.330 1393.960 ;
        RECT 1513.930 1393.900 1514.250 1393.960 ;
        RECT 1513.010 1393.760 1514.250 1393.900 ;
        RECT 1513.010 1393.700 1513.330 1393.760 ;
        RECT 1513.930 1393.700 1514.250 1393.760 ;
        RECT 1513.470 1338.820 1513.790 1338.880 ;
        RECT 1513.930 1338.820 1514.250 1338.880 ;
        RECT 1513.470 1338.680 1514.250 1338.820 ;
        RECT 1513.470 1338.620 1513.790 1338.680 ;
        RECT 1513.930 1338.620 1514.250 1338.680 ;
        RECT 1513.010 1159.300 1513.330 1159.360 ;
        RECT 1513.470 1159.300 1513.790 1159.360 ;
        RECT 1513.010 1159.160 1513.790 1159.300 ;
        RECT 1513.010 1159.100 1513.330 1159.160 ;
        RECT 1513.470 1159.100 1513.790 1159.160 ;
        RECT 1513.930 1111.020 1514.250 1111.080 ;
        RECT 1513.560 1110.880 1514.250 1111.020 ;
        RECT 1513.560 1110.740 1513.700 1110.880 ;
        RECT 1513.930 1110.820 1514.250 1110.880 ;
        RECT 1513.470 1110.480 1513.790 1110.740 ;
        RECT 1513.930 1096.740 1514.250 1096.800 ;
        RECT 1514.850 1096.740 1515.170 1096.800 ;
        RECT 1513.930 1096.600 1515.170 1096.740 ;
        RECT 1513.930 1096.540 1514.250 1096.600 ;
        RECT 1514.850 1096.540 1515.170 1096.600 ;
        RECT 1513.470 1028.540 1513.790 1028.800 ;
        RECT 1513.560 1028.120 1513.700 1028.540 ;
        RECT 1513.470 1027.860 1513.790 1028.120 ;
        RECT 1513.010 966.180 1513.330 966.240 ;
        RECT 1513.470 966.180 1513.790 966.240 ;
        RECT 1513.010 966.040 1513.790 966.180 ;
        RECT 1513.010 965.980 1513.330 966.040 ;
        RECT 1513.470 965.980 1513.790 966.040 ;
        RECT 1513.930 917.900 1514.250 917.960 ;
        RECT 1515.310 917.900 1515.630 917.960 ;
        RECT 1513.930 917.760 1515.630 917.900 ;
        RECT 1513.930 917.700 1514.250 917.760 ;
        RECT 1515.310 917.700 1515.630 917.760 ;
        RECT 1513.930 883.560 1514.250 883.620 ;
        RECT 1515.310 883.560 1515.630 883.620 ;
        RECT 1513.930 883.420 1515.630 883.560 ;
        RECT 1513.930 883.360 1514.250 883.420 ;
        RECT 1515.310 883.360 1515.630 883.420 ;
        RECT 1513.010 838.340 1513.330 838.400 ;
        RECT 1513.930 838.340 1514.250 838.400 ;
        RECT 1513.010 838.200 1514.250 838.340 ;
        RECT 1513.010 838.140 1513.330 838.200 ;
        RECT 1513.930 838.140 1514.250 838.200 ;
        RECT 1513.010 790.060 1513.330 790.120 ;
        RECT 1512.815 789.920 1513.330 790.060 ;
        RECT 1513.010 789.860 1513.330 789.920 ;
        RECT 1513.025 766.260 1513.315 766.305 ;
        RECT 1513.930 766.260 1514.250 766.320 ;
        RECT 1513.025 766.120 1514.250 766.260 ;
        RECT 1513.025 766.075 1513.315 766.120 ;
        RECT 1513.930 766.060 1514.250 766.120 ;
        RECT 1513.010 717.640 1513.330 717.700 ;
        RECT 1513.470 717.640 1513.790 717.700 ;
        RECT 1513.010 717.500 1513.790 717.640 ;
        RECT 1513.010 717.440 1513.330 717.500 ;
        RECT 1513.470 717.440 1513.790 717.500 ;
        RECT 1513.010 710.500 1513.330 710.560 ;
        RECT 1513.930 710.500 1514.250 710.560 ;
        RECT 1513.010 710.360 1514.250 710.500 ;
        RECT 1513.010 710.300 1513.330 710.360 ;
        RECT 1513.930 710.300 1514.250 710.360 ;
        RECT 1513.025 596.940 1513.315 596.985 ;
        RECT 1513.930 596.940 1514.250 597.000 ;
        RECT 1513.025 596.800 1514.250 596.940 ;
        RECT 1513.025 596.755 1513.315 596.800 ;
        RECT 1513.930 596.740 1514.250 596.800 ;
        RECT 1513.025 544.920 1513.315 544.965 ;
        RECT 1513.470 544.920 1513.790 544.980 ;
        RECT 1513.025 544.780 1513.790 544.920 ;
        RECT 1513.025 544.735 1513.315 544.780 ;
        RECT 1513.470 544.720 1513.790 544.780 ;
        RECT 1513.470 524.180 1513.790 524.240 ;
        RECT 1513.275 524.040 1513.790 524.180 ;
        RECT 1513.470 523.980 1513.790 524.040 ;
        RECT 1513.485 448.020 1513.775 448.065 ;
        RECT 1513.930 448.020 1514.250 448.080 ;
        RECT 1513.485 447.880 1514.250 448.020 ;
        RECT 1513.485 447.835 1513.775 447.880 ;
        RECT 1513.930 447.820 1514.250 447.880 ;
        RECT 1513.930 331.060 1514.250 331.120 ;
        RECT 1514.850 331.060 1515.170 331.120 ;
        RECT 1513.930 330.920 1515.170 331.060 ;
        RECT 1513.930 330.860 1514.250 330.920 ;
        RECT 1514.850 330.860 1515.170 330.920 ;
        RECT 1513.485 234.500 1513.775 234.545 ;
        RECT 1513.930 234.500 1514.250 234.560 ;
        RECT 1513.485 234.360 1514.250 234.500 ;
        RECT 1513.485 234.315 1513.775 234.360 ;
        RECT 1513.930 234.300 1514.250 234.360 ;
        RECT 1513.485 158.000 1513.775 158.045 ;
        RECT 1513.930 158.000 1514.250 158.060 ;
        RECT 1513.485 157.860 1514.250 158.000 ;
        RECT 1513.485 157.815 1513.775 157.860 ;
        RECT 1513.930 157.800 1514.250 157.860 ;
        RECT 1513.930 137.940 1514.250 138.000 ;
        RECT 1513.735 137.800 1514.250 137.940 ;
        RECT 1513.930 137.740 1514.250 137.800 ;
        RECT 1513.930 90.000 1514.250 90.060 ;
        RECT 1513.735 89.860 1514.250 90.000 ;
        RECT 1513.930 89.800 1514.250 89.860 ;
        RECT 1358.450 19.960 1358.770 20.020 ;
        RECT 1513.930 19.960 1514.250 20.020 ;
        RECT 1358.450 19.820 1514.250 19.960 ;
        RECT 1358.450 19.760 1358.770 19.820 ;
        RECT 1513.930 19.760 1514.250 19.820 ;
      LAYER via ;
        RECT 1513.040 1666.380 1513.300 1666.640 ;
        RECT 1515.340 1666.380 1515.600 1666.640 ;
        RECT 1513.040 1641.900 1513.300 1642.160 ;
        RECT 1513.960 1593.960 1514.220 1594.220 ;
        RECT 1513.960 1569.480 1514.220 1569.740 ;
        RECT 1514.880 1569.480 1515.140 1569.740 ;
        RECT 1513.960 1511.000 1514.220 1511.260 ;
        RECT 1513.960 1497.400 1514.220 1497.660 ;
        RECT 1513.040 1435.180 1513.300 1435.440 ;
        RECT 1513.960 1435.180 1514.220 1435.440 ;
        RECT 1513.040 1393.700 1513.300 1393.960 ;
        RECT 1513.960 1393.700 1514.220 1393.960 ;
        RECT 1513.500 1338.620 1513.760 1338.880 ;
        RECT 1513.960 1338.620 1514.220 1338.880 ;
        RECT 1513.040 1159.100 1513.300 1159.360 ;
        RECT 1513.500 1159.100 1513.760 1159.360 ;
        RECT 1513.960 1110.820 1514.220 1111.080 ;
        RECT 1513.500 1110.480 1513.760 1110.740 ;
        RECT 1513.960 1096.540 1514.220 1096.800 ;
        RECT 1514.880 1096.540 1515.140 1096.800 ;
        RECT 1513.500 1028.540 1513.760 1028.800 ;
        RECT 1513.500 1027.860 1513.760 1028.120 ;
        RECT 1513.040 965.980 1513.300 966.240 ;
        RECT 1513.500 965.980 1513.760 966.240 ;
        RECT 1513.960 917.700 1514.220 917.960 ;
        RECT 1515.340 917.700 1515.600 917.960 ;
        RECT 1513.960 883.360 1514.220 883.620 ;
        RECT 1515.340 883.360 1515.600 883.620 ;
        RECT 1513.040 838.140 1513.300 838.400 ;
        RECT 1513.960 838.140 1514.220 838.400 ;
        RECT 1513.040 789.860 1513.300 790.120 ;
        RECT 1513.960 766.060 1514.220 766.320 ;
        RECT 1513.040 717.440 1513.300 717.700 ;
        RECT 1513.500 717.440 1513.760 717.700 ;
        RECT 1513.040 710.300 1513.300 710.560 ;
        RECT 1513.960 710.300 1514.220 710.560 ;
        RECT 1513.960 596.740 1514.220 597.000 ;
        RECT 1513.500 544.720 1513.760 544.980 ;
        RECT 1513.500 523.980 1513.760 524.240 ;
        RECT 1513.960 447.820 1514.220 448.080 ;
        RECT 1513.960 330.860 1514.220 331.120 ;
        RECT 1514.880 330.860 1515.140 331.120 ;
        RECT 1513.960 234.300 1514.220 234.560 ;
        RECT 1513.960 157.800 1514.220 158.060 ;
        RECT 1513.960 137.740 1514.220 138.000 ;
        RECT 1513.960 89.800 1514.220 90.060 ;
        RECT 1358.480 19.760 1358.740 20.020 ;
        RECT 1513.960 19.760 1514.220 20.020 ;
      LAYER met2 ;
        RECT 1516.710 1700.410 1516.990 1704.000 ;
        RECT 1515.400 1700.270 1516.990 1700.410 ;
        RECT 1515.400 1666.670 1515.540 1700.270 ;
        RECT 1516.710 1700.000 1516.990 1700.270 ;
        RECT 1513.040 1666.350 1513.300 1666.670 ;
        RECT 1515.340 1666.350 1515.600 1666.670 ;
        RECT 1513.100 1642.190 1513.240 1666.350 ;
        RECT 1513.040 1641.870 1513.300 1642.190 ;
        RECT 1513.960 1593.930 1514.220 1594.250 ;
        RECT 1514.020 1593.765 1514.160 1593.930 ;
        RECT 1513.950 1593.395 1514.230 1593.765 ;
        RECT 1514.870 1593.395 1515.150 1593.765 ;
        RECT 1514.940 1569.770 1515.080 1593.395 ;
        RECT 1513.960 1569.450 1514.220 1569.770 ;
        RECT 1514.880 1569.450 1515.140 1569.770 ;
        RECT 1514.020 1511.290 1514.160 1569.450 ;
        RECT 1513.960 1510.970 1514.220 1511.290 ;
        RECT 1513.960 1497.370 1514.220 1497.690 ;
        RECT 1514.020 1435.470 1514.160 1497.370 ;
        RECT 1513.040 1435.150 1513.300 1435.470 ;
        RECT 1513.960 1435.150 1514.220 1435.470 ;
        RECT 1513.100 1393.990 1513.240 1435.150 ;
        RECT 1513.040 1393.670 1513.300 1393.990 ;
        RECT 1513.960 1393.670 1514.220 1393.990 ;
        RECT 1514.020 1338.910 1514.160 1393.670 ;
        RECT 1513.500 1338.765 1513.760 1338.910 ;
        RECT 1513.490 1338.395 1513.770 1338.765 ;
        RECT 1513.960 1338.590 1514.220 1338.910 ;
        RECT 1513.030 1289.435 1513.310 1289.805 ;
        RECT 1513.100 1242.205 1513.240 1289.435 ;
        RECT 1513.030 1241.835 1513.310 1242.205 ;
        RECT 1513.950 1241.835 1514.230 1242.205 ;
        RECT 1514.020 1225.090 1514.160 1241.835 ;
        RECT 1513.560 1224.950 1514.160 1225.090 ;
        RECT 1513.560 1173.410 1513.700 1224.950 ;
        RECT 1513.100 1173.270 1513.700 1173.410 ;
        RECT 1513.100 1159.390 1513.240 1173.270 ;
        RECT 1513.040 1159.070 1513.300 1159.390 ;
        RECT 1513.500 1159.070 1513.760 1159.390 ;
        RECT 1513.560 1124.960 1513.700 1159.070 ;
        RECT 1513.560 1124.820 1514.160 1124.960 ;
        RECT 1514.020 1111.110 1514.160 1124.820 ;
        RECT 1513.960 1110.790 1514.220 1111.110 ;
        RECT 1513.500 1110.450 1513.760 1110.770 ;
        RECT 1513.560 1097.250 1513.700 1110.450 ;
        RECT 1513.560 1097.110 1514.160 1097.250 ;
        RECT 1514.020 1096.830 1514.160 1097.110 ;
        RECT 1513.960 1096.510 1514.220 1096.830 ;
        RECT 1514.880 1096.510 1515.140 1096.830 ;
        RECT 1514.940 1049.085 1515.080 1096.510 ;
        RECT 1513.490 1048.715 1513.770 1049.085 ;
        RECT 1514.870 1048.715 1515.150 1049.085 ;
        RECT 1513.560 1028.830 1513.700 1048.715 ;
        RECT 1513.500 1028.510 1513.760 1028.830 ;
        RECT 1513.500 1027.830 1513.760 1028.150 ;
        RECT 1513.560 980.290 1513.700 1027.830 ;
        RECT 1513.100 980.150 1513.700 980.290 ;
        RECT 1513.100 966.270 1513.240 980.150 ;
        RECT 1513.040 965.950 1513.300 966.270 ;
        RECT 1513.500 966.125 1513.760 966.270 ;
        RECT 1513.490 965.755 1513.770 966.125 ;
        RECT 1515.330 965.755 1515.610 966.125 ;
        RECT 1515.400 917.990 1515.540 965.755 ;
        RECT 1513.960 917.845 1514.220 917.990 ;
        RECT 1515.340 917.845 1515.600 917.990 ;
        RECT 1513.950 917.475 1514.230 917.845 ;
        RECT 1515.330 917.475 1515.610 917.845 ;
        RECT 1515.400 883.650 1515.540 917.475 ;
        RECT 1513.960 883.330 1514.220 883.650 ;
        RECT 1515.340 883.330 1515.600 883.650 ;
        RECT 1514.020 838.430 1514.160 883.330 ;
        RECT 1513.040 838.110 1513.300 838.430 ;
        RECT 1513.960 838.110 1514.220 838.430 ;
        RECT 1513.100 790.150 1513.240 838.110 ;
        RECT 1513.040 789.830 1513.300 790.150 ;
        RECT 1513.960 766.030 1514.220 766.350 ;
        RECT 1514.020 717.810 1514.160 766.030 ;
        RECT 1513.560 717.730 1514.160 717.810 ;
        RECT 1513.040 717.410 1513.300 717.730 ;
        RECT 1513.500 717.670 1514.160 717.730 ;
        RECT 1513.500 717.410 1513.760 717.670 ;
        RECT 1513.100 710.590 1513.240 717.410 ;
        RECT 1513.040 710.270 1513.300 710.590 ;
        RECT 1513.960 710.270 1514.220 710.590 ;
        RECT 1514.020 597.030 1514.160 710.270 ;
        RECT 1513.960 596.710 1514.220 597.030 ;
        RECT 1513.500 544.690 1513.760 545.010 ;
        RECT 1513.560 524.270 1513.700 544.690 ;
        RECT 1513.500 523.950 1513.760 524.270 ;
        RECT 1513.960 447.790 1514.220 448.110 ;
        RECT 1514.020 434.365 1514.160 447.790 ;
        RECT 1513.950 433.995 1514.230 434.365 ;
        RECT 1513.490 386.395 1513.770 386.765 ;
        RECT 1513.560 362.170 1513.700 386.395 ;
        RECT 1513.100 362.030 1513.700 362.170 ;
        RECT 1513.100 339.165 1513.240 362.030 ;
        RECT 1513.030 338.795 1513.310 339.165 ;
        RECT 1513.950 338.115 1514.230 338.485 ;
        RECT 1514.020 331.150 1514.160 338.115 ;
        RECT 1513.960 330.830 1514.220 331.150 ;
        RECT 1514.880 330.830 1515.140 331.150 ;
        RECT 1514.940 241.925 1515.080 330.830 ;
        RECT 1513.950 241.555 1514.230 241.925 ;
        RECT 1514.870 241.555 1515.150 241.925 ;
        RECT 1514.020 234.590 1514.160 241.555 ;
        RECT 1513.960 234.270 1514.220 234.590 ;
        RECT 1513.960 157.770 1514.220 158.090 ;
        RECT 1514.020 138.030 1514.160 157.770 ;
        RECT 1513.960 137.710 1514.220 138.030 ;
        RECT 1513.960 89.770 1514.220 90.090 ;
        RECT 1514.020 20.050 1514.160 89.770 ;
        RECT 1358.480 19.730 1358.740 20.050 ;
        RECT 1513.960 19.730 1514.220 20.050 ;
        RECT 1358.540 2.400 1358.680 19.730 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
      LAYER via2 ;
        RECT 1513.950 1593.440 1514.230 1593.720 ;
        RECT 1514.870 1593.440 1515.150 1593.720 ;
        RECT 1513.490 1338.440 1513.770 1338.720 ;
        RECT 1513.030 1289.480 1513.310 1289.760 ;
        RECT 1513.030 1241.880 1513.310 1242.160 ;
        RECT 1513.950 1241.880 1514.230 1242.160 ;
        RECT 1513.490 1048.760 1513.770 1049.040 ;
        RECT 1514.870 1048.760 1515.150 1049.040 ;
        RECT 1513.490 965.800 1513.770 966.080 ;
        RECT 1515.330 965.800 1515.610 966.080 ;
        RECT 1513.950 917.520 1514.230 917.800 ;
        RECT 1515.330 917.520 1515.610 917.800 ;
        RECT 1513.950 434.040 1514.230 434.320 ;
        RECT 1513.490 386.440 1513.770 386.720 ;
        RECT 1513.030 338.840 1513.310 339.120 ;
        RECT 1513.950 338.160 1514.230 338.440 ;
        RECT 1513.950 241.600 1514.230 241.880 ;
        RECT 1514.870 241.600 1515.150 241.880 ;
      LAYER met3 ;
        RECT 1513.925 1593.730 1514.255 1593.745 ;
        RECT 1514.845 1593.730 1515.175 1593.745 ;
        RECT 1513.925 1593.430 1515.175 1593.730 ;
        RECT 1513.925 1593.415 1514.255 1593.430 ;
        RECT 1514.845 1593.415 1515.175 1593.430 ;
        RECT 1513.465 1338.740 1513.795 1338.745 ;
        RECT 1513.465 1338.730 1514.050 1338.740 ;
        RECT 1513.465 1338.430 1514.250 1338.730 ;
        RECT 1513.465 1338.420 1514.050 1338.430 ;
        RECT 1513.465 1338.415 1513.795 1338.420 ;
        RECT 1513.670 1290.140 1514.050 1290.460 ;
        RECT 1513.005 1289.770 1513.335 1289.785 ;
        RECT 1513.710 1289.770 1514.010 1290.140 ;
        RECT 1513.005 1289.470 1514.010 1289.770 ;
        RECT 1513.005 1289.455 1513.335 1289.470 ;
        RECT 1513.005 1242.170 1513.335 1242.185 ;
        RECT 1513.925 1242.170 1514.255 1242.185 ;
        RECT 1513.005 1241.870 1514.255 1242.170 ;
        RECT 1513.005 1241.855 1513.335 1241.870 ;
        RECT 1513.925 1241.855 1514.255 1241.870 ;
        RECT 1513.465 1049.050 1513.795 1049.065 ;
        RECT 1514.845 1049.050 1515.175 1049.065 ;
        RECT 1513.465 1048.750 1515.175 1049.050 ;
        RECT 1513.465 1048.735 1513.795 1048.750 ;
        RECT 1514.845 1048.735 1515.175 1048.750 ;
        RECT 1513.465 966.090 1513.795 966.105 ;
        RECT 1515.305 966.090 1515.635 966.105 ;
        RECT 1513.465 965.790 1515.635 966.090 ;
        RECT 1513.465 965.775 1513.795 965.790 ;
        RECT 1515.305 965.775 1515.635 965.790 ;
        RECT 1513.925 917.810 1514.255 917.825 ;
        RECT 1515.305 917.810 1515.635 917.825 ;
        RECT 1513.925 917.510 1515.635 917.810 ;
        RECT 1513.925 917.495 1514.255 917.510 ;
        RECT 1515.305 917.495 1515.635 917.510 ;
        RECT 1513.925 434.340 1514.255 434.345 ;
        RECT 1513.670 434.330 1514.255 434.340 ;
        RECT 1513.470 434.030 1514.255 434.330 ;
        RECT 1513.670 434.020 1514.255 434.030 ;
        RECT 1513.925 434.015 1514.255 434.020 ;
        RECT 1513.465 386.740 1513.795 386.745 ;
        RECT 1513.465 386.730 1514.050 386.740 ;
        RECT 1513.240 386.430 1514.050 386.730 ;
        RECT 1513.465 386.420 1514.050 386.430 ;
        RECT 1513.465 386.415 1513.795 386.420 ;
        RECT 1513.005 339.130 1513.335 339.145 ;
        RECT 1513.005 338.830 1514.930 339.130 ;
        RECT 1513.005 338.815 1513.335 338.830 ;
        RECT 1513.925 338.450 1514.255 338.465 ;
        RECT 1514.630 338.450 1514.930 338.830 ;
        RECT 1513.925 338.150 1514.930 338.450 ;
        RECT 1513.925 338.135 1514.255 338.150 ;
        RECT 1513.925 241.890 1514.255 241.905 ;
        RECT 1514.845 241.890 1515.175 241.905 ;
        RECT 1513.925 241.590 1515.175 241.890 ;
        RECT 1513.925 241.575 1514.255 241.590 ;
        RECT 1514.845 241.575 1515.175 241.590 ;
      LAYER via3 ;
        RECT 1513.700 1338.420 1514.020 1338.740 ;
        RECT 1513.700 1290.140 1514.020 1290.460 ;
        RECT 1513.700 434.020 1514.020 434.340 ;
        RECT 1513.700 386.420 1514.020 386.740 ;
      LAYER met4 ;
        RECT 1513.695 1338.415 1514.025 1338.745 ;
        RECT 1513.710 1290.465 1514.010 1338.415 ;
        RECT 1513.695 1290.135 1514.025 1290.465 ;
        RECT 1513.695 434.015 1514.025 434.345 ;
        RECT 1513.710 386.745 1514.010 434.015 ;
        RECT 1513.695 386.415 1514.025 386.745 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 0.300 ;
=======
      LAYER met1 ;
        RECT 1518.530 1678.480 1518.850 1678.540 ;
        RECT 1520.370 1678.480 1520.690 1678.540 ;
        RECT 1518.530 1678.340 1520.690 1678.480 ;
        RECT 1518.530 1678.280 1518.850 1678.340 ;
        RECT 1520.370 1678.280 1520.690 1678.340 ;
        RECT 1376.390 16.900 1376.710 16.960 ;
        RECT 1376.390 16.760 1487.020 16.900 ;
        RECT 1376.390 16.700 1376.710 16.760 ;
        RECT 1486.880 16.560 1487.020 16.760 ;
        RECT 1518.070 16.560 1518.390 16.620 ;
        RECT 1486.880 16.420 1518.390 16.560 ;
        RECT 1518.070 16.360 1518.390 16.420 ;
      LAYER via ;
        RECT 1518.560 1678.280 1518.820 1678.540 ;
        RECT 1520.400 1678.280 1520.660 1678.540 ;
        RECT 1376.420 16.700 1376.680 16.960 ;
        RECT 1518.100 16.360 1518.360 16.620 ;
      LAYER met2 ;
        RECT 1521.310 1700.410 1521.590 1704.000 ;
        RECT 1520.460 1700.270 1521.590 1700.410 ;
        RECT 1520.460 1678.570 1520.600 1700.270 ;
        RECT 1521.310 1700.000 1521.590 1700.270 ;
        RECT 1518.560 1678.250 1518.820 1678.570 ;
        RECT 1520.400 1678.250 1520.660 1678.570 ;
        RECT 1518.620 20.810 1518.760 1678.250 ;
        RECT 1518.160 20.670 1518.760 20.810 ;
        RECT 1376.420 16.670 1376.680 16.990 ;
        RECT 1376.480 2.400 1376.620 16.670 ;
        RECT 1518.160 16.650 1518.300 20.670 ;
        RECT 1518.100 16.330 1518.360 16.650 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 0.300 ;
=======
      LAYER li1 ;
        RECT 1486.405 1685.465 1486.575 1686.315 ;
      LAYER mcon ;
        RECT 1486.405 1686.145 1486.575 1686.315 ;
      LAYER met1 ;
        RECT 1400.310 1686.300 1400.630 1686.360 ;
        RECT 1486.345 1686.300 1486.635 1686.345 ;
        RECT 1400.310 1686.160 1486.635 1686.300 ;
        RECT 1400.310 1686.100 1400.630 1686.160 ;
        RECT 1486.345 1686.115 1486.635 1686.160 ;
        RECT 1486.345 1685.620 1486.635 1685.665 ;
        RECT 1526.350 1685.620 1526.670 1685.680 ;
        RECT 1486.345 1685.480 1526.670 1685.620 ;
        RECT 1486.345 1685.435 1486.635 1685.480 ;
        RECT 1526.350 1685.420 1526.670 1685.480 ;
        RECT 1394.330 16.560 1394.650 16.620 ;
        RECT 1400.310 16.560 1400.630 16.620 ;
        RECT 1394.330 16.420 1400.630 16.560 ;
        RECT 1394.330 16.360 1394.650 16.420 ;
        RECT 1400.310 16.360 1400.630 16.420 ;
      LAYER via ;
        RECT 1400.340 1686.100 1400.600 1686.360 ;
        RECT 1526.380 1685.420 1526.640 1685.680 ;
        RECT 1394.360 16.360 1394.620 16.620 ;
        RECT 1400.340 16.360 1400.600 16.620 ;
      LAYER met2 ;
        RECT 1526.370 1700.000 1526.650 1704.000 ;
        RECT 1400.340 1686.070 1400.600 1686.390 ;
        RECT 1400.400 16.650 1400.540 1686.070 ;
        RECT 1526.440 1685.710 1526.580 1700.000 ;
        RECT 1526.380 1685.390 1526.640 1685.710 ;
        RECT 1394.360 16.330 1394.620 16.650 ;
        RECT 1400.340 16.330 1400.600 16.650 ;
        RECT 1394.420 2.400 1394.560 16.330 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 0.300 ;
=======
      LAYER li1 ;
        RECT 1486.865 15.725 1487.035 19.295 ;
      LAYER mcon ;
        RECT 1486.865 19.125 1487.035 19.295 ;
      LAYER met1 ;
        RECT 1525.430 1678.140 1525.750 1678.200 ;
        RECT 1530.030 1678.140 1530.350 1678.200 ;
        RECT 1525.430 1678.000 1530.350 1678.140 ;
        RECT 1525.430 1677.940 1525.750 1678.000 ;
        RECT 1530.030 1677.940 1530.350 1678.000 ;
        RECT 1486.805 19.280 1487.095 19.325 ;
        RECT 1525.430 19.280 1525.750 19.340 ;
        RECT 1486.805 19.140 1525.750 19.280 ;
        RECT 1486.805 19.095 1487.095 19.140 ;
        RECT 1525.430 19.080 1525.750 19.140 ;
        RECT 1486.805 15.880 1487.095 15.925 ;
        RECT 1438.580 15.740 1487.095 15.880 ;
        RECT 1412.270 14.860 1412.590 14.920 ;
        RECT 1438.580 14.860 1438.720 15.740 ;
        RECT 1486.805 15.695 1487.095 15.740 ;
        RECT 1412.270 14.720 1438.720 14.860 ;
        RECT 1412.270 14.660 1412.590 14.720 ;
      LAYER via ;
        RECT 1525.460 1677.940 1525.720 1678.200 ;
        RECT 1530.060 1677.940 1530.320 1678.200 ;
        RECT 1525.460 19.080 1525.720 19.340 ;
        RECT 1412.300 14.660 1412.560 14.920 ;
      LAYER met2 ;
        RECT 1530.970 1700.410 1531.250 1704.000 ;
        RECT 1530.120 1700.270 1531.250 1700.410 ;
        RECT 1530.120 1678.230 1530.260 1700.270 ;
        RECT 1530.970 1700.000 1531.250 1700.270 ;
        RECT 1525.460 1677.910 1525.720 1678.230 ;
        RECT 1530.060 1677.910 1530.320 1678.230 ;
        RECT 1525.520 19.370 1525.660 1677.910 ;
        RECT 1525.460 19.050 1525.720 19.370 ;
        RECT 1412.300 14.630 1412.560 14.950 ;
        RECT 1412.360 2.400 1412.500 14.630 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 0.300 ;
=======
      LAYER li1 ;
        RECT 1533.785 1449.165 1533.955 1497.275 ;
        RECT 1533.325 496.485 1533.495 531.335 ;
        RECT 1533.325 338.045 1533.495 386.155 ;
        RECT 1533.325 241.485 1533.495 289.595 ;
        RECT 1533.325 89.845 1533.495 137.955 ;
      LAYER mcon ;
        RECT 1533.785 1497.105 1533.955 1497.275 ;
        RECT 1533.325 531.165 1533.495 531.335 ;
        RECT 1533.325 385.985 1533.495 386.155 ;
        RECT 1533.325 289.425 1533.495 289.595 ;
        RECT 1533.325 137.785 1533.495 137.955 ;
      LAYER met1 ;
        RECT 1533.710 1607.900 1534.030 1608.160 ;
        RECT 1533.800 1607.420 1533.940 1607.900 ;
        RECT 1534.170 1607.420 1534.490 1607.480 ;
        RECT 1533.800 1607.280 1534.490 1607.420 ;
        RECT 1534.170 1607.220 1534.490 1607.280 ;
        RECT 1532.330 1593.820 1532.650 1593.880 ;
        RECT 1534.170 1593.820 1534.490 1593.880 ;
        RECT 1532.330 1593.680 1534.490 1593.820 ;
        RECT 1532.330 1593.620 1532.650 1593.680 ;
        RECT 1534.170 1593.620 1534.490 1593.680 ;
        RECT 1532.330 1545.540 1532.650 1545.600 ;
        RECT 1532.790 1545.540 1533.110 1545.600 ;
        RECT 1532.330 1545.400 1533.110 1545.540 ;
        RECT 1532.330 1545.340 1532.650 1545.400 ;
        RECT 1532.790 1545.340 1533.110 1545.400 ;
        RECT 1533.725 1497.260 1534.015 1497.305 ;
        RECT 1534.170 1497.260 1534.490 1497.320 ;
        RECT 1533.725 1497.120 1534.490 1497.260 ;
        RECT 1533.725 1497.075 1534.015 1497.120 ;
        RECT 1534.170 1497.060 1534.490 1497.120 ;
        RECT 1533.710 1449.320 1534.030 1449.380 ;
        RECT 1533.515 1449.180 1534.030 1449.320 ;
        RECT 1533.710 1449.120 1534.030 1449.180 ;
        RECT 1532.790 1414.640 1533.110 1414.700 ;
        RECT 1533.710 1414.640 1534.030 1414.700 ;
        RECT 1532.790 1414.500 1534.030 1414.640 ;
        RECT 1532.790 1414.440 1533.110 1414.500 ;
        RECT 1533.710 1414.440 1534.030 1414.500 ;
        RECT 1532.790 1318.080 1533.110 1318.140 ;
        RECT 1533.710 1318.080 1534.030 1318.140 ;
        RECT 1532.790 1317.940 1534.030 1318.080 ;
        RECT 1532.790 1317.880 1533.110 1317.940 ;
        RECT 1533.710 1317.880 1534.030 1317.940 ;
        RECT 1532.790 1221.520 1533.110 1221.580 ;
        RECT 1533.710 1221.520 1534.030 1221.580 ;
        RECT 1532.790 1221.380 1534.030 1221.520 ;
        RECT 1532.790 1221.320 1533.110 1221.380 ;
        RECT 1533.710 1221.320 1534.030 1221.380 ;
        RECT 1532.790 1124.960 1533.110 1125.020 ;
        RECT 1533.710 1124.960 1534.030 1125.020 ;
        RECT 1532.790 1124.820 1534.030 1124.960 ;
        RECT 1532.790 1124.760 1533.110 1124.820 ;
        RECT 1533.710 1124.760 1534.030 1124.820 ;
        RECT 1532.790 1028.400 1533.110 1028.460 ;
        RECT 1533.710 1028.400 1534.030 1028.460 ;
        RECT 1532.790 1028.260 1534.030 1028.400 ;
        RECT 1532.790 1028.200 1533.110 1028.260 ;
        RECT 1533.710 1028.200 1534.030 1028.260 ;
        RECT 1532.790 931.840 1533.110 931.900 ;
        RECT 1533.710 931.840 1534.030 931.900 ;
        RECT 1532.790 931.700 1534.030 931.840 ;
        RECT 1532.790 931.640 1533.110 931.700 ;
        RECT 1533.710 931.640 1534.030 931.700 ;
        RECT 1533.250 883.360 1533.570 883.620 ;
        RECT 1533.340 882.880 1533.480 883.360 ;
        RECT 1533.710 882.880 1534.030 882.940 ;
        RECT 1533.340 882.740 1534.030 882.880 ;
        RECT 1533.710 882.680 1534.030 882.740 ;
        RECT 1532.790 835.280 1533.110 835.340 ;
        RECT 1533.710 835.280 1534.030 835.340 ;
        RECT 1532.790 835.140 1534.030 835.280 ;
        RECT 1532.790 835.080 1533.110 835.140 ;
        RECT 1533.710 835.080 1534.030 835.140 ;
        RECT 1532.790 738.380 1533.110 738.440 ;
        RECT 1533.710 738.380 1534.030 738.440 ;
        RECT 1532.790 738.240 1534.030 738.380 ;
        RECT 1532.790 738.180 1533.110 738.240 ;
        RECT 1533.710 738.180 1534.030 738.240 ;
        RECT 1533.250 689.900 1533.570 690.160 ;
        RECT 1533.340 689.760 1533.480 689.900 ;
        RECT 1533.710 689.760 1534.030 689.820 ;
        RECT 1533.340 689.620 1534.030 689.760 ;
        RECT 1533.710 689.560 1534.030 689.620 ;
        RECT 1532.790 641.820 1533.110 641.880 ;
        RECT 1533.710 641.820 1534.030 641.880 ;
        RECT 1532.790 641.680 1534.030 641.820 ;
        RECT 1532.790 641.620 1533.110 641.680 ;
        RECT 1533.710 641.620 1534.030 641.680 ;
        RECT 1533.250 593.340 1533.570 593.600 ;
        RECT 1533.340 593.200 1533.480 593.340 ;
        RECT 1533.710 593.200 1534.030 593.260 ;
        RECT 1533.340 593.060 1534.030 593.200 ;
        RECT 1533.710 593.000 1534.030 593.060 ;
        RECT 1532.790 545.260 1533.110 545.320 ;
        RECT 1533.710 545.260 1534.030 545.320 ;
        RECT 1532.790 545.120 1534.030 545.260 ;
        RECT 1532.790 545.060 1533.110 545.120 ;
        RECT 1533.710 545.060 1534.030 545.120 ;
        RECT 1533.250 531.320 1533.570 531.380 ;
        RECT 1533.055 531.180 1533.570 531.320 ;
        RECT 1533.250 531.120 1533.570 531.180 ;
        RECT 1533.250 496.640 1533.570 496.700 ;
        RECT 1533.055 496.500 1533.570 496.640 ;
        RECT 1533.250 496.440 1533.570 496.500 ;
        RECT 1532.790 448.700 1533.110 448.760 ;
        RECT 1533.710 448.700 1534.030 448.760 ;
        RECT 1532.790 448.560 1534.030 448.700 ;
        RECT 1532.790 448.500 1533.110 448.560 ;
        RECT 1533.710 448.500 1534.030 448.560 ;
        RECT 1533.250 400.220 1533.570 400.480 ;
        RECT 1533.340 399.740 1533.480 400.220 ;
        RECT 1533.710 399.740 1534.030 399.800 ;
        RECT 1533.340 399.600 1534.030 399.740 ;
        RECT 1533.710 399.540 1534.030 399.600 ;
        RECT 1533.265 386.140 1533.555 386.185 ;
        RECT 1533.710 386.140 1534.030 386.200 ;
        RECT 1533.265 386.000 1534.030 386.140 ;
        RECT 1533.265 385.955 1533.555 386.000 ;
        RECT 1533.710 385.940 1534.030 386.000 ;
        RECT 1533.250 338.200 1533.570 338.260 ;
        RECT 1533.055 338.060 1533.570 338.200 ;
        RECT 1533.250 338.000 1533.570 338.060 ;
        RECT 1533.265 289.580 1533.555 289.625 ;
        RECT 1533.710 289.580 1534.030 289.640 ;
        RECT 1533.265 289.440 1534.030 289.580 ;
        RECT 1533.265 289.395 1533.555 289.440 ;
        RECT 1533.710 289.380 1534.030 289.440 ;
        RECT 1533.250 241.640 1533.570 241.700 ;
        RECT 1533.055 241.500 1533.570 241.640 ;
        RECT 1533.250 241.440 1533.570 241.500 ;
        RECT 1533.250 145.080 1533.570 145.140 ;
        RECT 1534.170 145.080 1534.490 145.140 ;
        RECT 1533.250 144.940 1534.490 145.080 ;
        RECT 1533.250 144.880 1533.570 144.940 ;
        RECT 1534.170 144.880 1534.490 144.940 ;
        RECT 1533.250 137.940 1533.570 138.000 ;
        RECT 1533.055 137.800 1533.570 137.940 ;
        RECT 1533.250 137.740 1533.570 137.800 ;
        RECT 1533.250 90.000 1533.570 90.060 ;
        RECT 1533.055 89.860 1533.570 90.000 ;
        RECT 1533.250 89.800 1533.570 89.860 ;
        RECT 1532.330 15.540 1532.650 15.600 ;
        RECT 1439.040 15.400 1532.650 15.540 ;
        RECT 1429.750 14.520 1430.070 14.580 ;
        RECT 1439.040 14.520 1439.180 15.400 ;
        RECT 1532.330 15.340 1532.650 15.400 ;
        RECT 1429.750 14.380 1439.180 14.520 ;
        RECT 1429.750 14.320 1430.070 14.380 ;
      LAYER via ;
        RECT 1533.740 1607.900 1534.000 1608.160 ;
        RECT 1534.200 1607.220 1534.460 1607.480 ;
        RECT 1532.360 1593.620 1532.620 1593.880 ;
        RECT 1534.200 1593.620 1534.460 1593.880 ;
        RECT 1532.360 1545.340 1532.620 1545.600 ;
        RECT 1532.820 1545.340 1533.080 1545.600 ;
        RECT 1534.200 1497.060 1534.460 1497.320 ;
        RECT 1533.740 1449.120 1534.000 1449.380 ;
        RECT 1532.820 1414.440 1533.080 1414.700 ;
        RECT 1533.740 1414.440 1534.000 1414.700 ;
        RECT 1532.820 1317.880 1533.080 1318.140 ;
        RECT 1533.740 1317.880 1534.000 1318.140 ;
        RECT 1532.820 1221.320 1533.080 1221.580 ;
        RECT 1533.740 1221.320 1534.000 1221.580 ;
        RECT 1532.820 1124.760 1533.080 1125.020 ;
        RECT 1533.740 1124.760 1534.000 1125.020 ;
        RECT 1532.820 1028.200 1533.080 1028.460 ;
        RECT 1533.740 1028.200 1534.000 1028.460 ;
        RECT 1532.820 931.640 1533.080 931.900 ;
        RECT 1533.740 931.640 1534.000 931.900 ;
        RECT 1533.280 883.360 1533.540 883.620 ;
        RECT 1533.740 882.680 1534.000 882.940 ;
        RECT 1532.820 835.080 1533.080 835.340 ;
        RECT 1533.740 835.080 1534.000 835.340 ;
        RECT 1532.820 738.180 1533.080 738.440 ;
        RECT 1533.740 738.180 1534.000 738.440 ;
        RECT 1533.280 689.900 1533.540 690.160 ;
        RECT 1533.740 689.560 1534.000 689.820 ;
        RECT 1532.820 641.620 1533.080 641.880 ;
        RECT 1533.740 641.620 1534.000 641.880 ;
        RECT 1533.280 593.340 1533.540 593.600 ;
        RECT 1533.740 593.000 1534.000 593.260 ;
        RECT 1532.820 545.060 1533.080 545.320 ;
        RECT 1533.740 545.060 1534.000 545.320 ;
        RECT 1533.280 531.120 1533.540 531.380 ;
        RECT 1533.280 496.440 1533.540 496.700 ;
        RECT 1532.820 448.500 1533.080 448.760 ;
        RECT 1533.740 448.500 1534.000 448.760 ;
        RECT 1533.280 400.220 1533.540 400.480 ;
        RECT 1533.740 399.540 1534.000 399.800 ;
        RECT 1533.740 385.940 1534.000 386.200 ;
        RECT 1533.280 338.000 1533.540 338.260 ;
        RECT 1533.740 289.380 1534.000 289.640 ;
        RECT 1533.280 241.440 1533.540 241.700 ;
        RECT 1533.280 144.880 1533.540 145.140 ;
        RECT 1534.200 144.880 1534.460 145.140 ;
        RECT 1533.280 137.740 1533.540 138.000 ;
        RECT 1533.280 89.800 1533.540 90.060 ;
        RECT 1429.780 14.320 1430.040 14.580 ;
        RECT 1532.360 15.340 1532.620 15.600 ;
      LAYER met2 ;
        RECT 1536.030 1700.410 1536.310 1704.000 ;
        RECT 1535.180 1700.270 1536.310 1700.410 ;
        RECT 1535.180 1666.410 1535.320 1700.270 ;
        RECT 1536.030 1700.000 1536.310 1700.270 ;
        RECT 1533.800 1666.270 1535.320 1666.410 ;
        RECT 1533.800 1608.190 1533.940 1666.270 ;
        RECT 1533.740 1607.870 1534.000 1608.190 ;
        RECT 1534.200 1607.190 1534.460 1607.510 ;
        RECT 1534.260 1593.910 1534.400 1607.190 ;
        RECT 1532.360 1593.590 1532.620 1593.910 ;
        RECT 1534.200 1593.590 1534.460 1593.910 ;
        RECT 1532.420 1545.630 1532.560 1593.590 ;
        RECT 1532.360 1545.310 1532.620 1545.630 ;
        RECT 1532.820 1545.310 1533.080 1545.630 ;
        RECT 1532.880 1497.770 1533.020 1545.310 ;
        RECT 1532.880 1497.630 1534.400 1497.770 ;
        RECT 1534.260 1497.350 1534.400 1497.630 ;
        RECT 1534.200 1497.030 1534.460 1497.350 ;
        RECT 1533.740 1449.090 1534.000 1449.410 ;
        RECT 1533.800 1414.730 1533.940 1449.090 ;
        RECT 1532.820 1414.410 1533.080 1414.730 ;
        RECT 1533.740 1414.410 1534.000 1414.730 ;
        RECT 1532.880 1414.130 1533.020 1414.410 ;
        RECT 1532.880 1413.990 1533.480 1414.130 ;
        RECT 1533.340 1366.530 1533.480 1413.990 ;
        RECT 1533.340 1366.390 1533.940 1366.530 ;
        RECT 1533.800 1318.170 1533.940 1366.390 ;
        RECT 1532.820 1317.850 1533.080 1318.170 ;
        RECT 1533.740 1317.850 1534.000 1318.170 ;
        RECT 1532.880 1317.570 1533.020 1317.850 ;
        RECT 1532.880 1317.430 1533.480 1317.570 ;
        RECT 1533.340 1269.970 1533.480 1317.430 ;
        RECT 1533.340 1269.830 1533.940 1269.970 ;
        RECT 1533.800 1221.610 1533.940 1269.830 ;
        RECT 1532.820 1221.290 1533.080 1221.610 ;
        RECT 1533.740 1221.290 1534.000 1221.610 ;
        RECT 1532.880 1221.010 1533.020 1221.290 ;
        RECT 1532.880 1220.870 1533.480 1221.010 ;
        RECT 1533.340 1173.410 1533.480 1220.870 ;
        RECT 1533.340 1173.270 1533.940 1173.410 ;
        RECT 1533.800 1125.050 1533.940 1173.270 ;
        RECT 1532.820 1124.730 1533.080 1125.050 ;
        RECT 1533.740 1124.730 1534.000 1125.050 ;
        RECT 1532.880 1124.450 1533.020 1124.730 ;
        RECT 1532.880 1124.310 1533.480 1124.450 ;
        RECT 1533.340 1076.850 1533.480 1124.310 ;
        RECT 1533.340 1076.710 1533.940 1076.850 ;
        RECT 1533.800 1028.490 1533.940 1076.710 ;
        RECT 1532.820 1028.170 1533.080 1028.490 ;
        RECT 1533.740 1028.170 1534.000 1028.490 ;
        RECT 1532.880 1027.890 1533.020 1028.170 ;
        RECT 1532.880 1027.750 1533.480 1027.890 ;
        RECT 1533.340 980.290 1533.480 1027.750 ;
        RECT 1533.340 980.150 1533.940 980.290 ;
        RECT 1533.800 931.930 1533.940 980.150 ;
        RECT 1532.820 931.610 1533.080 931.930 ;
        RECT 1533.740 931.610 1534.000 931.930 ;
        RECT 1532.880 931.330 1533.020 931.610 ;
        RECT 1532.880 931.190 1533.480 931.330 ;
        RECT 1533.340 883.650 1533.480 931.190 ;
        RECT 1533.280 883.330 1533.540 883.650 ;
        RECT 1533.740 882.650 1534.000 882.970 ;
        RECT 1533.800 835.370 1533.940 882.650 ;
        RECT 1532.820 835.050 1533.080 835.370 ;
        RECT 1533.740 835.050 1534.000 835.370 ;
        RECT 1532.880 834.770 1533.020 835.050 ;
        RECT 1532.880 834.630 1533.480 834.770 ;
        RECT 1533.340 796.690 1533.480 834.630 ;
        RECT 1533.340 796.550 1533.940 796.690 ;
        RECT 1533.800 738.470 1533.940 796.550 ;
        RECT 1532.820 738.210 1533.080 738.470 ;
        RECT 1532.820 738.150 1533.480 738.210 ;
        RECT 1533.740 738.150 1534.000 738.470 ;
        RECT 1532.880 738.070 1533.480 738.150 ;
        RECT 1533.340 690.190 1533.480 738.070 ;
        RECT 1533.280 689.870 1533.540 690.190 ;
        RECT 1533.740 689.530 1534.000 689.850 ;
        RECT 1533.800 641.910 1533.940 689.530 ;
        RECT 1532.820 641.650 1533.080 641.910 ;
        RECT 1532.820 641.590 1533.480 641.650 ;
        RECT 1533.740 641.590 1534.000 641.910 ;
        RECT 1532.880 641.510 1533.480 641.590 ;
        RECT 1533.340 593.630 1533.480 641.510 ;
        RECT 1533.280 593.310 1533.540 593.630 ;
        RECT 1533.740 592.970 1534.000 593.290 ;
        RECT 1533.800 545.350 1533.940 592.970 ;
        RECT 1532.820 545.090 1533.080 545.350 ;
        RECT 1532.820 545.030 1533.480 545.090 ;
        RECT 1533.740 545.030 1534.000 545.350 ;
        RECT 1532.880 544.950 1533.480 545.030 ;
        RECT 1533.340 531.410 1533.480 544.950 ;
        RECT 1533.280 531.090 1533.540 531.410 ;
        RECT 1533.280 496.410 1533.540 496.730 ;
        RECT 1533.340 483.210 1533.480 496.410 ;
        RECT 1533.340 483.070 1533.940 483.210 ;
        RECT 1533.800 448.790 1533.940 483.070 ;
        RECT 1532.820 448.530 1533.080 448.790 ;
        RECT 1532.820 448.470 1533.480 448.530 ;
        RECT 1533.740 448.470 1534.000 448.790 ;
        RECT 1532.880 448.390 1533.480 448.470 ;
        RECT 1533.340 400.510 1533.480 448.390 ;
        RECT 1533.280 400.190 1533.540 400.510 ;
        RECT 1533.740 399.510 1534.000 399.830 ;
        RECT 1533.800 386.230 1533.940 399.510 ;
        RECT 1533.740 385.910 1534.000 386.230 ;
        RECT 1533.280 337.970 1533.540 338.290 ;
        RECT 1533.340 303.690 1533.480 337.970 ;
        RECT 1533.340 303.550 1533.940 303.690 ;
        RECT 1533.800 289.670 1533.940 303.550 ;
        RECT 1533.740 289.350 1534.000 289.670 ;
        RECT 1533.280 241.410 1533.540 241.730 ;
        RECT 1533.340 207.130 1533.480 241.410 ;
        RECT 1533.340 206.990 1533.940 207.130 ;
        RECT 1533.800 168.370 1533.940 206.990 ;
        RECT 1533.800 168.230 1534.400 168.370 ;
        RECT 1534.260 145.170 1534.400 168.230 ;
        RECT 1533.280 144.850 1533.540 145.170 ;
        RECT 1534.200 144.850 1534.460 145.170 ;
        RECT 1533.340 138.030 1533.480 144.850 ;
        RECT 1533.280 137.710 1533.540 138.030 ;
        RECT 1533.280 89.770 1533.540 90.090 ;
        RECT 1533.340 62.290 1533.480 89.770 ;
        RECT 1532.420 62.150 1533.480 62.290 ;
        RECT 1532.420 15.630 1532.560 62.150 ;
        RECT 1532.360 15.310 1532.620 15.630 ;
        RECT 1429.780 14.290 1430.040 14.610 ;
        RECT 1429.840 2.400 1429.980 14.290 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 0.300 ;
=======
      LAYER met1 ;
        RECT 1447.690 15.200 1448.010 15.260 ;
        RECT 1540.150 15.200 1540.470 15.260 ;
        RECT 1447.690 15.060 1540.470 15.200 ;
        RECT 1447.690 15.000 1448.010 15.060 ;
        RECT 1540.150 15.000 1540.470 15.060 ;
      LAYER via ;
        RECT 1447.720 15.000 1447.980 15.260 ;
        RECT 1540.180 15.000 1540.440 15.260 ;
      LAYER met2 ;
        RECT 1540.630 1700.410 1540.910 1704.000 ;
        RECT 1540.240 1700.270 1540.910 1700.410 ;
        RECT 1540.240 15.290 1540.380 1700.270 ;
        RECT 1540.630 1700.000 1540.910 1700.270 ;
        RECT 1447.720 14.970 1447.980 15.290 ;
        RECT 1540.180 14.970 1540.440 15.290 ;
        RECT 1447.780 2.400 1447.920 14.970 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 0.300 ;
=======
      LAYER li1 ;
        RECT 1488.245 16.065 1488.415 17.255 ;
      LAYER mcon ;
        RECT 1488.245 17.085 1488.415 17.255 ;
      LAYER met1 ;
        RECT 1488.185 17.240 1488.475 17.285 ;
        RECT 1546.130 17.240 1546.450 17.300 ;
        RECT 1488.185 17.100 1546.450 17.240 ;
        RECT 1488.185 17.055 1488.475 17.100 ;
        RECT 1546.130 17.040 1546.450 17.100 ;
        RECT 1465.630 16.220 1465.950 16.280 ;
        RECT 1488.185 16.220 1488.475 16.265 ;
        RECT 1465.630 16.080 1488.475 16.220 ;
        RECT 1465.630 16.020 1465.950 16.080 ;
        RECT 1488.185 16.035 1488.475 16.080 ;
      LAYER via ;
        RECT 1546.160 17.040 1546.420 17.300 ;
        RECT 1465.660 16.020 1465.920 16.280 ;
      LAYER met2 ;
        RECT 1545.690 1700.410 1545.970 1704.000 ;
        RECT 1545.690 1700.270 1546.360 1700.410 ;
        RECT 1545.690 1700.000 1545.970 1700.270 ;
        RECT 1546.220 17.330 1546.360 1700.270 ;
        RECT 1546.160 17.010 1546.420 17.330 ;
        RECT 1465.660 15.990 1465.920 16.310 ;
        RECT 1465.720 2.400 1465.860 15.990 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1546.590 1678.140 1546.910 1678.200 ;
        RECT 1549.350 1678.140 1549.670 1678.200 ;
        RECT 1546.590 1678.000 1549.670 1678.140 ;
        RECT 1546.590 1677.940 1546.910 1678.000 ;
        RECT 1549.350 1677.940 1549.670 1678.000 ;
        RECT 1484.490 17.240 1484.810 17.300 ;
        RECT 1484.490 17.100 1487.940 17.240 ;
        RECT 1484.490 17.040 1484.810 17.100 ;
        RECT 1487.800 16.900 1487.940 17.100 ;
        RECT 1487.800 16.760 1528.880 16.900 ;
        RECT 1528.740 16.560 1528.880 16.760 ;
        RECT 1546.590 16.560 1546.910 16.620 ;
        RECT 1528.740 16.420 1546.910 16.560 ;
        RECT 1546.590 16.360 1546.910 16.420 ;
      LAYER via ;
        RECT 1546.620 1677.940 1546.880 1678.200 ;
        RECT 1549.380 1677.940 1549.640 1678.200 ;
        RECT 1484.520 17.040 1484.780 17.300 ;
        RECT 1546.620 16.360 1546.880 16.620 ;
      LAYER met2 ;
        RECT 1550.290 1700.410 1550.570 1704.000 ;
        RECT 1549.440 1700.270 1550.570 1700.410 ;
        RECT 1549.440 1678.230 1549.580 1700.270 ;
        RECT 1550.290 1700.000 1550.570 1700.270 ;
        RECT 1546.620 1677.910 1546.880 1678.230 ;
        RECT 1549.380 1677.910 1549.640 1678.230 ;
        RECT 1484.520 17.010 1484.780 17.330 ;
        RECT 1484.580 9.250 1484.720 17.010 ;
        RECT 1546.680 16.650 1546.820 1677.910 ;
        RECT 1546.620 16.330 1546.880 16.650 ;
        RECT 1483.660 9.110 1484.720 9.250 ;
        RECT 1483.660 2.400 1483.800 9.110 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 0.300 ;
=======
      LAYER met1 ;
        RECT 1501.510 18.260 1501.830 18.320 ;
        RECT 1553.950 18.260 1554.270 18.320 ;
        RECT 1501.510 18.120 1554.270 18.260 ;
        RECT 1501.510 18.060 1501.830 18.120 ;
        RECT 1553.950 18.060 1554.270 18.120 ;
      LAYER via ;
        RECT 1501.540 18.060 1501.800 18.320 ;
        RECT 1553.980 18.060 1554.240 18.320 ;
      LAYER met2 ;
        RECT 1554.890 1700.410 1555.170 1704.000 ;
        RECT 1554.040 1700.270 1555.170 1700.410 ;
        RECT 1554.040 18.350 1554.180 1700.270 ;
        RECT 1554.890 1700.000 1555.170 1700.270 ;
        RECT 1501.540 18.030 1501.800 18.350 ;
        RECT 1553.980 18.030 1554.240 18.350 ;
        RECT 1501.600 2.400 1501.740 18.030 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1560.390 96.940 1560.710 97.200 ;
        RECT 1560.480 96.520 1560.620 96.940 ;
        RECT 1560.390 96.260 1560.710 96.520 ;
        RECT 1518.990 19.620 1519.310 19.680 ;
        RECT 1560.390 19.620 1560.710 19.680 ;
        RECT 1518.990 19.480 1560.710 19.620 ;
        RECT 1518.990 19.420 1519.310 19.480 ;
        RECT 1560.390 19.420 1560.710 19.480 ;
      LAYER via ;
        RECT 1560.420 96.940 1560.680 97.200 ;
        RECT 1560.420 96.260 1560.680 96.520 ;
        RECT 1519.020 19.420 1519.280 19.680 ;
        RECT 1560.420 19.420 1560.680 19.680 ;
      LAYER met2 ;
        RECT 1559.950 1700.410 1560.230 1704.000 ;
        RECT 1559.950 1700.270 1560.620 1700.410 ;
        RECT 1559.950 1700.000 1560.230 1700.270 ;
        RECT 1560.480 97.230 1560.620 1700.270 ;
        RECT 1560.420 96.910 1560.680 97.230 ;
        RECT 1560.420 96.230 1560.680 96.550 ;
        RECT 1560.480 19.710 1560.620 96.230 ;
        RECT 1519.020 19.390 1519.280 19.710 ;
        RECT 1560.420 19.390 1560.680 19.710 ;
        RECT 1519.080 2.400 1519.220 19.390 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1339.130 1677.460 1339.450 1677.520 ;
        RECT 1341.890 1677.460 1342.210 1677.520 ;
        RECT 1339.130 1677.320 1342.210 1677.460 ;
        RECT 1339.130 1677.260 1339.450 1677.320 ;
        RECT 1341.890 1677.260 1342.210 1677.320 ;
        RECT 716.290 47.160 716.610 47.220 ;
        RECT 1339.130 47.160 1339.450 47.220 ;
        RECT 716.290 47.020 1339.450 47.160 ;
        RECT 716.290 46.960 716.610 47.020 ;
        RECT 1339.130 46.960 1339.450 47.020 ;
      LAYER via ;
        RECT 1339.160 1677.260 1339.420 1677.520 ;
        RECT 1341.920 1677.260 1342.180 1677.520 ;
        RECT 716.320 46.960 716.580 47.220 ;
        RECT 1339.160 46.960 1339.420 47.220 ;
      LAYER met2 ;
        RECT 1343.290 1700.410 1343.570 1704.000 ;
        RECT 1341.980 1700.270 1343.570 1700.410 ;
        RECT 1341.980 1677.550 1342.120 1700.270 ;
        RECT 1343.290 1700.000 1343.570 1700.270 ;
        RECT 1339.160 1677.230 1339.420 1677.550 ;
        RECT 1341.920 1677.230 1342.180 1677.550 ;
        RECT 1339.220 47.250 1339.360 1677.230 ;
        RECT 716.320 46.930 716.580 47.250 ;
        RECT 1339.160 46.930 1339.420 47.250 ;
        RECT 716.380 2.400 716.520 46.930 ;
        RECT 716.170 -4.800 716.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 0.300 ;
=======
      LAYER li1 ;
        RECT 1562.305 1490.645 1562.475 1529.915 ;
        RECT 1561.845 1200.625 1562.015 1248.735 ;
        RECT 1561.845 689.605 1562.015 724.455 ;
        RECT 1561.845 593.045 1562.015 627.895 ;
        RECT 1561.845 496.485 1562.015 531.335 ;
        RECT 1562.305 179.605 1562.475 227.715 ;
        RECT 1560.005 65.365 1560.175 110.755 ;
      LAYER mcon ;
        RECT 1562.305 1529.745 1562.475 1529.915 ;
        RECT 1561.845 1248.565 1562.015 1248.735 ;
        RECT 1561.845 724.285 1562.015 724.455 ;
        RECT 1561.845 627.725 1562.015 627.895 ;
        RECT 1561.845 531.165 1562.015 531.335 ;
        RECT 1562.305 227.545 1562.475 227.715 ;
        RECT 1560.005 110.585 1560.175 110.755 ;
      LAYER met1 ;
        RECT 1562.230 1692.080 1562.550 1692.140 ;
        RECT 1564.530 1692.080 1564.850 1692.140 ;
        RECT 1562.230 1691.940 1564.850 1692.080 ;
        RECT 1562.230 1691.880 1562.550 1691.940 ;
        RECT 1564.530 1691.880 1564.850 1691.940 ;
        RECT 1561.770 1594.160 1562.090 1594.220 ;
        RECT 1562.230 1594.160 1562.550 1594.220 ;
        RECT 1561.770 1594.020 1562.550 1594.160 ;
        RECT 1561.770 1593.960 1562.090 1594.020 ;
        RECT 1562.230 1593.960 1562.550 1594.020 ;
        RECT 1562.230 1529.900 1562.550 1529.960 ;
        RECT 1562.035 1529.760 1562.550 1529.900 ;
        RECT 1562.230 1529.700 1562.550 1529.760 ;
        RECT 1562.245 1490.800 1562.535 1490.845 ;
        RECT 1562.690 1490.800 1563.010 1490.860 ;
        RECT 1562.245 1490.660 1563.010 1490.800 ;
        RECT 1562.245 1490.615 1562.535 1490.660 ;
        RECT 1562.690 1490.600 1563.010 1490.660 ;
        RECT 1561.770 1442.180 1562.090 1442.240 ;
        RECT 1562.690 1442.180 1563.010 1442.240 ;
        RECT 1561.770 1442.040 1563.010 1442.180 ;
        RECT 1561.770 1441.980 1562.090 1442.040 ;
        RECT 1562.690 1441.980 1563.010 1442.040 ;
        RECT 1561.770 1414.440 1562.090 1414.700 ;
        RECT 1561.860 1414.300 1562.000 1414.440 ;
        RECT 1562.230 1414.300 1562.550 1414.360 ;
        RECT 1561.860 1414.160 1562.550 1414.300 ;
        RECT 1562.230 1414.100 1562.550 1414.160 ;
        RECT 1561.770 1248.720 1562.090 1248.780 ;
        RECT 1561.575 1248.580 1562.090 1248.720 ;
        RECT 1561.770 1248.520 1562.090 1248.580 ;
        RECT 1561.770 1200.780 1562.090 1200.840 ;
        RECT 1561.575 1200.640 1562.090 1200.780 ;
        RECT 1561.770 1200.580 1562.090 1200.640 ;
        RECT 1561.310 1124.960 1561.630 1125.020 ;
        RECT 1562.230 1124.960 1562.550 1125.020 ;
        RECT 1561.310 1124.820 1562.550 1124.960 ;
        RECT 1561.310 1124.760 1561.630 1124.820 ;
        RECT 1562.230 1124.760 1562.550 1124.820 ;
        RECT 1561.310 1028.400 1561.630 1028.460 ;
        RECT 1562.230 1028.400 1562.550 1028.460 ;
        RECT 1561.310 1028.260 1562.550 1028.400 ;
        RECT 1561.310 1028.200 1561.630 1028.260 ;
        RECT 1562.230 1028.200 1562.550 1028.260 ;
        RECT 1561.310 931.840 1561.630 931.900 ;
        RECT 1562.230 931.840 1562.550 931.900 ;
        RECT 1561.310 931.700 1562.550 931.840 ;
        RECT 1561.310 931.640 1561.630 931.700 ;
        RECT 1562.230 931.640 1562.550 931.700 ;
        RECT 1560.850 869.620 1561.170 869.680 ;
        RECT 1562.230 869.620 1562.550 869.680 ;
        RECT 1560.850 869.480 1562.550 869.620 ;
        RECT 1560.850 869.420 1561.170 869.480 ;
        RECT 1562.230 869.420 1562.550 869.480 ;
        RECT 1561.310 818.280 1561.630 818.340 ;
        RECT 1562.230 818.280 1562.550 818.340 ;
        RECT 1561.310 818.140 1562.550 818.280 ;
        RECT 1561.310 818.080 1561.630 818.140 ;
        RECT 1562.230 818.080 1562.550 818.140 ;
        RECT 1561.770 724.440 1562.090 724.500 ;
        RECT 1561.575 724.300 1562.090 724.440 ;
        RECT 1561.770 724.240 1562.090 724.300 ;
        RECT 1561.770 689.760 1562.090 689.820 ;
        RECT 1561.575 689.620 1562.090 689.760 ;
        RECT 1561.770 689.560 1562.090 689.620 ;
        RECT 1561.310 641.820 1561.630 641.880 ;
        RECT 1562.230 641.820 1562.550 641.880 ;
        RECT 1561.310 641.680 1562.550 641.820 ;
        RECT 1561.310 641.620 1561.630 641.680 ;
        RECT 1562.230 641.620 1562.550 641.680 ;
        RECT 1561.770 627.880 1562.090 627.940 ;
        RECT 1561.575 627.740 1562.090 627.880 ;
        RECT 1561.770 627.680 1562.090 627.740 ;
        RECT 1561.770 593.200 1562.090 593.260 ;
        RECT 1561.575 593.060 1562.090 593.200 ;
        RECT 1561.770 593.000 1562.090 593.060 ;
        RECT 1561.310 545.260 1561.630 545.320 ;
        RECT 1562.230 545.260 1562.550 545.320 ;
        RECT 1561.310 545.120 1562.550 545.260 ;
        RECT 1561.310 545.060 1561.630 545.120 ;
        RECT 1562.230 545.060 1562.550 545.120 ;
        RECT 1561.770 531.320 1562.090 531.380 ;
        RECT 1561.575 531.180 1562.090 531.320 ;
        RECT 1561.770 531.120 1562.090 531.180 ;
        RECT 1561.770 496.640 1562.090 496.700 ;
        RECT 1561.575 496.500 1562.090 496.640 ;
        RECT 1561.770 496.440 1562.090 496.500 ;
        RECT 1561.310 448.360 1561.630 448.420 ;
        RECT 1562.230 448.360 1562.550 448.420 ;
        RECT 1561.310 448.220 1562.550 448.360 ;
        RECT 1561.310 448.160 1561.630 448.220 ;
        RECT 1562.230 448.160 1562.550 448.220 ;
        RECT 1560.850 338.200 1561.170 338.260 ;
        RECT 1561.310 338.200 1561.630 338.260 ;
        RECT 1560.850 338.060 1561.630 338.200 ;
        RECT 1560.850 338.000 1561.170 338.060 ;
        RECT 1561.310 338.000 1561.630 338.060 ;
        RECT 1560.850 302.840 1561.170 302.900 ;
        RECT 1561.770 302.840 1562.090 302.900 ;
        RECT 1560.850 302.700 1562.090 302.840 ;
        RECT 1560.850 302.640 1561.170 302.700 ;
        RECT 1561.770 302.640 1562.090 302.700 ;
        RECT 1561.770 255.380 1562.090 255.640 ;
        RECT 1561.860 254.900 1562.000 255.380 ;
        RECT 1562.690 254.900 1563.010 254.960 ;
        RECT 1561.860 254.760 1563.010 254.900 ;
        RECT 1562.690 254.700 1563.010 254.760 ;
        RECT 1562.245 227.700 1562.535 227.745 ;
        RECT 1562.690 227.700 1563.010 227.760 ;
        RECT 1562.245 227.560 1563.010 227.700 ;
        RECT 1562.245 227.515 1562.535 227.560 ;
        RECT 1562.690 227.500 1563.010 227.560 ;
        RECT 1562.230 179.760 1562.550 179.820 ;
        RECT 1562.035 179.620 1562.550 179.760 ;
        RECT 1562.230 179.560 1562.550 179.620 ;
        RECT 1559.945 110.740 1560.235 110.785 ;
        RECT 1561.310 110.740 1561.630 110.800 ;
        RECT 1559.945 110.600 1561.630 110.740 ;
        RECT 1559.945 110.555 1560.235 110.600 ;
        RECT 1561.310 110.540 1561.630 110.600 ;
        RECT 1559.945 65.520 1560.235 65.565 ;
        RECT 1561.770 65.520 1562.090 65.580 ;
        RECT 1559.945 65.380 1562.090 65.520 ;
        RECT 1559.945 65.335 1560.235 65.380 ;
        RECT 1561.770 65.320 1562.090 65.380 ;
        RECT 1536.930 16.900 1537.250 16.960 ;
        RECT 1561.770 16.900 1562.090 16.960 ;
        RECT 1536.930 16.760 1562.090 16.900 ;
        RECT 1536.930 16.700 1537.250 16.760 ;
        RECT 1561.770 16.700 1562.090 16.760 ;
      LAYER via ;
        RECT 1562.260 1691.880 1562.520 1692.140 ;
        RECT 1564.560 1691.880 1564.820 1692.140 ;
        RECT 1561.800 1593.960 1562.060 1594.220 ;
        RECT 1562.260 1593.960 1562.520 1594.220 ;
        RECT 1562.260 1529.700 1562.520 1529.960 ;
        RECT 1562.720 1490.600 1562.980 1490.860 ;
        RECT 1561.800 1441.980 1562.060 1442.240 ;
        RECT 1562.720 1441.980 1562.980 1442.240 ;
        RECT 1561.800 1414.440 1562.060 1414.700 ;
        RECT 1562.260 1414.100 1562.520 1414.360 ;
        RECT 1561.800 1248.520 1562.060 1248.780 ;
        RECT 1561.800 1200.580 1562.060 1200.840 ;
        RECT 1561.340 1124.760 1561.600 1125.020 ;
        RECT 1562.260 1124.760 1562.520 1125.020 ;
        RECT 1561.340 1028.200 1561.600 1028.460 ;
        RECT 1562.260 1028.200 1562.520 1028.460 ;
        RECT 1561.340 931.640 1561.600 931.900 ;
        RECT 1562.260 931.640 1562.520 931.900 ;
        RECT 1560.880 869.420 1561.140 869.680 ;
        RECT 1562.260 869.420 1562.520 869.680 ;
        RECT 1561.340 818.080 1561.600 818.340 ;
        RECT 1562.260 818.080 1562.520 818.340 ;
        RECT 1561.800 724.240 1562.060 724.500 ;
        RECT 1561.800 689.560 1562.060 689.820 ;
        RECT 1561.340 641.620 1561.600 641.880 ;
        RECT 1562.260 641.620 1562.520 641.880 ;
        RECT 1561.800 627.680 1562.060 627.940 ;
        RECT 1561.800 593.000 1562.060 593.260 ;
        RECT 1561.340 545.060 1561.600 545.320 ;
        RECT 1562.260 545.060 1562.520 545.320 ;
        RECT 1561.800 531.120 1562.060 531.380 ;
        RECT 1561.800 496.440 1562.060 496.700 ;
        RECT 1561.340 448.160 1561.600 448.420 ;
        RECT 1562.260 448.160 1562.520 448.420 ;
        RECT 1560.880 338.000 1561.140 338.260 ;
        RECT 1561.340 338.000 1561.600 338.260 ;
        RECT 1560.880 302.640 1561.140 302.900 ;
        RECT 1561.800 302.640 1562.060 302.900 ;
        RECT 1561.800 255.380 1562.060 255.640 ;
        RECT 1562.720 254.700 1562.980 254.960 ;
        RECT 1562.720 227.500 1562.980 227.760 ;
        RECT 1562.260 179.560 1562.520 179.820 ;
        RECT 1561.340 110.540 1561.600 110.800 ;
        RECT 1561.800 65.320 1562.060 65.580 ;
        RECT 1536.960 16.700 1537.220 16.960 ;
        RECT 1561.800 16.700 1562.060 16.960 ;
      LAYER met2 ;
        RECT 1564.550 1700.000 1564.830 1704.000 ;
        RECT 1564.620 1692.170 1564.760 1700.000 ;
        RECT 1562.260 1691.850 1562.520 1692.170 ;
        RECT 1564.560 1691.850 1564.820 1692.170 ;
        RECT 1562.320 1594.250 1562.460 1691.850 ;
        RECT 1561.800 1593.930 1562.060 1594.250 ;
        RECT 1562.260 1593.930 1562.520 1594.250 ;
        RECT 1561.860 1559.650 1562.000 1593.930 ;
        RECT 1561.860 1559.510 1562.460 1559.650 ;
        RECT 1562.320 1529.990 1562.460 1559.510 ;
        RECT 1562.260 1529.670 1562.520 1529.990 ;
        RECT 1562.720 1490.570 1562.980 1490.890 ;
        RECT 1562.780 1442.270 1562.920 1490.570 ;
        RECT 1561.800 1441.950 1562.060 1442.270 ;
        RECT 1562.720 1441.950 1562.980 1442.270 ;
        RECT 1561.860 1414.730 1562.000 1441.950 ;
        RECT 1561.800 1414.410 1562.060 1414.730 ;
        RECT 1562.260 1414.070 1562.520 1414.390 ;
        RECT 1562.320 1316.890 1562.460 1414.070 ;
        RECT 1561.400 1316.750 1562.460 1316.890 ;
        RECT 1561.400 1248.890 1561.540 1316.750 ;
        RECT 1561.400 1248.810 1562.000 1248.890 ;
        RECT 1561.400 1248.750 1562.060 1248.810 ;
        RECT 1561.800 1248.490 1562.060 1248.750 ;
        RECT 1561.800 1200.550 1562.060 1200.870 ;
        RECT 1561.860 1173.410 1562.000 1200.550 ;
        RECT 1561.860 1173.270 1562.460 1173.410 ;
        RECT 1562.320 1125.050 1562.460 1173.270 ;
        RECT 1561.340 1124.730 1561.600 1125.050 ;
        RECT 1562.260 1124.730 1562.520 1125.050 ;
        RECT 1561.400 1124.450 1561.540 1124.730 ;
        RECT 1561.400 1124.310 1562.000 1124.450 ;
        RECT 1561.860 1076.850 1562.000 1124.310 ;
        RECT 1561.860 1076.710 1562.460 1076.850 ;
        RECT 1562.320 1028.490 1562.460 1076.710 ;
        RECT 1561.340 1028.170 1561.600 1028.490 ;
        RECT 1562.260 1028.170 1562.520 1028.490 ;
        RECT 1561.400 1027.890 1561.540 1028.170 ;
        RECT 1561.400 1027.750 1562.000 1027.890 ;
        RECT 1561.860 980.290 1562.000 1027.750 ;
        RECT 1561.860 980.150 1562.460 980.290 ;
        RECT 1562.320 931.930 1562.460 980.150 ;
        RECT 1561.340 931.610 1561.600 931.930 ;
        RECT 1562.260 931.610 1562.520 931.930 ;
        RECT 1561.400 931.330 1561.540 931.610 ;
        RECT 1561.400 931.190 1562.000 931.330 ;
        RECT 1561.860 917.845 1562.000 931.190 ;
        RECT 1560.870 917.475 1561.150 917.845 ;
        RECT 1561.790 917.475 1562.070 917.845 ;
        RECT 1560.940 869.710 1561.080 917.475 ;
        RECT 1560.880 869.390 1561.140 869.710 ;
        RECT 1562.260 869.390 1562.520 869.710 ;
        RECT 1562.320 818.370 1562.460 869.390 ;
        RECT 1561.340 818.050 1561.600 818.370 ;
        RECT 1562.260 818.050 1562.520 818.370 ;
        RECT 1561.400 787.170 1561.540 818.050 ;
        RECT 1560.940 787.030 1561.540 787.170 ;
        RECT 1560.940 766.090 1561.080 787.030 ;
        RECT 1560.940 765.950 1561.540 766.090 ;
        RECT 1561.400 738.210 1561.540 765.950 ;
        RECT 1561.400 738.070 1562.000 738.210 ;
        RECT 1561.860 724.530 1562.000 738.070 ;
        RECT 1561.800 724.210 1562.060 724.530 ;
        RECT 1561.800 689.530 1562.060 689.850 ;
        RECT 1561.860 676.330 1562.000 689.530 ;
        RECT 1561.860 676.190 1562.460 676.330 ;
        RECT 1562.320 641.910 1562.460 676.190 ;
        RECT 1561.340 641.650 1561.600 641.910 ;
        RECT 1561.340 641.590 1562.000 641.650 ;
        RECT 1562.260 641.590 1562.520 641.910 ;
        RECT 1561.400 641.510 1562.000 641.590 ;
        RECT 1561.860 627.970 1562.000 641.510 ;
        RECT 1561.800 627.650 1562.060 627.970 ;
        RECT 1561.800 592.970 1562.060 593.290 ;
        RECT 1561.860 579.770 1562.000 592.970 ;
        RECT 1561.860 579.630 1562.460 579.770 ;
        RECT 1562.320 545.350 1562.460 579.630 ;
        RECT 1561.340 545.090 1561.600 545.350 ;
        RECT 1561.340 545.030 1562.000 545.090 ;
        RECT 1562.260 545.030 1562.520 545.350 ;
        RECT 1561.400 544.950 1562.000 545.030 ;
        RECT 1561.860 531.410 1562.000 544.950 ;
        RECT 1561.800 531.090 1562.060 531.410 ;
        RECT 1561.800 496.410 1562.060 496.730 ;
        RECT 1561.860 483.210 1562.000 496.410 ;
        RECT 1561.860 483.070 1562.460 483.210 ;
        RECT 1562.320 448.450 1562.460 483.070 ;
        RECT 1561.340 448.130 1561.600 448.450 ;
        RECT 1562.260 448.130 1562.520 448.450 ;
        RECT 1561.400 400.930 1561.540 448.130 ;
        RECT 1560.940 400.790 1561.540 400.930 ;
        RECT 1560.940 400.250 1561.080 400.790 ;
        RECT 1560.940 400.110 1561.540 400.250 ;
        RECT 1561.400 338.290 1561.540 400.110 ;
        RECT 1560.880 337.970 1561.140 338.290 ;
        RECT 1561.340 337.970 1561.600 338.290 ;
        RECT 1560.940 302.930 1561.080 337.970 ;
        RECT 1560.880 302.610 1561.140 302.930 ;
        RECT 1561.800 302.610 1562.060 302.930 ;
        RECT 1561.860 255.670 1562.000 302.610 ;
        RECT 1561.800 255.350 1562.060 255.670 ;
        RECT 1562.720 254.670 1562.980 254.990 ;
        RECT 1562.780 227.790 1562.920 254.670 ;
        RECT 1562.720 227.470 1562.980 227.790 ;
        RECT 1562.260 179.530 1562.520 179.850 ;
        RECT 1562.320 154.770 1562.460 179.530 ;
        RECT 1561.400 154.630 1562.460 154.770 ;
        RECT 1561.400 110.830 1561.540 154.630 ;
        RECT 1561.340 110.510 1561.600 110.830 ;
        RECT 1561.800 65.290 1562.060 65.610 ;
        RECT 1561.860 16.990 1562.000 65.290 ;
        RECT 1536.960 16.670 1537.220 16.990 ;
        RECT 1561.800 16.670 1562.060 16.990 ;
        RECT 1537.020 2.400 1537.160 16.670 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
      LAYER via2 ;
        RECT 1560.870 917.520 1561.150 917.800 ;
        RECT 1561.790 917.520 1562.070 917.800 ;
      LAYER met3 ;
        RECT 1560.845 917.810 1561.175 917.825 ;
        RECT 1561.765 917.810 1562.095 917.825 ;
        RECT 1560.845 917.510 1562.095 917.810 ;
        RECT 1560.845 917.495 1561.175 917.510 ;
        RECT 1561.765 917.495 1562.095 917.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1559.010 1688.340 1559.330 1688.400 ;
        RECT 1569.590 1688.340 1569.910 1688.400 ;
        RECT 1559.010 1688.200 1569.910 1688.340 ;
        RECT 1559.010 1688.140 1559.330 1688.200 ;
        RECT 1569.590 1688.140 1569.910 1688.200 ;
        RECT 1554.870 15.540 1555.190 15.600 ;
        RECT 1559.010 15.540 1559.330 15.600 ;
        RECT 1554.870 15.400 1559.330 15.540 ;
        RECT 1554.870 15.340 1555.190 15.400 ;
        RECT 1559.010 15.340 1559.330 15.400 ;
      LAYER via ;
        RECT 1559.040 1688.140 1559.300 1688.400 ;
        RECT 1569.620 1688.140 1569.880 1688.400 ;
        RECT 1554.900 15.340 1555.160 15.600 ;
        RECT 1559.040 15.340 1559.300 15.600 ;
      LAYER met2 ;
        RECT 1569.610 1700.000 1569.890 1704.000 ;
        RECT 1569.680 1688.430 1569.820 1700.000 ;
        RECT 1559.040 1688.110 1559.300 1688.430 ;
        RECT 1569.620 1688.110 1569.880 1688.430 ;
        RECT 1559.100 15.630 1559.240 1688.110 ;
        RECT 1554.900 15.310 1555.160 15.630 ;
        RECT 1559.040 15.310 1559.300 15.630 ;
        RECT 1554.960 2.400 1555.100 15.310 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 0.300 ;
=======
      LAYER li1 ;
        RECT 1573.805 1635.485 1573.975 1683.595 ;
        RECT 1573.805 1538.925 1573.975 1587.035 ;
        RECT 1573.805 766.105 1573.975 814.215 ;
        RECT 1573.805 669.545 1573.975 717.655 ;
        RECT 1573.805 572.645 1573.975 620.755 ;
        RECT 1573.805 476.085 1573.975 524.195 ;
        RECT 1573.805 379.525 1573.975 427.635 ;
        RECT 1573.805 282.965 1573.975 331.075 ;
        RECT 1573.345 48.365 1573.515 137.955 ;
      LAYER mcon ;
        RECT 1573.805 1683.425 1573.975 1683.595 ;
        RECT 1573.805 1586.865 1573.975 1587.035 ;
        RECT 1573.805 814.045 1573.975 814.215 ;
        RECT 1573.805 717.485 1573.975 717.655 ;
        RECT 1573.805 620.585 1573.975 620.755 ;
        RECT 1573.805 524.025 1573.975 524.195 ;
        RECT 1573.805 427.465 1573.975 427.635 ;
        RECT 1573.805 330.905 1573.975 331.075 ;
        RECT 1573.345 137.785 1573.515 137.955 ;
      LAYER met1 ;
        RECT 1573.730 1683.580 1574.050 1683.640 ;
        RECT 1573.535 1683.440 1574.050 1683.580 ;
        RECT 1573.730 1683.380 1574.050 1683.440 ;
        RECT 1573.730 1635.640 1574.050 1635.700 ;
        RECT 1573.535 1635.500 1574.050 1635.640 ;
        RECT 1573.730 1635.440 1574.050 1635.500 ;
        RECT 1573.730 1587.020 1574.050 1587.080 ;
        RECT 1573.535 1586.880 1574.050 1587.020 ;
        RECT 1573.730 1586.820 1574.050 1586.880 ;
        RECT 1573.730 1539.080 1574.050 1539.140 ;
        RECT 1573.535 1538.940 1574.050 1539.080 ;
        RECT 1573.730 1538.880 1574.050 1538.940 ;
        RECT 1572.810 1152.500 1573.130 1152.560 ;
        RECT 1573.730 1152.500 1574.050 1152.560 ;
        RECT 1572.810 1152.360 1574.050 1152.500 ;
        RECT 1572.810 1152.300 1573.130 1152.360 ;
        RECT 1573.730 1152.300 1574.050 1152.360 ;
        RECT 1572.810 1007.320 1573.130 1007.380 ;
        RECT 1573.730 1007.320 1574.050 1007.380 ;
        RECT 1572.810 1007.180 1574.050 1007.320 ;
        RECT 1572.810 1007.120 1573.130 1007.180 ;
        RECT 1573.730 1007.120 1574.050 1007.180 ;
        RECT 1572.810 910.760 1573.130 910.820 ;
        RECT 1573.730 910.760 1574.050 910.820 ;
        RECT 1572.810 910.620 1574.050 910.760 ;
        RECT 1572.810 910.560 1573.130 910.620 ;
        RECT 1573.730 910.560 1574.050 910.620 ;
        RECT 1573.730 814.200 1574.050 814.260 ;
        RECT 1573.535 814.060 1574.050 814.200 ;
        RECT 1573.730 814.000 1574.050 814.060 ;
        RECT 1573.730 766.260 1574.050 766.320 ;
        RECT 1573.535 766.120 1574.050 766.260 ;
        RECT 1573.730 766.060 1574.050 766.120 ;
        RECT 1573.730 717.640 1574.050 717.700 ;
        RECT 1573.535 717.500 1574.050 717.640 ;
        RECT 1573.730 717.440 1574.050 717.500 ;
        RECT 1573.730 669.700 1574.050 669.760 ;
        RECT 1573.535 669.560 1574.050 669.700 ;
        RECT 1573.730 669.500 1574.050 669.560 ;
        RECT 1573.730 620.740 1574.050 620.800 ;
        RECT 1573.535 620.600 1574.050 620.740 ;
        RECT 1573.730 620.540 1574.050 620.600 ;
        RECT 1573.730 572.800 1574.050 572.860 ;
        RECT 1573.535 572.660 1574.050 572.800 ;
        RECT 1573.730 572.600 1574.050 572.660 ;
        RECT 1573.730 524.180 1574.050 524.240 ;
        RECT 1573.535 524.040 1574.050 524.180 ;
        RECT 1573.730 523.980 1574.050 524.040 ;
        RECT 1573.730 476.240 1574.050 476.300 ;
        RECT 1573.535 476.100 1574.050 476.240 ;
        RECT 1573.730 476.040 1574.050 476.100 ;
        RECT 1573.730 427.620 1574.050 427.680 ;
        RECT 1573.535 427.480 1574.050 427.620 ;
        RECT 1573.730 427.420 1574.050 427.480 ;
        RECT 1573.730 379.680 1574.050 379.740 ;
        RECT 1573.535 379.540 1574.050 379.680 ;
        RECT 1573.730 379.480 1574.050 379.540 ;
        RECT 1573.730 338.680 1574.050 338.940 ;
        RECT 1573.820 338.260 1573.960 338.680 ;
        RECT 1573.730 338.000 1574.050 338.260 ;
        RECT 1573.730 331.060 1574.050 331.120 ;
        RECT 1573.535 330.920 1574.050 331.060 ;
        RECT 1573.730 330.860 1574.050 330.920 ;
        RECT 1573.730 283.120 1574.050 283.180 ;
        RECT 1573.535 282.980 1574.050 283.120 ;
        RECT 1573.730 282.920 1574.050 282.980 ;
        RECT 1573.285 137.940 1573.575 137.985 ;
        RECT 1573.730 137.940 1574.050 138.000 ;
        RECT 1573.285 137.800 1574.050 137.940 ;
        RECT 1573.285 137.755 1573.575 137.800 ;
        RECT 1573.730 137.740 1574.050 137.800 ;
        RECT 1573.270 48.520 1573.590 48.580 ;
        RECT 1573.075 48.380 1573.590 48.520 ;
        RECT 1573.270 48.320 1573.590 48.380 ;
      LAYER via ;
        RECT 1573.760 1683.380 1574.020 1683.640 ;
        RECT 1573.760 1635.440 1574.020 1635.700 ;
        RECT 1573.760 1586.820 1574.020 1587.080 ;
        RECT 1573.760 1538.880 1574.020 1539.140 ;
        RECT 1572.840 1152.300 1573.100 1152.560 ;
        RECT 1573.760 1152.300 1574.020 1152.560 ;
        RECT 1572.840 1007.120 1573.100 1007.380 ;
        RECT 1573.760 1007.120 1574.020 1007.380 ;
        RECT 1572.840 910.560 1573.100 910.820 ;
        RECT 1573.760 910.560 1574.020 910.820 ;
        RECT 1573.760 814.000 1574.020 814.260 ;
        RECT 1573.760 766.060 1574.020 766.320 ;
        RECT 1573.760 717.440 1574.020 717.700 ;
        RECT 1573.760 669.500 1574.020 669.760 ;
        RECT 1573.760 620.540 1574.020 620.800 ;
        RECT 1573.760 572.600 1574.020 572.860 ;
        RECT 1573.760 523.980 1574.020 524.240 ;
        RECT 1573.760 476.040 1574.020 476.300 ;
        RECT 1573.760 427.420 1574.020 427.680 ;
        RECT 1573.760 379.480 1574.020 379.740 ;
        RECT 1573.760 338.680 1574.020 338.940 ;
        RECT 1573.760 338.000 1574.020 338.260 ;
        RECT 1573.760 330.860 1574.020 331.120 ;
        RECT 1573.760 282.920 1574.020 283.180 ;
        RECT 1573.760 137.740 1574.020 138.000 ;
        RECT 1573.300 48.320 1573.560 48.580 ;
      LAYER met2 ;
        RECT 1574.210 1700.410 1574.490 1704.000 ;
        RECT 1573.820 1700.270 1574.490 1700.410 ;
        RECT 1573.820 1683.670 1573.960 1700.270 ;
        RECT 1574.210 1700.000 1574.490 1700.270 ;
        RECT 1573.760 1683.350 1574.020 1683.670 ;
        RECT 1573.760 1635.410 1574.020 1635.730 ;
        RECT 1573.820 1587.110 1573.960 1635.410 ;
        RECT 1573.760 1586.790 1574.020 1587.110 ;
        RECT 1573.760 1538.850 1574.020 1539.170 ;
        RECT 1573.820 1200.725 1573.960 1538.850 ;
        RECT 1572.830 1200.355 1573.110 1200.725 ;
        RECT 1573.750 1200.355 1574.030 1200.725 ;
        RECT 1572.900 1152.590 1573.040 1200.355 ;
        RECT 1572.840 1152.270 1573.100 1152.590 ;
        RECT 1573.760 1152.270 1574.020 1152.590 ;
        RECT 1573.820 1104.165 1573.960 1152.270 ;
        RECT 1572.830 1103.795 1573.110 1104.165 ;
        RECT 1573.750 1103.795 1574.030 1104.165 ;
        RECT 1572.900 1055.885 1573.040 1103.795 ;
        RECT 1572.830 1055.515 1573.110 1055.885 ;
        RECT 1573.750 1055.515 1574.030 1055.885 ;
        RECT 1573.820 1007.410 1573.960 1055.515 ;
        RECT 1572.840 1007.090 1573.100 1007.410 ;
        RECT 1573.760 1007.090 1574.020 1007.410 ;
        RECT 1572.900 959.325 1573.040 1007.090 ;
        RECT 1572.830 958.955 1573.110 959.325 ;
        RECT 1573.750 958.955 1574.030 959.325 ;
        RECT 1573.820 910.850 1573.960 958.955 ;
        RECT 1572.840 910.530 1573.100 910.850 ;
        RECT 1573.760 910.530 1574.020 910.850 ;
        RECT 1572.900 862.765 1573.040 910.530 ;
        RECT 1572.830 862.395 1573.110 862.765 ;
        RECT 1573.750 862.395 1574.030 862.765 ;
        RECT 1573.820 814.290 1573.960 862.395 ;
        RECT 1573.760 813.970 1574.020 814.290 ;
        RECT 1573.760 766.030 1574.020 766.350 ;
        RECT 1573.820 717.730 1573.960 766.030 ;
        RECT 1573.760 717.410 1574.020 717.730 ;
        RECT 1573.760 669.470 1574.020 669.790 ;
        RECT 1573.820 620.830 1573.960 669.470 ;
        RECT 1573.760 620.510 1574.020 620.830 ;
        RECT 1573.760 572.570 1574.020 572.890 ;
        RECT 1573.820 524.270 1573.960 572.570 ;
        RECT 1573.760 523.950 1574.020 524.270 ;
        RECT 1573.760 476.010 1574.020 476.330 ;
        RECT 1573.820 427.710 1573.960 476.010 ;
        RECT 1573.760 427.390 1574.020 427.710 ;
        RECT 1573.760 379.450 1574.020 379.770 ;
        RECT 1573.820 338.970 1573.960 379.450 ;
        RECT 1573.760 338.650 1574.020 338.970 ;
        RECT 1573.760 337.970 1574.020 338.290 ;
        RECT 1573.820 331.150 1573.960 337.970 ;
        RECT 1573.760 330.830 1574.020 331.150 ;
        RECT 1573.760 282.890 1574.020 283.210 ;
        RECT 1573.820 138.030 1573.960 282.890 ;
        RECT 1573.760 137.710 1574.020 138.030 ;
        RECT 1573.300 48.290 1573.560 48.610 ;
        RECT 1573.360 14.010 1573.500 48.290 ;
        RECT 1572.900 13.870 1573.500 14.010 ;
        RECT 1572.900 2.400 1573.040 13.870 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
      LAYER via2 ;
        RECT 1572.830 1200.400 1573.110 1200.680 ;
        RECT 1573.750 1200.400 1574.030 1200.680 ;
        RECT 1572.830 1103.840 1573.110 1104.120 ;
        RECT 1573.750 1103.840 1574.030 1104.120 ;
        RECT 1572.830 1055.560 1573.110 1055.840 ;
        RECT 1573.750 1055.560 1574.030 1055.840 ;
        RECT 1572.830 959.000 1573.110 959.280 ;
        RECT 1573.750 959.000 1574.030 959.280 ;
        RECT 1572.830 862.440 1573.110 862.720 ;
        RECT 1573.750 862.440 1574.030 862.720 ;
      LAYER met3 ;
        RECT 1572.805 1200.690 1573.135 1200.705 ;
        RECT 1573.725 1200.690 1574.055 1200.705 ;
        RECT 1572.805 1200.390 1574.055 1200.690 ;
        RECT 1572.805 1200.375 1573.135 1200.390 ;
        RECT 1573.725 1200.375 1574.055 1200.390 ;
        RECT 1572.805 1104.130 1573.135 1104.145 ;
        RECT 1573.725 1104.130 1574.055 1104.145 ;
        RECT 1572.805 1103.830 1574.055 1104.130 ;
        RECT 1572.805 1103.815 1573.135 1103.830 ;
        RECT 1573.725 1103.815 1574.055 1103.830 ;
        RECT 1572.805 1055.850 1573.135 1055.865 ;
        RECT 1573.725 1055.850 1574.055 1055.865 ;
        RECT 1572.805 1055.550 1574.055 1055.850 ;
        RECT 1572.805 1055.535 1573.135 1055.550 ;
        RECT 1573.725 1055.535 1574.055 1055.550 ;
        RECT 1572.805 959.290 1573.135 959.305 ;
        RECT 1573.725 959.290 1574.055 959.305 ;
        RECT 1572.805 958.990 1574.055 959.290 ;
        RECT 1572.805 958.975 1573.135 958.990 ;
        RECT 1573.725 958.975 1574.055 958.990 ;
        RECT 1572.805 862.730 1573.135 862.745 ;
        RECT 1573.725 862.730 1574.055 862.745 ;
        RECT 1572.805 862.430 1574.055 862.730 ;
        RECT 1572.805 862.415 1573.135 862.430 ;
        RECT 1573.725 862.415 1574.055 862.430 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1579.710 20.640 1580.030 20.700 ;
        RECT 1590.290 20.640 1590.610 20.700 ;
        RECT 1579.710 20.500 1590.610 20.640 ;
        RECT 1579.710 20.440 1580.030 20.500 ;
        RECT 1590.290 20.440 1590.610 20.500 ;
      LAYER via ;
        RECT 1579.740 20.440 1580.000 20.700 ;
        RECT 1590.320 20.440 1590.580 20.700 ;
      LAYER met2 ;
        RECT 1579.270 1700.410 1579.550 1704.000 ;
        RECT 1579.270 1700.270 1579.940 1700.410 ;
        RECT 1579.270 1700.000 1579.550 1700.270 ;
        RECT 1579.800 20.730 1579.940 1700.270 ;
        RECT 1579.740 20.410 1580.000 20.730 ;
        RECT 1590.320 20.410 1590.580 20.730 ;
        RECT 1590.380 2.400 1590.520 20.410 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1583.850 1684.260 1584.170 1684.320 ;
        RECT 1585.690 1684.260 1586.010 1684.320 ;
        RECT 1583.850 1684.120 1586.010 1684.260 ;
        RECT 1583.850 1684.060 1584.170 1684.120 ;
        RECT 1585.690 1684.060 1586.010 1684.120 ;
        RECT 1585.690 17.240 1586.010 17.300 ;
        RECT 1608.230 17.240 1608.550 17.300 ;
        RECT 1585.690 17.100 1608.550 17.240 ;
        RECT 1585.690 17.040 1586.010 17.100 ;
        RECT 1608.230 17.040 1608.550 17.100 ;
      LAYER via ;
        RECT 1583.880 1684.060 1584.140 1684.320 ;
        RECT 1585.720 1684.060 1585.980 1684.320 ;
        RECT 1585.720 17.040 1585.980 17.300 ;
        RECT 1608.260 17.040 1608.520 17.300 ;
      LAYER met2 ;
        RECT 1583.870 1700.000 1584.150 1704.000 ;
        RECT 1583.940 1684.350 1584.080 1700.000 ;
        RECT 1583.880 1684.030 1584.140 1684.350 ;
        RECT 1585.720 1684.030 1585.980 1684.350 ;
        RECT 1585.780 17.330 1585.920 1684.030 ;
        RECT 1585.720 17.010 1585.980 17.330 ;
        RECT 1608.260 17.010 1608.520 17.330 ;
        RECT 1608.320 2.400 1608.460 17.010 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1588.910 1683.920 1589.230 1683.980 ;
        RECT 1593.510 1683.920 1593.830 1683.980 ;
        RECT 1588.910 1683.780 1593.830 1683.920 ;
        RECT 1588.910 1683.720 1589.230 1683.780 ;
        RECT 1593.510 1683.720 1593.830 1683.780 ;
        RECT 1593.510 14.520 1593.830 14.580 ;
        RECT 1626.170 14.520 1626.490 14.580 ;
        RECT 1593.510 14.380 1626.490 14.520 ;
        RECT 1593.510 14.320 1593.830 14.380 ;
        RECT 1626.170 14.320 1626.490 14.380 ;
      LAYER via ;
        RECT 1588.940 1683.720 1589.200 1683.980 ;
        RECT 1593.540 1683.720 1593.800 1683.980 ;
        RECT 1593.540 14.320 1593.800 14.580 ;
        RECT 1626.200 14.320 1626.460 14.580 ;
      LAYER met2 ;
        RECT 1588.930 1700.000 1589.210 1704.000 ;
        RECT 1589.000 1684.010 1589.140 1700.000 ;
        RECT 1588.940 1683.690 1589.200 1684.010 ;
        RECT 1593.540 1683.690 1593.800 1684.010 ;
        RECT 1593.600 14.610 1593.740 1683.690 ;
        RECT 1593.540 14.290 1593.800 14.610 ;
        RECT 1626.200 14.290 1626.460 14.610 ;
        RECT 1626.260 2.400 1626.400 14.290 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1593.510 1689.700 1593.830 1689.760 ;
        RECT 1610.990 1689.700 1611.310 1689.760 ;
        RECT 1593.510 1689.560 1611.310 1689.700 ;
        RECT 1593.510 1689.500 1593.830 1689.560 ;
        RECT 1610.990 1689.500 1611.310 1689.560 ;
        RECT 1610.990 17.580 1611.310 17.640 ;
        RECT 1644.110 17.580 1644.430 17.640 ;
        RECT 1610.990 17.440 1644.430 17.580 ;
        RECT 1610.990 17.380 1611.310 17.440 ;
        RECT 1644.110 17.380 1644.430 17.440 ;
      LAYER via ;
        RECT 1593.540 1689.500 1593.800 1689.760 ;
        RECT 1611.020 1689.500 1611.280 1689.760 ;
        RECT 1611.020 17.380 1611.280 17.640 ;
        RECT 1644.140 17.380 1644.400 17.640 ;
      LAYER met2 ;
        RECT 1593.530 1700.000 1593.810 1704.000 ;
        RECT 1593.600 1689.790 1593.740 1700.000 ;
        RECT 1593.540 1689.470 1593.800 1689.790 ;
        RECT 1611.020 1689.470 1611.280 1689.790 ;
        RECT 1611.080 17.670 1611.220 1689.470 ;
        RECT 1611.020 17.350 1611.280 17.670 ;
        RECT 1644.140 17.350 1644.400 17.670 ;
        RECT 1644.200 2.400 1644.340 17.350 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1599.490 19.280 1599.810 19.340 ;
        RECT 1662.050 19.280 1662.370 19.340 ;
        RECT 1599.490 19.140 1662.370 19.280 ;
        RECT 1599.490 19.080 1599.810 19.140 ;
        RECT 1662.050 19.080 1662.370 19.140 ;
      LAYER via ;
        RECT 1599.520 19.080 1599.780 19.340 ;
        RECT 1662.080 19.080 1662.340 19.340 ;
      LAYER met2 ;
        RECT 1598.590 1700.410 1598.870 1704.000 ;
        RECT 1598.590 1700.270 1599.720 1700.410 ;
        RECT 1598.590 1700.000 1598.870 1700.270 ;
        RECT 1599.580 19.370 1599.720 1700.270 ;
        RECT 1599.520 19.050 1599.780 19.370 ;
        RECT 1662.080 19.050 1662.340 19.370 ;
        RECT 1662.140 2.400 1662.280 19.050 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 0.300 ;
=======
      LAYER met1 ;
        RECT 1603.170 1687.660 1603.490 1687.720 ;
        RECT 1673.090 1687.660 1673.410 1687.720 ;
        RECT 1603.170 1687.520 1673.410 1687.660 ;
        RECT 1603.170 1687.460 1603.490 1687.520 ;
        RECT 1673.090 1687.460 1673.410 1687.520 ;
        RECT 1673.090 20.640 1673.410 20.700 ;
        RECT 1679.530 20.640 1679.850 20.700 ;
        RECT 1673.090 20.500 1679.850 20.640 ;
        RECT 1673.090 20.440 1673.410 20.500 ;
        RECT 1679.530 20.440 1679.850 20.500 ;
      LAYER via ;
        RECT 1603.200 1687.460 1603.460 1687.720 ;
        RECT 1673.120 1687.460 1673.380 1687.720 ;
        RECT 1673.120 20.440 1673.380 20.700 ;
        RECT 1679.560 20.440 1679.820 20.700 ;
      LAYER met2 ;
        RECT 1603.190 1700.000 1603.470 1704.000 ;
        RECT 1603.260 1687.750 1603.400 1700.000 ;
        RECT 1603.200 1687.430 1603.460 1687.750 ;
        RECT 1673.120 1687.430 1673.380 1687.750 ;
        RECT 1673.180 20.730 1673.320 1687.430 ;
        RECT 1673.120 20.410 1673.380 20.730 ;
        RECT 1679.560 20.410 1679.820 20.730 ;
        RECT 1679.620 2.400 1679.760 20.410 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1693.790 1687.660 1694.110 1687.720 ;
        RECT 1680.080 1687.520 1694.110 1687.660 ;
        RECT 1608.230 1687.320 1608.550 1687.380 ;
        RECT 1680.080 1687.320 1680.220 1687.520 ;
        RECT 1693.790 1687.460 1694.110 1687.520 ;
        RECT 1608.230 1687.180 1680.220 1687.320 ;
        RECT 1608.230 1687.120 1608.550 1687.180 ;
        RECT 1693.790 17.580 1694.110 17.640 ;
        RECT 1697.470 17.580 1697.790 17.640 ;
        RECT 1693.790 17.440 1697.790 17.580 ;
        RECT 1693.790 17.380 1694.110 17.440 ;
        RECT 1697.470 17.380 1697.790 17.440 ;
      LAYER via ;
        RECT 1608.260 1687.120 1608.520 1687.380 ;
        RECT 1693.820 1687.460 1694.080 1687.720 ;
        RECT 1693.820 17.380 1694.080 17.640 ;
        RECT 1697.500 17.380 1697.760 17.640 ;
      LAYER met2 ;
        RECT 1608.250 1700.000 1608.530 1704.000 ;
        RECT 1608.320 1687.410 1608.460 1700.000 ;
        RECT 1693.820 1687.430 1694.080 1687.750 ;
        RECT 1608.260 1687.090 1608.520 1687.410 ;
        RECT 1693.880 17.670 1694.020 1687.430 ;
        RECT 1693.820 17.350 1694.080 17.670 ;
        RECT 1697.500 17.350 1697.760 17.670 ;
        RECT 1697.560 2.400 1697.700 17.350 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 0.300 ;
=======
      LAYER met1 ;
        RECT 734.230 47.500 734.550 47.560 ;
        RECT 1346.950 47.500 1347.270 47.560 ;
        RECT 734.230 47.360 1347.270 47.500 ;
        RECT 734.230 47.300 734.550 47.360 ;
        RECT 1346.950 47.300 1347.270 47.360 ;
      LAYER via ;
        RECT 734.260 47.300 734.520 47.560 ;
        RECT 1346.980 47.300 1347.240 47.560 ;
      LAYER met2 ;
        RECT 1347.890 1700.410 1348.170 1704.000 ;
        RECT 1347.040 1700.270 1348.170 1700.410 ;
        RECT 1347.040 47.590 1347.180 1700.270 ;
        RECT 1347.890 1700.000 1348.170 1700.270 ;
        RECT 734.260 47.270 734.520 47.590 ;
        RECT 1346.980 47.270 1347.240 47.590 ;
        RECT 734.320 2.400 734.460 47.270 ;
        RECT 734.110 -4.800 734.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 0.300 ;
=======
      LAYER li1 ;
        RECT 1652.925 15.385 1653.095 16.575 ;
      LAYER mcon ;
        RECT 1652.925 16.405 1653.095 16.575 ;
      LAYER met1 ;
        RECT 1613.290 16.900 1613.610 16.960 ;
        RECT 1613.290 16.760 1620.880 16.900 ;
        RECT 1613.290 16.700 1613.610 16.760 ;
        RECT 1620.740 16.560 1620.880 16.760 ;
        RECT 1652.865 16.560 1653.155 16.605 ;
        RECT 1620.740 16.420 1653.155 16.560 ;
        RECT 1652.865 16.375 1653.155 16.420 ;
        RECT 1652.865 15.540 1653.155 15.585 ;
        RECT 1715.410 15.540 1715.730 15.600 ;
        RECT 1652.865 15.400 1715.730 15.540 ;
        RECT 1652.865 15.355 1653.155 15.400 ;
        RECT 1715.410 15.340 1715.730 15.400 ;
      LAYER via ;
        RECT 1613.320 16.700 1613.580 16.960 ;
        RECT 1715.440 15.340 1715.700 15.600 ;
      LAYER met2 ;
        RECT 1612.850 1700.410 1613.130 1704.000 ;
        RECT 1612.850 1700.270 1613.520 1700.410 ;
        RECT 1612.850 1700.000 1613.130 1700.270 ;
        RECT 1613.380 16.990 1613.520 1700.270 ;
        RECT 1613.320 16.670 1613.580 16.990 ;
        RECT 1715.440 15.310 1715.700 15.630 ;
        RECT 1715.500 2.400 1715.640 15.310 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 0.300 ;
=======
      LAYER met1 ;
        RECT 1617.890 1688.680 1618.210 1688.740 ;
        RECT 1620.190 1688.680 1620.510 1688.740 ;
        RECT 1617.890 1688.540 1620.510 1688.680 ;
        RECT 1617.890 1688.480 1618.210 1688.540 ;
        RECT 1620.190 1688.480 1620.510 1688.540 ;
        RECT 1619.730 14.860 1620.050 14.920 ;
        RECT 1733.350 14.860 1733.670 14.920 ;
        RECT 1619.730 14.720 1733.670 14.860 ;
        RECT 1619.730 14.660 1620.050 14.720 ;
        RECT 1733.350 14.660 1733.670 14.720 ;
      LAYER via ;
        RECT 1617.920 1688.480 1618.180 1688.740 ;
        RECT 1620.220 1688.480 1620.480 1688.740 ;
        RECT 1619.760 14.660 1620.020 14.920 ;
        RECT 1733.380 14.660 1733.640 14.920 ;
      LAYER met2 ;
        RECT 1617.910 1700.000 1618.190 1704.000 ;
        RECT 1617.980 1688.770 1618.120 1700.000 ;
        RECT 1617.920 1688.450 1618.180 1688.770 ;
        RECT 1620.220 1688.450 1620.480 1688.770 ;
        RECT 1620.280 20.130 1620.420 1688.450 ;
        RECT 1619.820 19.990 1620.420 20.130 ;
        RECT 1619.820 14.950 1619.960 19.990 ;
        RECT 1619.760 14.630 1620.020 14.950 ;
        RECT 1733.380 14.630 1733.640 14.950 ;
        RECT 1733.440 2.400 1733.580 14.630 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1622.490 1688.340 1622.810 1688.400 ;
        RECT 1627.550 1688.340 1627.870 1688.400 ;
        RECT 1622.490 1688.200 1627.870 1688.340 ;
        RECT 1622.490 1688.140 1622.810 1688.200 ;
        RECT 1627.550 1688.140 1627.870 1688.200 ;
        RECT 1627.550 18.260 1627.870 18.320 ;
        RECT 1751.290 18.260 1751.610 18.320 ;
        RECT 1627.550 18.120 1751.610 18.260 ;
        RECT 1627.550 18.060 1627.870 18.120 ;
        RECT 1751.290 18.060 1751.610 18.120 ;
      LAYER via ;
        RECT 1622.520 1688.140 1622.780 1688.400 ;
        RECT 1627.580 1688.140 1627.840 1688.400 ;
        RECT 1627.580 18.060 1627.840 18.320 ;
        RECT 1751.320 18.060 1751.580 18.320 ;
      LAYER met2 ;
        RECT 1622.510 1700.000 1622.790 1704.000 ;
        RECT 1622.580 1688.430 1622.720 1700.000 ;
        RECT 1622.520 1688.110 1622.780 1688.430 ;
        RECT 1627.580 1688.110 1627.840 1688.430 ;
        RECT 1627.640 18.350 1627.780 1688.110 ;
        RECT 1627.580 18.030 1627.840 18.350 ;
        RECT 1751.320 18.030 1751.580 18.350 ;
        RECT 1751.380 2.400 1751.520 18.030 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 0.300 ;
=======
      LAYER met1 ;
        RECT 1627.090 15.880 1627.410 15.940 ;
        RECT 1768.770 15.880 1769.090 15.940 ;
        RECT 1627.090 15.740 1769.090 15.880 ;
        RECT 1627.090 15.680 1627.410 15.740 ;
        RECT 1768.770 15.680 1769.090 15.740 ;
      LAYER via ;
        RECT 1627.120 15.680 1627.380 15.940 ;
        RECT 1768.800 15.680 1769.060 15.940 ;
      LAYER met2 ;
        RECT 1627.570 1700.410 1627.850 1704.000 ;
        RECT 1627.180 1700.270 1627.850 1700.410 ;
        RECT 1627.180 15.970 1627.320 1700.270 ;
        RECT 1627.570 1700.000 1627.850 1700.270 ;
        RECT 1627.120 15.650 1627.380 15.970 ;
        RECT 1768.800 15.650 1769.060 15.970 ;
        RECT 1768.860 2.400 1769.000 15.650 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 0.300 ;
=======
      LAYER li1 ;
        RECT 1675.005 14.365 1675.175 19.975 ;
      LAYER mcon ;
        RECT 1675.005 19.805 1675.175 19.975 ;
      LAYER met1 ;
        RECT 1632.150 1688.680 1632.470 1688.740 ;
        RECT 1634.450 1688.680 1634.770 1688.740 ;
        RECT 1632.150 1688.540 1634.770 1688.680 ;
        RECT 1632.150 1688.480 1632.470 1688.540 ;
        RECT 1634.450 1688.480 1634.770 1688.540 ;
        RECT 1674.945 19.960 1675.235 20.005 ;
        RECT 1786.710 19.960 1787.030 20.020 ;
        RECT 1674.945 19.820 1787.030 19.960 ;
        RECT 1674.945 19.775 1675.235 19.820 ;
        RECT 1786.710 19.760 1787.030 19.820 ;
        RECT 1634.450 14.520 1634.770 14.580 ;
        RECT 1674.945 14.520 1675.235 14.565 ;
        RECT 1634.450 14.380 1675.235 14.520 ;
        RECT 1634.450 14.320 1634.770 14.380 ;
        RECT 1674.945 14.335 1675.235 14.380 ;
      LAYER via ;
        RECT 1632.180 1688.480 1632.440 1688.740 ;
        RECT 1634.480 1688.480 1634.740 1688.740 ;
        RECT 1786.740 19.760 1787.000 20.020 ;
        RECT 1634.480 14.320 1634.740 14.580 ;
      LAYER met2 ;
        RECT 1632.170 1700.000 1632.450 1704.000 ;
        RECT 1632.240 1688.770 1632.380 1700.000 ;
        RECT 1632.180 1688.450 1632.440 1688.770 ;
        RECT 1634.480 1688.450 1634.740 1688.770 ;
        RECT 1634.540 14.610 1634.680 1688.450 ;
        RECT 1786.740 19.730 1787.000 20.050 ;
        RECT 1634.480 14.290 1634.740 14.610 ;
        RECT 1786.800 2.400 1786.940 19.730 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 0.300 ;
=======
      LAYER li1 ;
        RECT 1641.425 1256.045 1641.595 1257.575 ;
        RECT 1662.585 16.065 1662.755 19.295 ;
      LAYER mcon ;
        RECT 1641.425 1257.405 1641.595 1257.575 ;
        RECT 1662.585 19.125 1662.755 19.295 ;
      LAYER met1 ;
        RECT 1637.210 1688.340 1637.530 1688.400 ;
        RECT 1641.350 1688.340 1641.670 1688.400 ;
        RECT 1637.210 1688.200 1641.670 1688.340 ;
        RECT 1637.210 1688.140 1637.530 1688.200 ;
        RECT 1641.350 1688.140 1641.670 1688.200 ;
        RECT 1641.350 1257.560 1641.670 1257.620 ;
        RECT 1641.155 1257.420 1641.670 1257.560 ;
        RECT 1641.350 1257.360 1641.670 1257.420 ;
        RECT 1641.350 1256.200 1641.670 1256.260 ;
        RECT 1641.155 1256.060 1641.670 1256.200 ;
        RECT 1641.350 1256.000 1641.670 1256.060 ;
        RECT 1641.350 435.920 1641.670 436.180 ;
        RECT 1641.440 435.160 1641.580 435.920 ;
        RECT 1641.350 434.900 1641.670 435.160 ;
        RECT 1641.350 146.240 1641.670 146.500 ;
        RECT 1641.440 145.140 1641.580 146.240 ;
        RECT 1641.350 144.880 1641.670 145.140 ;
        RECT 1662.525 19.280 1662.815 19.325 ;
        RECT 1804.650 19.280 1804.970 19.340 ;
        RECT 1662.525 19.140 1804.970 19.280 ;
        RECT 1662.525 19.095 1662.815 19.140 ;
        RECT 1804.650 19.080 1804.970 19.140 ;
        RECT 1641.350 16.220 1641.670 16.280 ;
        RECT 1662.525 16.220 1662.815 16.265 ;
        RECT 1641.350 16.080 1662.815 16.220 ;
        RECT 1641.350 16.020 1641.670 16.080 ;
        RECT 1662.525 16.035 1662.815 16.080 ;
      LAYER via ;
        RECT 1637.240 1688.140 1637.500 1688.400 ;
        RECT 1641.380 1688.140 1641.640 1688.400 ;
        RECT 1641.380 1257.360 1641.640 1257.620 ;
        RECT 1641.380 1256.000 1641.640 1256.260 ;
        RECT 1641.380 435.920 1641.640 436.180 ;
        RECT 1641.380 434.900 1641.640 435.160 ;
        RECT 1641.380 146.240 1641.640 146.500 ;
        RECT 1641.380 144.880 1641.640 145.140 ;
        RECT 1804.680 19.080 1804.940 19.340 ;
        RECT 1641.380 16.020 1641.640 16.280 ;
      LAYER met2 ;
        RECT 1637.230 1700.000 1637.510 1704.000 ;
        RECT 1637.300 1688.430 1637.440 1700.000 ;
        RECT 1637.240 1688.110 1637.500 1688.430 ;
        RECT 1641.380 1688.110 1641.640 1688.430 ;
        RECT 1641.440 1257.650 1641.580 1688.110 ;
        RECT 1641.380 1257.330 1641.640 1257.650 ;
        RECT 1641.380 1255.970 1641.640 1256.290 ;
        RECT 1641.440 436.210 1641.580 1255.970 ;
        RECT 1641.380 435.890 1641.640 436.210 ;
        RECT 1641.380 434.870 1641.640 435.190 ;
        RECT 1641.440 146.530 1641.580 434.870 ;
        RECT 1641.380 146.210 1641.640 146.530 ;
        RECT 1641.380 144.850 1641.640 145.170 ;
        RECT 1641.440 16.310 1641.580 144.850 ;
        RECT 1804.680 19.050 1804.940 19.370 ;
        RECT 1641.380 15.990 1641.640 16.310 ;
        RECT 1804.740 2.400 1804.880 19.050 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1641.810 1257.020 1642.130 1257.280 ;
        RECT 1641.900 1256.260 1642.040 1257.020 ;
        RECT 1641.810 1256.000 1642.130 1256.260 ;
        RECT 1641.810 145.560 1642.130 145.820 ;
        RECT 1641.900 145.140 1642.040 145.560 ;
        RECT 1641.810 144.880 1642.130 145.140 ;
      LAYER via ;
        RECT 1641.840 1257.020 1642.100 1257.280 ;
        RECT 1641.840 1256.000 1642.100 1256.260 ;
        RECT 1641.840 145.560 1642.100 145.820 ;
        RECT 1641.840 144.880 1642.100 145.140 ;
      LAYER met2 ;
        RECT 1641.830 1700.000 1642.110 1704.000 ;
        RECT 1641.900 1257.310 1642.040 1700.000 ;
        RECT 1641.840 1256.990 1642.100 1257.310 ;
        RECT 1641.840 1255.970 1642.100 1256.290 ;
        RECT 1641.900 145.850 1642.040 1255.970 ;
        RECT 1641.840 145.530 1642.100 145.850 ;
        RECT 1641.840 144.850 1642.100 145.170 ;
        RECT 1641.900 16.845 1642.040 144.850 ;
        RECT 1641.830 16.475 1642.110 16.845 ;
        RECT 1822.610 16.475 1822.890 16.845 ;
        RECT 1822.680 2.400 1822.820 16.475 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
      LAYER via2 ;
        RECT 1641.830 16.520 1642.110 16.800 ;
        RECT 1822.610 16.520 1822.890 16.800 ;
      LAYER met3 ;
        RECT 1641.805 16.810 1642.135 16.825 ;
        RECT 1822.585 16.810 1822.915 16.825 ;
        RECT 1641.805 16.510 1822.915 16.810 ;
        RECT 1641.805 16.495 1642.135 16.510 ;
        RECT 1822.585 16.495 1822.915 16.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 0.300 ;
=======
      LAYER li1 ;
        RECT 1700.765 17.425 1700.935 20.315 ;
        RECT 1820.365 17.425 1820.535 18.955 ;
      LAYER mcon ;
        RECT 1700.765 20.145 1700.935 20.315 ;
        RECT 1820.365 18.785 1820.535 18.955 ;
      LAYER met1 ;
        RECT 1646.870 1685.620 1647.190 1685.680 ;
        RECT 1648.710 1685.620 1649.030 1685.680 ;
        RECT 1646.870 1685.480 1649.030 1685.620 ;
        RECT 1646.870 1685.420 1647.190 1685.480 ;
        RECT 1648.710 1685.420 1649.030 1685.480 ;
        RECT 1700.705 20.300 1700.995 20.345 ;
        RECT 1674.560 20.160 1700.995 20.300 ;
        RECT 1648.710 19.960 1649.030 20.020 ;
        RECT 1674.560 19.960 1674.700 20.160 ;
        RECT 1700.705 20.115 1700.995 20.160 ;
        RECT 1648.710 19.820 1674.700 19.960 ;
        RECT 1648.710 19.760 1649.030 19.820 ;
        RECT 1820.305 18.940 1820.595 18.985 ;
        RECT 1840.070 18.940 1840.390 19.000 ;
        RECT 1820.305 18.800 1840.390 18.940 ;
        RECT 1820.305 18.755 1820.595 18.800 ;
        RECT 1840.070 18.740 1840.390 18.800 ;
        RECT 1700.705 17.580 1700.995 17.625 ;
        RECT 1820.305 17.580 1820.595 17.625 ;
        RECT 1700.705 17.440 1820.595 17.580 ;
        RECT 1700.705 17.395 1700.995 17.440 ;
        RECT 1820.305 17.395 1820.595 17.440 ;
      LAYER via ;
        RECT 1646.900 1685.420 1647.160 1685.680 ;
        RECT 1648.740 1685.420 1649.000 1685.680 ;
        RECT 1648.740 19.760 1649.000 20.020 ;
        RECT 1840.100 18.740 1840.360 19.000 ;
      LAYER met2 ;
        RECT 1646.890 1700.000 1647.170 1704.000 ;
        RECT 1646.960 1685.710 1647.100 1700.000 ;
        RECT 1646.900 1685.390 1647.160 1685.710 ;
        RECT 1648.740 1685.390 1649.000 1685.710 ;
        RECT 1648.800 20.050 1648.940 1685.390 ;
        RECT 1648.740 19.730 1649.000 20.050 ;
        RECT 1840.100 18.710 1840.360 19.030 ;
        RECT 1840.160 2.400 1840.300 18.710 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1651.470 1688.680 1651.790 1688.740 ;
        RECT 1655.610 1688.680 1655.930 1688.740 ;
        RECT 1651.470 1688.540 1655.930 1688.680 ;
        RECT 1651.470 1688.480 1651.790 1688.540 ;
        RECT 1655.610 1688.480 1655.930 1688.540 ;
        RECT 1655.610 17.240 1655.930 17.300 ;
        RECT 1858.010 17.240 1858.330 17.300 ;
        RECT 1655.610 17.100 1858.330 17.240 ;
        RECT 1655.610 17.040 1655.930 17.100 ;
        RECT 1858.010 17.040 1858.330 17.100 ;
      LAYER via ;
        RECT 1651.500 1688.480 1651.760 1688.740 ;
        RECT 1655.640 1688.480 1655.900 1688.740 ;
        RECT 1655.640 17.040 1655.900 17.300 ;
        RECT 1858.040 17.040 1858.300 17.300 ;
      LAYER met2 ;
        RECT 1651.490 1700.000 1651.770 1704.000 ;
        RECT 1651.560 1688.770 1651.700 1700.000 ;
        RECT 1651.500 1688.450 1651.760 1688.770 ;
        RECT 1655.640 1688.450 1655.900 1688.770 ;
        RECT 1655.700 17.330 1655.840 1688.450 ;
        RECT 1655.640 17.010 1655.900 17.330 ;
        RECT 1858.040 17.010 1858.300 17.330 ;
        RECT 1858.100 2.400 1858.240 17.010 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 0.300 ;
=======
      LAYER li1 ;
        RECT 1763.325 14.365 1763.495 15.215 ;
      LAYER mcon ;
        RECT 1763.325 15.045 1763.495 15.215 ;
      LAYER met1 ;
        RECT 1656.070 1686.980 1656.390 1687.040 ;
        RECT 1742.090 1686.980 1742.410 1687.040 ;
        RECT 1656.070 1686.840 1742.410 1686.980 ;
        RECT 1656.070 1686.780 1656.390 1686.840 ;
        RECT 1742.090 1686.780 1742.410 1686.840 ;
        RECT 1763.265 15.200 1763.555 15.245 ;
        RECT 1875.950 15.200 1876.270 15.260 ;
        RECT 1763.265 15.060 1876.270 15.200 ;
        RECT 1763.265 15.015 1763.555 15.060 ;
        RECT 1875.950 15.000 1876.270 15.060 ;
        RECT 1763.265 14.520 1763.555 14.565 ;
        RECT 1745.860 14.380 1763.555 14.520 ;
        RECT 1742.090 14.180 1742.410 14.240 ;
        RECT 1745.860 14.180 1746.000 14.380 ;
        RECT 1763.265 14.335 1763.555 14.380 ;
        RECT 1742.090 14.040 1746.000 14.180 ;
        RECT 1742.090 13.980 1742.410 14.040 ;
      LAYER via ;
        RECT 1656.100 1686.780 1656.360 1687.040 ;
        RECT 1742.120 1686.780 1742.380 1687.040 ;
        RECT 1875.980 15.000 1876.240 15.260 ;
        RECT 1742.120 13.980 1742.380 14.240 ;
      LAYER met2 ;
        RECT 1656.090 1700.000 1656.370 1704.000 ;
        RECT 1656.160 1687.070 1656.300 1700.000 ;
        RECT 1656.100 1686.750 1656.360 1687.070 ;
        RECT 1742.120 1686.750 1742.380 1687.070 ;
        RECT 1742.180 14.270 1742.320 1686.750 ;
        RECT 1875.980 14.970 1876.240 15.290 ;
        RECT 1742.120 13.950 1742.380 14.270 ;
        RECT 1876.040 2.400 1876.180 14.970 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 0.300 ;
=======
      LAYER met1 ;
        RECT 752.170 47.840 752.490 47.900 ;
        RECT 1352.470 47.840 1352.790 47.900 ;
        RECT 752.170 47.700 1352.790 47.840 ;
        RECT 752.170 47.640 752.490 47.700 ;
        RECT 1352.470 47.640 1352.790 47.700 ;
      LAYER via ;
        RECT 752.200 47.640 752.460 47.900 ;
        RECT 1352.500 47.640 1352.760 47.900 ;
      LAYER met2 ;
        RECT 1352.490 1700.000 1352.770 1704.000 ;
        RECT 1352.560 47.930 1352.700 1700.000 ;
        RECT 752.200 47.610 752.460 47.930 ;
        RECT 1352.500 47.610 1352.760 47.930 ;
        RECT 752.260 2.400 752.400 47.610 ;
        RECT 752.050 -4.800 752.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1669.500 1688.200 1677.000 1688.340 ;
        RECT 1661.130 1688.000 1661.450 1688.060 ;
        RECT 1669.500 1688.000 1669.640 1688.200 ;
        RECT 1661.130 1687.860 1669.640 1688.000 ;
        RECT 1676.860 1688.000 1677.000 1688.200 ;
        RECT 1676.860 1687.860 1694.480 1688.000 ;
        RECT 1661.130 1687.800 1661.450 1687.860 ;
        RECT 1694.340 1687.660 1694.480 1687.860 ;
        RECT 1721.390 1687.660 1721.710 1687.720 ;
        RECT 1694.340 1687.520 1721.710 1687.660 ;
        RECT 1721.390 1687.460 1721.710 1687.520 ;
        RECT 1721.390 15.540 1721.710 15.600 ;
        RECT 1893.890 15.540 1894.210 15.600 ;
        RECT 1721.390 15.400 1894.210 15.540 ;
        RECT 1721.390 15.340 1721.710 15.400 ;
        RECT 1893.890 15.340 1894.210 15.400 ;
      LAYER via ;
        RECT 1661.160 1687.800 1661.420 1688.060 ;
        RECT 1721.420 1687.460 1721.680 1687.720 ;
        RECT 1721.420 15.340 1721.680 15.600 ;
        RECT 1893.920 15.340 1894.180 15.600 ;
      LAYER met2 ;
        RECT 1661.150 1700.000 1661.430 1704.000 ;
        RECT 1661.220 1688.090 1661.360 1700.000 ;
        RECT 1661.160 1687.770 1661.420 1688.090 ;
        RECT 1721.420 1687.430 1721.680 1687.750 ;
        RECT 1721.480 15.630 1721.620 1687.430 ;
        RECT 1721.420 15.310 1721.680 15.630 ;
        RECT 1893.920 15.310 1894.180 15.630 ;
        RECT 1893.980 2.400 1894.120 15.310 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1665.730 1689.020 1666.050 1689.080 ;
        RECT 1669.410 1689.020 1669.730 1689.080 ;
        RECT 1665.730 1688.880 1669.730 1689.020 ;
        RECT 1665.730 1688.820 1666.050 1688.880 ;
        RECT 1669.410 1688.820 1669.730 1688.880 ;
        RECT 1669.410 16.220 1669.730 16.280 ;
        RECT 1911.830 16.220 1912.150 16.280 ;
        RECT 1669.410 16.080 1912.150 16.220 ;
        RECT 1669.410 16.020 1669.730 16.080 ;
        RECT 1911.830 16.020 1912.150 16.080 ;
      LAYER via ;
        RECT 1665.760 1688.820 1666.020 1689.080 ;
        RECT 1669.440 1688.820 1669.700 1689.080 ;
        RECT 1669.440 16.020 1669.700 16.280 ;
        RECT 1911.860 16.020 1912.120 16.280 ;
      LAYER met2 ;
        RECT 1665.750 1700.000 1666.030 1704.000 ;
        RECT 1665.820 1689.110 1665.960 1700.000 ;
        RECT 1665.760 1688.790 1666.020 1689.110 ;
        RECT 1669.440 1688.790 1669.700 1689.110 ;
        RECT 1669.500 16.310 1669.640 1688.790 ;
        RECT 1669.440 15.990 1669.700 16.310 ;
        RECT 1911.860 15.990 1912.120 16.310 ;
        RECT 1911.920 2.400 1912.060 15.990 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1670.790 1689.020 1671.110 1689.080 ;
        RECT 1676.310 1689.020 1676.630 1689.080 ;
        RECT 1670.790 1688.880 1676.630 1689.020 ;
        RECT 1670.790 1688.820 1671.110 1688.880 ;
        RECT 1676.310 1688.820 1676.630 1688.880 ;
        RECT 1676.310 16.560 1676.630 16.620 ;
        RECT 1929.310 16.560 1929.630 16.620 ;
        RECT 1676.310 16.420 1929.630 16.560 ;
        RECT 1676.310 16.360 1676.630 16.420 ;
        RECT 1929.310 16.360 1929.630 16.420 ;
      LAYER via ;
        RECT 1670.820 1688.820 1671.080 1689.080 ;
        RECT 1676.340 1688.820 1676.600 1689.080 ;
        RECT 1676.340 16.360 1676.600 16.620 ;
        RECT 1929.340 16.360 1929.600 16.620 ;
      LAYER met2 ;
        RECT 1670.810 1700.000 1671.090 1704.000 ;
        RECT 1670.880 1689.110 1671.020 1700.000 ;
        RECT 1670.820 1688.790 1671.080 1689.110 ;
        RECT 1676.340 1688.790 1676.600 1689.110 ;
        RECT 1676.400 16.650 1676.540 1688.790 ;
        RECT 1676.340 16.330 1676.600 16.650 ;
        RECT 1929.340 16.330 1929.600 16.650 ;
        RECT 1929.400 2.400 1929.540 16.330 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1947.130 -4.800 1947.690 0.300 ;
=======
        RECT 1675.410 1700.410 1675.690 1704.000 ;
        RECT 1675.410 1700.270 1676.080 1700.410 ;
        RECT 1675.410 1700.000 1675.690 1700.270 ;
        RECT 1675.940 15.485 1676.080 1700.270 ;
        RECT 1675.870 15.115 1676.150 15.485 ;
        RECT 1947.270 15.115 1947.550 15.485 ;
        RECT 1947.340 2.400 1947.480 15.115 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
      LAYER via2 ;
        RECT 1675.870 15.160 1676.150 15.440 ;
        RECT 1947.270 15.160 1947.550 15.440 ;
      LAYER met3 ;
        RECT 1675.845 15.450 1676.175 15.465 ;
        RECT 1947.245 15.450 1947.575 15.465 ;
        RECT 1675.845 15.150 1947.575 15.450 ;
        RECT 1675.845 15.135 1676.175 15.150 ;
        RECT 1947.245 15.135 1947.575 15.150 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 0.300 ;
=======
      LAYER li1 ;
        RECT 1689.265 19.635 1689.435 20.655 ;
        RECT 1703.525 20.485 1705.535 20.655 ;
        RECT 1689.265 19.465 1692.195 19.635 ;
        RECT 1703.525 19.465 1703.695 20.485 ;
      LAYER mcon ;
        RECT 1689.265 20.485 1689.435 20.655 ;
        RECT 1705.365 20.485 1705.535 20.655 ;
        RECT 1692.025 19.465 1692.195 19.635 ;
      LAYER met1 ;
        RECT 1680.450 1687.320 1680.770 1687.380 ;
        RECT 1683.210 1687.320 1683.530 1687.380 ;
        RECT 1680.450 1687.180 1683.530 1687.320 ;
        RECT 1680.450 1687.120 1680.770 1687.180 ;
        RECT 1683.210 1687.120 1683.530 1687.180 ;
        RECT 1683.210 20.640 1683.530 20.700 ;
        RECT 1689.205 20.640 1689.495 20.685 ;
        RECT 1683.210 20.500 1689.495 20.640 ;
        RECT 1683.210 20.440 1683.530 20.500 ;
        RECT 1689.205 20.455 1689.495 20.500 ;
        RECT 1705.305 20.640 1705.595 20.685 ;
        RECT 1965.190 20.640 1965.510 20.700 ;
        RECT 1705.305 20.500 1965.510 20.640 ;
        RECT 1705.305 20.455 1705.595 20.500 ;
        RECT 1965.190 20.440 1965.510 20.500 ;
        RECT 1691.965 19.620 1692.255 19.665 ;
        RECT 1703.465 19.620 1703.755 19.665 ;
        RECT 1691.965 19.480 1703.755 19.620 ;
        RECT 1691.965 19.435 1692.255 19.480 ;
        RECT 1703.465 19.435 1703.755 19.480 ;
      LAYER via ;
        RECT 1680.480 1687.120 1680.740 1687.380 ;
        RECT 1683.240 1687.120 1683.500 1687.380 ;
        RECT 1683.240 20.440 1683.500 20.700 ;
        RECT 1965.220 20.440 1965.480 20.700 ;
      LAYER met2 ;
        RECT 1680.470 1700.000 1680.750 1704.000 ;
        RECT 1680.540 1687.410 1680.680 1700.000 ;
        RECT 1680.480 1687.090 1680.740 1687.410 ;
        RECT 1683.240 1687.090 1683.500 1687.410 ;
        RECT 1683.300 20.730 1683.440 1687.090 ;
        RECT 1683.240 20.410 1683.500 20.730 ;
        RECT 1965.220 20.410 1965.480 20.730 ;
        RECT 1965.280 2.400 1965.420 20.410 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1685.050 1684.600 1685.370 1684.660 ;
        RECT 1689.650 1684.600 1689.970 1684.660 ;
        RECT 1685.050 1684.460 1689.970 1684.600 ;
        RECT 1685.050 1684.400 1685.370 1684.460 ;
        RECT 1689.650 1684.400 1689.970 1684.460 ;
        RECT 1689.650 20.640 1689.970 20.700 ;
        RECT 1689.650 20.500 1705.060 20.640 ;
        RECT 1689.650 20.440 1689.970 20.500 ;
        RECT 1704.920 20.300 1705.060 20.500 ;
        RECT 1983.130 20.300 1983.450 20.360 ;
        RECT 1704.920 20.160 1983.450 20.300 ;
        RECT 1983.130 20.100 1983.450 20.160 ;
      LAYER via ;
        RECT 1685.080 1684.400 1685.340 1684.660 ;
        RECT 1689.680 1684.400 1689.940 1684.660 ;
        RECT 1689.680 20.440 1689.940 20.700 ;
        RECT 1983.160 20.100 1983.420 20.360 ;
      LAYER met2 ;
        RECT 1685.070 1700.000 1685.350 1704.000 ;
        RECT 1685.140 1684.690 1685.280 1700.000 ;
        RECT 1685.080 1684.370 1685.340 1684.690 ;
        RECT 1689.680 1684.370 1689.940 1684.690 ;
        RECT 1689.740 20.730 1689.880 1684.370 ;
        RECT 1689.680 20.410 1689.940 20.730 ;
        RECT 1983.160 20.070 1983.420 20.390 ;
        RECT 1983.220 2.400 1983.360 20.070 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2000.950 -4.800 2001.510 0.300 ;
=======
        RECT 1690.130 1700.000 1690.410 1704.000 ;
        RECT 1690.200 16.165 1690.340 1700.000 ;
        RECT 1690.130 15.795 1690.410 16.165 ;
        RECT 2001.090 15.795 2001.370 16.165 ;
        RECT 2001.160 2.400 2001.300 15.795 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
      LAYER via2 ;
        RECT 1690.130 15.840 1690.410 16.120 ;
        RECT 2001.090 15.840 2001.370 16.120 ;
      LAYER met3 ;
        RECT 1690.105 16.130 1690.435 16.145 ;
        RECT 2001.065 16.130 2001.395 16.145 ;
        RECT 1690.105 15.830 2001.395 16.130 ;
        RECT 1690.105 15.815 1690.435 15.830 ;
        RECT 2001.065 15.815 2001.395 15.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1694.710 1685.960 1695.030 1686.020 ;
        RECT 1697.010 1685.960 1697.330 1686.020 ;
        RECT 1694.710 1685.820 1697.330 1685.960 ;
        RECT 1694.710 1685.760 1695.030 1685.820 ;
        RECT 1697.010 1685.760 1697.330 1685.820 ;
      LAYER via ;
        RECT 1694.740 1685.760 1695.000 1686.020 ;
        RECT 1697.040 1685.760 1697.300 1686.020 ;
      LAYER met2 ;
        RECT 1694.730 1700.000 1695.010 1704.000 ;
        RECT 1694.800 1686.050 1694.940 1700.000 ;
        RECT 1694.740 1685.730 1695.000 1686.050 ;
        RECT 1697.040 1685.730 1697.300 1686.050 ;
        RECT 1697.100 20.245 1697.240 1685.730 ;
        RECT 1697.030 19.875 1697.310 20.245 ;
        RECT 2018.570 19.875 2018.850 20.245 ;
        RECT 2018.640 2.400 2018.780 19.875 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
      LAYER via2 ;
        RECT 1697.030 19.920 1697.310 20.200 ;
        RECT 2018.570 19.920 2018.850 20.200 ;
      LAYER met3 ;
        RECT 1697.005 20.210 1697.335 20.225 ;
        RECT 2018.545 20.210 2018.875 20.225 ;
        RECT 1697.005 19.910 2018.875 20.210 ;
        RECT 1697.005 19.895 1697.335 19.910 ;
        RECT 2018.545 19.895 2018.875 19.910 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1699.770 1689.020 1700.090 1689.080 ;
        RECT 1703.910 1689.020 1704.230 1689.080 ;
        RECT 1699.770 1688.880 1704.230 1689.020 ;
        RECT 1699.770 1688.820 1700.090 1688.880 ;
        RECT 1703.910 1688.820 1704.230 1688.880 ;
        RECT 1703.910 19.620 1704.230 19.680 ;
        RECT 2036.490 19.620 2036.810 19.680 ;
        RECT 1703.910 19.480 2036.810 19.620 ;
        RECT 1703.910 19.420 1704.230 19.480 ;
        RECT 2036.490 19.420 2036.810 19.480 ;
      LAYER via ;
        RECT 1699.800 1688.820 1700.060 1689.080 ;
        RECT 1703.940 1688.820 1704.200 1689.080 ;
        RECT 1703.940 19.420 1704.200 19.680 ;
        RECT 2036.520 19.420 2036.780 19.680 ;
      LAYER met2 ;
        RECT 1699.790 1700.000 1700.070 1704.000 ;
        RECT 1699.860 1689.110 1700.000 1700.000 ;
        RECT 1699.800 1688.790 1700.060 1689.110 ;
        RECT 1703.940 1688.790 1704.200 1689.110 ;
        RECT 1704.000 19.710 1704.140 1688.790 ;
        RECT 1703.940 19.390 1704.200 19.710 ;
        RECT 2036.520 19.390 2036.780 19.710 ;
        RECT 2036.580 2.400 2036.720 19.390 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 0.300 ;
=======
      LAYER li1 ;
        RECT 1725.145 14.025 1725.315 18.955 ;
        RECT 1772.985 14.875 1773.155 18.955 ;
        RECT 1773.445 15.725 1773.615 18.955 ;
        RECT 1785.865 15.725 1786.035 16.915 ;
        RECT 1797.365 16.745 1797.535 19.975 ;
        RECT 1824.965 17.425 1825.135 19.975 ;
        RECT 1873.265 17.425 1873.435 18.955 ;
        RECT 1918.345 16.065 1918.515 18.955 ;
        RECT 1966.185 16.065 1966.355 18.955 ;
        RECT 2028.285 18.615 2028.455 18.955 ;
        RECT 2029.205 18.615 2029.375 20.315 ;
        RECT 2028.285 18.445 2029.375 18.615 ;
        RECT 1772.525 14.705 1773.155 14.875 ;
      LAYER mcon ;
        RECT 2029.205 20.145 2029.375 20.315 ;
        RECT 1797.365 19.805 1797.535 19.975 ;
        RECT 1725.145 18.785 1725.315 18.955 ;
        RECT 1772.985 18.785 1773.155 18.955 ;
        RECT 1773.445 18.785 1773.615 18.955 ;
        RECT 1824.965 19.805 1825.135 19.975 ;
        RECT 1873.265 18.785 1873.435 18.955 ;
        RECT 1918.345 18.785 1918.515 18.955 ;
        RECT 1785.865 16.745 1786.035 16.915 ;
        RECT 1966.185 18.785 1966.355 18.955 ;
        RECT 2028.285 18.785 2028.455 18.955 ;
      LAYER met1 ;
        RECT 1704.370 1688.680 1704.690 1688.740 ;
        RECT 1710.350 1688.680 1710.670 1688.740 ;
        RECT 1704.370 1688.540 1710.670 1688.680 ;
        RECT 1704.370 1688.480 1704.690 1688.540 ;
        RECT 1710.350 1688.480 1710.670 1688.540 ;
        RECT 2029.145 20.300 2029.435 20.345 ;
        RECT 2054.430 20.300 2054.750 20.360 ;
        RECT 2029.145 20.160 2054.750 20.300 ;
        RECT 2029.145 20.115 2029.435 20.160 ;
        RECT 2054.430 20.100 2054.750 20.160 ;
        RECT 1797.305 19.960 1797.595 20.005 ;
        RECT 1824.905 19.960 1825.195 20.005 ;
        RECT 1797.305 19.820 1825.195 19.960 ;
        RECT 1797.305 19.775 1797.595 19.820 ;
        RECT 1824.905 19.775 1825.195 19.820 ;
        RECT 1710.350 18.940 1710.670 19.000 ;
        RECT 1725.085 18.940 1725.375 18.985 ;
        RECT 1710.350 18.800 1725.375 18.940 ;
        RECT 1710.350 18.740 1710.670 18.800 ;
        RECT 1725.085 18.755 1725.375 18.800 ;
        RECT 1772.925 18.940 1773.215 18.985 ;
        RECT 1773.385 18.940 1773.675 18.985 ;
        RECT 1772.925 18.800 1773.675 18.940 ;
        RECT 1772.925 18.755 1773.215 18.800 ;
        RECT 1773.385 18.755 1773.675 18.800 ;
        RECT 1873.205 18.940 1873.495 18.985 ;
        RECT 1918.285 18.940 1918.575 18.985 ;
        RECT 1873.205 18.800 1918.575 18.940 ;
        RECT 1873.205 18.755 1873.495 18.800 ;
        RECT 1918.285 18.755 1918.575 18.800 ;
        RECT 1966.125 18.940 1966.415 18.985 ;
        RECT 2028.225 18.940 2028.515 18.985 ;
        RECT 1966.125 18.800 2028.515 18.940 ;
        RECT 1966.125 18.755 1966.415 18.800 ;
        RECT 2028.225 18.755 2028.515 18.800 ;
        RECT 1824.905 17.580 1825.195 17.625 ;
        RECT 1873.205 17.580 1873.495 17.625 ;
        RECT 1824.905 17.440 1873.495 17.580 ;
        RECT 1824.905 17.395 1825.195 17.440 ;
        RECT 1873.205 17.395 1873.495 17.440 ;
        RECT 1785.805 16.900 1786.095 16.945 ;
        RECT 1797.305 16.900 1797.595 16.945 ;
        RECT 1785.805 16.760 1797.595 16.900 ;
        RECT 1785.805 16.715 1786.095 16.760 ;
        RECT 1797.305 16.715 1797.595 16.760 ;
        RECT 1918.285 16.220 1918.575 16.265 ;
        RECT 1966.125 16.220 1966.415 16.265 ;
        RECT 1918.285 16.080 1966.415 16.220 ;
        RECT 1918.285 16.035 1918.575 16.080 ;
        RECT 1966.125 16.035 1966.415 16.080 ;
        RECT 1773.385 15.880 1773.675 15.925 ;
        RECT 1785.805 15.880 1786.095 15.925 ;
        RECT 1773.385 15.740 1786.095 15.880 ;
        RECT 1773.385 15.695 1773.675 15.740 ;
        RECT 1785.805 15.695 1786.095 15.740 ;
        RECT 1772.465 14.860 1772.755 14.905 ;
        RECT 1733.900 14.720 1772.755 14.860 ;
        RECT 1725.085 14.180 1725.375 14.225 ;
        RECT 1733.900 14.180 1734.040 14.720 ;
        RECT 1772.465 14.675 1772.755 14.720 ;
        RECT 1725.085 14.040 1734.040 14.180 ;
        RECT 1725.085 13.995 1725.375 14.040 ;
      LAYER via ;
        RECT 1704.400 1688.480 1704.660 1688.740 ;
        RECT 1710.380 1688.480 1710.640 1688.740 ;
        RECT 2054.460 20.100 2054.720 20.360 ;
        RECT 1710.380 18.740 1710.640 19.000 ;
      LAYER met2 ;
        RECT 1704.390 1700.000 1704.670 1704.000 ;
        RECT 1704.460 1688.770 1704.600 1700.000 ;
        RECT 1704.400 1688.450 1704.660 1688.770 ;
        RECT 1710.380 1688.450 1710.640 1688.770 ;
        RECT 1710.440 19.030 1710.580 1688.450 ;
        RECT 2054.460 20.070 2054.720 20.390 ;
        RECT 1710.380 18.710 1710.640 19.030 ;
        RECT 2054.520 2.400 2054.660 20.070 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 0.300 ;
=======
      LAYER met1 ;
        RECT 769.650 48.180 769.970 48.240 ;
        RECT 1353.850 48.180 1354.170 48.240 ;
        RECT 769.650 48.040 1354.170 48.180 ;
        RECT 769.650 47.980 769.970 48.040 ;
        RECT 1353.850 47.980 1354.170 48.040 ;
      LAYER via ;
        RECT 769.680 47.980 769.940 48.240 ;
        RECT 1353.880 47.980 1354.140 48.240 ;
      LAYER met2 ;
        RECT 1357.550 1700.410 1357.830 1704.000 ;
        RECT 1356.240 1700.270 1357.830 1700.410 ;
        RECT 1356.240 1677.290 1356.380 1700.270 ;
        RECT 1357.550 1700.000 1357.830 1700.270 ;
        RECT 1353.940 1677.150 1356.380 1677.290 ;
        RECT 1353.940 48.270 1354.080 1677.150 ;
        RECT 769.680 47.950 769.940 48.270 ;
        RECT 1353.880 47.950 1354.140 48.270 ;
        RECT 769.740 2.400 769.880 47.950 ;
        RECT 769.530 -4.800 770.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 0.300 ;
=======
      LAYER li1 ;
        RECT 2038.865 16.405 2039.035 18.615 ;
      LAYER mcon ;
        RECT 2038.865 18.445 2039.035 18.615 ;
      LAYER met1 ;
        RECT 1709.430 1689.360 1709.750 1689.420 ;
        RECT 1710.810 1689.360 1711.130 1689.420 ;
        RECT 1709.430 1689.220 1711.130 1689.360 ;
        RECT 1709.430 1689.160 1709.750 1689.220 ;
        RECT 1710.810 1689.160 1711.130 1689.220 ;
        RECT 1710.810 18.600 1711.130 18.660 ;
        RECT 2038.805 18.600 2039.095 18.645 ;
        RECT 1710.810 18.460 2039.095 18.600 ;
        RECT 1710.810 18.400 1711.130 18.460 ;
        RECT 2038.805 18.415 2039.095 18.460 ;
        RECT 2038.805 16.560 2039.095 16.605 ;
        RECT 2072.370 16.560 2072.690 16.620 ;
        RECT 2038.805 16.420 2072.690 16.560 ;
        RECT 2038.805 16.375 2039.095 16.420 ;
        RECT 2072.370 16.360 2072.690 16.420 ;
      LAYER via ;
        RECT 1709.460 1689.160 1709.720 1689.420 ;
        RECT 1710.840 1689.160 1711.100 1689.420 ;
        RECT 1710.840 18.400 1711.100 18.660 ;
        RECT 2072.400 16.360 2072.660 16.620 ;
      LAYER met2 ;
        RECT 1709.450 1700.000 1709.730 1704.000 ;
        RECT 1709.520 1689.450 1709.660 1700.000 ;
        RECT 1709.460 1689.130 1709.720 1689.450 ;
        RECT 1710.840 1689.130 1711.100 1689.450 ;
        RECT 1710.900 18.690 1711.040 1689.130 ;
        RECT 1710.840 18.370 1711.100 18.690 ;
        RECT 2072.400 16.330 2072.660 16.650 ;
        RECT 2072.460 2.400 2072.600 16.330 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 0.300 ;
=======
      LAYER li1 ;
        RECT 2028.745 18.785 2028.915 20.315 ;
      LAYER mcon ;
        RECT 2028.745 20.145 2028.915 20.315 ;
      LAYER met1 ;
        RECT 1714.030 1690.380 1714.350 1690.440 ;
        RECT 2011.190 1690.380 2011.510 1690.440 ;
        RECT 1714.030 1690.240 2011.510 1690.380 ;
        RECT 1714.030 1690.180 1714.350 1690.240 ;
        RECT 2011.190 1690.180 2011.510 1690.240 ;
        RECT 2011.190 20.300 2011.510 20.360 ;
        RECT 2028.685 20.300 2028.975 20.345 ;
        RECT 2011.190 20.160 2028.975 20.300 ;
        RECT 2011.190 20.100 2011.510 20.160 ;
        RECT 2028.685 20.115 2028.975 20.160 ;
        RECT 2028.685 18.940 2028.975 18.985 ;
        RECT 2089.850 18.940 2090.170 19.000 ;
        RECT 2028.685 18.800 2090.170 18.940 ;
        RECT 2028.685 18.755 2028.975 18.800 ;
        RECT 2089.850 18.740 2090.170 18.800 ;
      LAYER via ;
        RECT 1714.060 1690.180 1714.320 1690.440 ;
        RECT 2011.220 1690.180 2011.480 1690.440 ;
        RECT 2011.220 20.100 2011.480 20.360 ;
        RECT 2089.880 18.740 2090.140 19.000 ;
      LAYER met2 ;
        RECT 1714.050 1700.000 1714.330 1704.000 ;
        RECT 1714.120 1690.470 1714.260 1700.000 ;
        RECT 1714.060 1690.150 1714.320 1690.470 ;
        RECT 2011.220 1690.150 2011.480 1690.470 ;
        RECT 2011.280 20.390 2011.420 1690.150 ;
        RECT 2011.220 20.070 2011.480 20.390 ;
        RECT 2089.880 18.710 2090.140 19.030 ;
        RECT 2089.940 2.400 2090.080 18.710 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 0.300 ;
=======
      LAYER li1 ;
        RECT 1965.725 16.405 1965.895 20.655 ;
      LAYER mcon ;
        RECT 1965.725 20.485 1965.895 20.655 ;
      LAYER met1 ;
        RECT 1719.090 1686.300 1719.410 1686.360 ;
        RECT 1924.710 1686.300 1925.030 1686.360 ;
        RECT 1942.190 1686.300 1942.510 1686.360 ;
        RECT 1719.090 1686.160 1897.800 1686.300 ;
        RECT 1719.090 1686.100 1719.410 1686.160 ;
        RECT 1897.660 1685.960 1897.800 1686.160 ;
        RECT 1924.710 1686.160 1942.510 1686.300 ;
        RECT 1924.710 1686.100 1925.030 1686.160 ;
        RECT 1942.190 1686.100 1942.510 1686.160 ;
        RECT 1898.490 1685.960 1898.810 1686.020 ;
        RECT 1897.660 1685.820 1898.810 1685.960 ;
        RECT 1898.490 1685.760 1898.810 1685.820 ;
        RECT 1965.665 20.640 1965.955 20.685 ;
        RECT 2107.790 20.640 2108.110 20.700 ;
        RECT 1965.665 20.500 2108.110 20.640 ;
        RECT 1965.665 20.455 1965.955 20.500 ;
        RECT 2107.790 20.440 2108.110 20.500 ;
        RECT 1942.190 16.560 1942.510 16.620 ;
        RECT 1965.665 16.560 1965.955 16.605 ;
        RECT 1942.190 16.420 1965.955 16.560 ;
        RECT 1942.190 16.360 1942.510 16.420 ;
        RECT 1965.665 16.375 1965.955 16.420 ;
      LAYER via ;
        RECT 1719.120 1686.100 1719.380 1686.360 ;
        RECT 1924.740 1686.100 1925.000 1686.360 ;
        RECT 1942.220 1686.100 1942.480 1686.360 ;
        RECT 1898.520 1685.760 1898.780 1686.020 ;
        RECT 2107.820 20.440 2108.080 20.700 ;
        RECT 1942.220 16.360 1942.480 16.620 ;
      LAYER met2 ;
        RECT 1719.110 1700.000 1719.390 1704.000 ;
        RECT 1719.180 1686.390 1719.320 1700.000 ;
        RECT 1719.120 1686.070 1719.380 1686.390 ;
        RECT 1924.740 1686.245 1925.000 1686.390 ;
        RECT 1898.510 1685.875 1898.790 1686.245 ;
        RECT 1924.730 1685.875 1925.010 1686.245 ;
        RECT 1942.220 1686.070 1942.480 1686.390 ;
        RECT 1898.520 1685.730 1898.780 1685.875 ;
        RECT 1942.280 16.650 1942.420 1686.070 ;
        RECT 2107.820 20.410 2108.080 20.730 ;
        RECT 1942.220 16.330 1942.480 16.650 ;
        RECT 2107.880 2.400 2108.020 20.410 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
      LAYER via2 ;
        RECT 1898.510 1685.920 1898.790 1686.200 ;
        RECT 1924.730 1685.920 1925.010 1686.200 ;
      LAYER met3 ;
        RECT 1898.485 1686.210 1898.815 1686.225 ;
        RECT 1924.705 1686.210 1925.035 1686.225 ;
        RECT 1898.485 1685.910 1925.035 1686.210 ;
        RECT 1898.485 1685.895 1898.815 1685.910 ;
        RECT 1924.705 1685.895 1925.035 1685.910 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1723.690 1689.700 1724.010 1689.760 ;
        RECT 2066.390 1689.700 2066.710 1689.760 ;
        RECT 1723.690 1689.560 2066.710 1689.700 ;
        RECT 1723.690 1689.500 1724.010 1689.560 ;
        RECT 2066.390 1689.500 2066.710 1689.560 ;
        RECT 2066.390 19.620 2066.710 19.680 ;
        RECT 2125.730 19.620 2126.050 19.680 ;
        RECT 2066.390 19.480 2126.050 19.620 ;
        RECT 2066.390 19.420 2066.710 19.480 ;
        RECT 2125.730 19.420 2126.050 19.480 ;
      LAYER via ;
        RECT 1723.720 1689.500 1723.980 1689.760 ;
        RECT 2066.420 1689.500 2066.680 1689.760 ;
        RECT 2066.420 19.420 2066.680 19.680 ;
        RECT 2125.760 19.420 2126.020 19.680 ;
      LAYER met2 ;
        RECT 1723.710 1700.000 1723.990 1704.000 ;
        RECT 1723.780 1689.790 1723.920 1700.000 ;
        RECT 1723.720 1689.470 1723.980 1689.790 ;
        RECT 2066.420 1689.470 2066.680 1689.790 ;
        RECT 2066.480 19.710 2066.620 1689.470 ;
        RECT 2066.420 19.390 2066.680 19.710 ;
        RECT 2125.760 19.390 2126.020 19.710 ;
        RECT 2125.820 2.400 2125.960 19.390 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1728.750 1688.680 1729.070 1688.740 ;
        RECT 1731.510 1688.680 1731.830 1688.740 ;
        RECT 1728.750 1688.540 1731.830 1688.680 ;
        RECT 1728.750 1688.480 1729.070 1688.540 ;
        RECT 1731.510 1688.480 1731.830 1688.540 ;
        RECT 1731.510 17.920 1731.830 17.980 ;
        RECT 2143.670 17.920 2143.990 17.980 ;
        RECT 1731.510 17.780 2143.990 17.920 ;
        RECT 1731.510 17.720 1731.830 17.780 ;
        RECT 2143.670 17.720 2143.990 17.780 ;
      LAYER via ;
        RECT 1728.780 1688.480 1729.040 1688.740 ;
        RECT 1731.540 1688.480 1731.800 1688.740 ;
        RECT 1731.540 17.720 1731.800 17.980 ;
        RECT 2143.700 17.720 2143.960 17.980 ;
      LAYER met2 ;
        RECT 1728.770 1700.000 1729.050 1704.000 ;
        RECT 1728.840 1688.770 1728.980 1700.000 ;
        RECT 1728.780 1688.450 1729.040 1688.770 ;
        RECT 1731.540 1688.450 1731.800 1688.770 ;
        RECT 1731.600 18.010 1731.740 1688.450 ;
        RECT 1731.540 17.690 1731.800 18.010 ;
        RECT 2143.700 17.690 2143.960 18.010 ;
        RECT 2143.760 2.400 2143.900 17.690 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 0.300 ;
=======
      LAYER li1 ;
        RECT 1771.605 1689.205 1772.695 1689.375 ;
        RECT 1771.605 1687.845 1771.775 1689.205 ;
      LAYER mcon ;
        RECT 1772.525 1689.205 1772.695 1689.375 ;
      LAYER met1 ;
        RECT 2159.770 1689.500 2160.090 1689.760 ;
        RECT 1772.465 1689.360 1772.755 1689.405 ;
        RECT 2159.860 1689.360 2160.000 1689.500 ;
        RECT 1772.465 1689.220 2160.000 1689.360 ;
        RECT 1772.465 1689.175 1772.755 1689.220 ;
        RECT 1733.350 1688.000 1733.670 1688.060 ;
        RECT 1771.545 1688.000 1771.835 1688.045 ;
        RECT 1733.350 1687.860 1771.835 1688.000 ;
        RECT 1733.350 1687.800 1733.670 1687.860 ;
        RECT 1771.545 1687.815 1771.835 1687.860 ;
      LAYER via ;
        RECT 2159.800 1689.500 2160.060 1689.760 ;
        RECT 1733.380 1687.800 1733.640 1688.060 ;
      LAYER met2 ;
        RECT 1733.370 1700.000 1733.650 1704.000 ;
        RECT 1733.440 1688.090 1733.580 1700.000 ;
        RECT 2159.800 1689.470 2160.060 1689.790 ;
        RECT 1733.380 1687.770 1733.640 1688.090 ;
        RECT 2159.860 17.410 2160.000 1689.470 ;
        RECT 2159.860 17.270 2161.840 17.410 ;
        RECT 2161.700 2.400 2161.840 17.270 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 0.300 ;
=======
      LAYER li1 ;
        RECT 2111.545 18.445 2111.715 20.655 ;
      LAYER mcon ;
        RECT 2111.545 20.485 2111.715 20.655 ;
      LAYER met1 ;
        RECT 1738.410 1690.040 1738.730 1690.100 ;
        RECT 2080.190 1690.040 2080.510 1690.100 ;
        RECT 1738.410 1689.900 2080.510 1690.040 ;
        RECT 1738.410 1689.840 1738.730 1689.900 ;
        RECT 2080.190 1689.840 2080.510 1689.900 ;
        RECT 2111.485 20.640 2111.775 20.685 ;
        RECT 2121.130 20.640 2121.450 20.700 ;
        RECT 2111.485 20.500 2121.450 20.640 ;
        RECT 2111.485 20.455 2111.775 20.500 ;
        RECT 2121.130 20.440 2121.450 20.500 ;
        RECT 2091.230 18.600 2091.550 18.660 ;
        RECT 2111.485 18.600 2111.775 18.645 ;
        RECT 2091.230 18.460 2111.775 18.600 ;
        RECT 2091.230 18.400 2091.550 18.460 ;
        RECT 2111.485 18.415 2111.775 18.460 ;
        RECT 2159.310 18.600 2159.630 18.660 ;
        RECT 2179.090 18.600 2179.410 18.660 ;
        RECT 2159.310 18.460 2179.410 18.600 ;
        RECT 2159.310 18.400 2159.630 18.460 ;
        RECT 2179.090 18.400 2179.410 18.460 ;
      LAYER via ;
        RECT 1738.440 1689.840 1738.700 1690.100 ;
        RECT 2080.220 1689.840 2080.480 1690.100 ;
        RECT 2121.160 20.440 2121.420 20.700 ;
        RECT 2091.260 18.400 2091.520 18.660 ;
        RECT 2159.340 18.400 2159.600 18.660 ;
        RECT 2179.120 18.400 2179.380 18.660 ;
      LAYER met2 ;
        RECT 1738.430 1700.000 1738.710 1704.000 ;
        RECT 1738.500 1690.130 1738.640 1700.000 ;
        RECT 1738.440 1689.810 1738.700 1690.130 ;
        RECT 2080.220 1689.810 2080.480 1690.130 ;
        RECT 2080.280 20.925 2080.420 1689.810 ;
        RECT 2080.210 20.555 2080.490 20.925 ;
        RECT 2091.250 20.555 2091.530 20.925 ;
        RECT 2121.150 20.555 2121.430 20.925 ;
        RECT 2159.330 20.555 2159.610 20.925 ;
        RECT 2091.320 18.690 2091.460 20.555 ;
        RECT 2121.160 20.410 2121.420 20.555 ;
        RECT 2159.400 18.690 2159.540 20.555 ;
        RECT 2091.260 18.370 2091.520 18.690 ;
        RECT 2159.340 18.370 2159.600 18.690 ;
        RECT 2179.120 18.370 2179.380 18.690 ;
        RECT 2179.180 2.400 2179.320 18.370 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
      LAYER via2 ;
        RECT 2080.210 20.600 2080.490 20.880 ;
        RECT 2091.250 20.600 2091.530 20.880 ;
        RECT 2121.150 20.600 2121.430 20.880 ;
        RECT 2159.330 20.600 2159.610 20.880 ;
      LAYER met3 ;
        RECT 2080.185 20.890 2080.515 20.905 ;
        RECT 2091.225 20.890 2091.555 20.905 ;
        RECT 2080.185 20.590 2091.555 20.890 ;
        RECT 2080.185 20.575 2080.515 20.590 ;
        RECT 2091.225 20.575 2091.555 20.590 ;
        RECT 2121.125 20.890 2121.455 20.905 ;
        RECT 2159.305 20.890 2159.635 20.905 ;
        RECT 2121.125 20.590 2159.635 20.890 ;
        RECT 2121.125 20.575 2121.455 20.590 ;
        RECT 2159.305 20.575 2159.635 20.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 0.300 ;
=======
      LAYER li1 ;
        RECT 1824.505 1686.825 1824.675 1689.035 ;
        RECT 1870.045 1688.865 1870.215 1691.075 ;
        RECT 1898.105 1688.865 1898.275 1691.075 ;
        RECT 1966.645 1686.145 1966.815 1689.035 ;
        RECT 2018.165 1686.145 2018.335 1689.035 ;
        RECT 2063.245 1688.865 2063.415 1690.395 ;
        RECT 2099.125 1688.865 2099.295 1690.395 ;
        RECT 2159.845 1686.485 2160.015 1689.035 ;
      LAYER mcon ;
        RECT 1870.045 1690.905 1870.215 1691.075 ;
        RECT 1824.505 1688.865 1824.675 1689.035 ;
        RECT 1898.105 1690.905 1898.275 1691.075 ;
        RECT 2063.245 1690.225 2063.415 1690.395 ;
        RECT 1966.645 1688.865 1966.815 1689.035 ;
        RECT 2018.165 1688.865 2018.335 1689.035 ;
        RECT 2099.125 1690.225 2099.295 1690.395 ;
        RECT 2159.845 1688.865 2160.015 1689.035 ;
      LAYER met1 ;
        RECT 1869.985 1691.060 1870.275 1691.105 ;
        RECT 1898.045 1691.060 1898.335 1691.105 ;
        RECT 1869.985 1690.920 1898.335 1691.060 ;
        RECT 1869.985 1690.875 1870.275 1690.920 ;
        RECT 1898.045 1690.875 1898.335 1690.920 ;
        RECT 2063.185 1690.380 2063.475 1690.425 ;
        RECT 2099.065 1690.380 2099.355 1690.425 ;
        RECT 2063.185 1690.240 2099.355 1690.380 ;
        RECT 2063.185 1690.195 2063.475 1690.240 ;
        RECT 2099.065 1690.195 2099.355 1690.240 ;
        RECT 1824.445 1689.020 1824.735 1689.065 ;
        RECT 1869.985 1689.020 1870.275 1689.065 ;
        RECT 1824.445 1688.880 1870.275 1689.020 ;
        RECT 1824.445 1688.835 1824.735 1688.880 ;
        RECT 1869.985 1688.835 1870.275 1688.880 ;
        RECT 1898.045 1689.020 1898.335 1689.065 ;
        RECT 1966.585 1689.020 1966.875 1689.065 ;
        RECT 1898.045 1688.880 1966.875 1689.020 ;
        RECT 1898.045 1688.835 1898.335 1688.880 ;
        RECT 1966.585 1688.835 1966.875 1688.880 ;
        RECT 2018.105 1689.020 2018.395 1689.065 ;
        RECT 2063.185 1689.020 2063.475 1689.065 ;
        RECT 2018.105 1688.880 2063.475 1689.020 ;
        RECT 2018.105 1688.835 2018.395 1688.880 ;
        RECT 2063.185 1688.835 2063.475 1688.880 ;
        RECT 2099.065 1689.020 2099.355 1689.065 ;
        RECT 2159.785 1689.020 2160.075 1689.065 ;
        RECT 2099.065 1688.880 2160.075 1689.020 ;
        RECT 2099.065 1688.835 2099.355 1688.880 ;
        RECT 2159.785 1688.835 2160.075 1688.880 ;
        RECT 1743.010 1687.320 1743.330 1687.380 ;
        RECT 1743.010 1687.180 1776.360 1687.320 ;
        RECT 1743.010 1687.120 1743.330 1687.180 ;
        RECT 1776.220 1686.640 1776.360 1687.180 ;
        RECT 1824.445 1686.980 1824.735 1687.025 ;
        RECT 1786.800 1686.840 1824.735 1686.980 ;
        RECT 1786.800 1686.640 1786.940 1686.840 ;
        RECT 1824.445 1686.795 1824.735 1686.840 ;
        RECT 1776.220 1686.500 1786.940 1686.640 ;
        RECT 2159.785 1686.640 2160.075 1686.685 ;
        RECT 2194.270 1686.640 2194.590 1686.700 ;
        RECT 2159.785 1686.500 2194.590 1686.640 ;
        RECT 2159.785 1686.455 2160.075 1686.500 ;
        RECT 2194.270 1686.440 2194.590 1686.500 ;
        RECT 1966.585 1686.300 1966.875 1686.345 ;
        RECT 2018.105 1686.300 2018.395 1686.345 ;
        RECT 1966.585 1686.160 2018.395 1686.300 ;
        RECT 1966.585 1686.115 1966.875 1686.160 ;
        RECT 2018.105 1686.115 2018.395 1686.160 ;
      LAYER via ;
        RECT 1743.040 1687.120 1743.300 1687.380 ;
        RECT 2194.300 1686.440 2194.560 1686.700 ;
      LAYER met2 ;
        RECT 1743.030 1700.000 1743.310 1704.000 ;
        RECT 1743.100 1687.410 1743.240 1700.000 ;
        RECT 1743.040 1687.090 1743.300 1687.410 ;
        RECT 2194.300 1686.410 2194.560 1686.730 ;
        RECT 2194.360 17.410 2194.500 1686.410 ;
        RECT 2194.360 17.270 2197.260 17.410 ;
        RECT 2197.120 2.400 2197.260 17.270 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1748.070 1689.020 1748.390 1689.080 ;
        RECT 1752.210 1689.020 1752.530 1689.080 ;
        RECT 1748.070 1688.880 1752.530 1689.020 ;
        RECT 1748.070 1688.820 1748.390 1688.880 ;
        RECT 1752.210 1688.820 1752.530 1688.880 ;
        RECT 1752.210 18.260 1752.530 18.320 ;
        RECT 2214.970 18.260 2215.290 18.320 ;
        RECT 1752.210 18.120 2215.290 18.260 ;
        RECT 1752.210 18.060 1752.530 18.120 ;
        RECT 2214.970 18.060 2215.290 18.120 ;
      LAYER via ;
        RECT 1748.100 1688.820 1748.360 1689.080 ;
        RECT 1752.240 1688.820 1752.500 1689.080 ;
        RECT 1752.240 18.060 1752.500 18.320 ;
        RECT 2215.000 18.060 2215.260 18.320 ;
      LAYER met2 ;
        RECT 1748.090 1700.000 1748.370 1704.000 ;
        RECT 1748.160 1689.110 1748.300 1700.000 ;
        RECT 1748.100 1688.790 1748.360 1689.110 ;
        RECT 1752.240 1688.790 1752.500 1689.110 ;
        RECT 1752.300 18.350 1752.440 1688.790 ;
        RECT 1752.240 18.030 1752.500 18.350 ;
        RECT 2215.000 18.030 2215.260 18.350 ;
        RECT 2215.060 2.400 2215.200 18.030 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1752.670 1689.020 1752.990 1689.080 ;
        RECT 1752.670 1688.880 1766.240 1689.020 ;
        RECT 1752.670 1688.820 1752.990 1688.880 ;
        RECT 1766.100 1688.680 1766.240 1688.880 ;
        RECT 2228.770 1688.680 2229.090 1688.740 ;
        RECT 1766.100 1688.540 2229.090 1688.680 ;
        RECT 2228.770 1688.480 2229.090 1688.540 ;
      LAYER via ;
        RECT 1752.700 1688.820 1752.960 1689.080 ;
        RECT 2228.800 1688.480 2229.060 1688.740 ;
      LAYER met2 ;
        RECT 1752.690 1700.000 1752.970 1704.000 ;
        RECT 1752.760 1689.110 1752.900 1700.000 ;
        RECT 1752.700 1688.790 1752.960 1689.110 ;
        RECT 2228.800 1688.450 2229.060 1688.770 ;
        RECT 2228.860 17.410 2229.000 1688.450 ;
        RECT 2228.860 17.270 2233.140 17.410 ;
        RECT 2233.000 2.400 2233.140 17.270 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 0.300 ;
=======
      LAYER met1 ;
        RECT 787.590 44.440 787.910 44.500 ;
        RECT 1360.290 44.440 1360.610 44.500 ;
        RECT 787.590 44.300 1360.610 44.440 ;
        RECT 787.590 44.240 787.910 44.300 ;
        RECT 1360.290 44.240 1360.610 44.300 ;
      LAYER via ;
        RECT 787.620 44.240 787.880 44.500 ;
        RECT 1360.320 44.240 1360.580 44.500 ;
      LAYER met2 ;
        RECT 1362.150 1700.410 1362.430 1704.000 ;
        RECT 1361.300 1700.270 1362.430 1700.410 ;
        RECT 1361.300 1677.970 1361.440 1700.270 ;
        RECT 1362.150 1700.000 1362.430 1700.270 ;
        RECT 1360.380 1677.830 1361.440 1677.970 ;
        RECT 1360.380 44.530 1360.520 1677.830 ;
        RECT 787.620 44.210 787.880 44.530 ;
        RECT 1360.320 44.210 1360.580 44.530 ;
        RECT 787.680 2.400 787.820 44.210 ;
        RECT 787.470 -4.800 788.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1757.270 1688.680 1757.590 1688.740 ;
        RECT 1759.110 1688.680 1759.430 1688.740 ;
        RECT 1757.270 1688.540 1759.430 1688.680 ;
        RECT 1757.270 1688.480 1757.590 1688.540 ;
        RECT 1759.110 1688.480 1759.430 1688.540 ;
        RECT 1759.110 14.180 1759.430 14.240 ;
        RECT 2250.850 14.180 2251.170 14.240 ;
        RECT 1759.110 14.040 2251.170 14.180 ;
        RECT 1759.110 13.980 1759.430 14.040 ;
        RECT 2250.850 13.980 2251.170 14.040 ;
      LAYER via ;
        RECT 1757.300 1688.480 1757.560 1688.740 ;
        RECT 1759.140 1688.480 1759.400 1688.740 ;
        RECT 1759.140 13.980 1759.400 14.240 ;
        RECT 2250.880 13.980 2251.140 14.240 ;
      LAYER met2 ;
        RECT 1757.290 1700.000 1757.570 1704.000 ;
        RECT 1757.360 1688.770 1757.500 1700.000 ;
        RECT 1757.300 1688.450 1757.560 1688.770 ;
        RECT 1759.140 1688.450 1759.400 1688.770 ;
        RECT 1759.200 14.270 1759.340 1688.450 ;
        RECT 1759.140 13.950 1759.400 14.270 ;
        RECT 2250.880 13.950 2251.140 14.270 ;
        RECT 2250.940 2.400 2251.080 13.950 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1762.330 1688.340 1762.650 1688.400 ;
        RECT 2252.690 1688.340 2253.010 1688.400 ;
        RECT 1762.330 1688.200 2253.010 1688.340 ;
        RECT 1762.330 1688.140 1762.650 1688.200 ;
        RECT 2252.690 1688.140 2253.010 1688.200 ;
        RECT 2252.690 14.180 2253.010 14.240 ;
        RECT 2268.330 14.180 2268.650 14.240 ;
        RECT 2252.690 14.040 2268.650 14.180 ;
        RECT 2252.690 13.980 2253.010 14.040 ;
        RECT 2268.330 13.980 2268.650 14.040 ;
      LAYER via ;
        RECT 1762.360 1688.140 1762.620 1688.400 ;
        RECT 2252.720 1688.140 2252.980 1688.400 ;
        RECT 2252.720 13.980 2252.980 14.240 ;
        RECT 2268.360 13.980 2268.620 14.240 ;
      LAYER met2 ;
        RECT 1762.350 1700.000 1762.630 1704.000 ;
        RECT 1762.420 1688.430 1762.560 1700.000 ;
        RECT 1762.360 1688.110 1762.620 1688.430 ;
        RECT 2252.720 1688.110 2252.980 1688.430 ;
        RECT 2252.780 14.270 2252.920 1688.110 ;
        RECT 2252.720 13.950 2252.980 14.270 ;
        RECT 2268.360 13.950 2268.620 14.270 ;
        RECT 2268.420 2.400 2268.560 13.950 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 0.300 ;
=======
      LAYER met1 ;
        RECT 1766.930 1686.980 1767.250 1687.040 ;
        RECT 1772.910 1686.980 1773.230 1687.040 ;
        RECT 1766.930 1686.840 1773.230 1686.980 ;
        RECT 1766.930 1686.780 1767.250 1686.840 ;
        RECT 1772.910 1686.780 1773.230 1686.840 ;
        RECT 1772.910 14.520 1773.230 14.580 ;
        RECT 2286.270 14.520 2286.590 14.580 ;
        RECT 1772.910 14.380 2286.590 14.520 ;
        RECT 1772.910 14.320 1773.230 14.380 ;
        RECT 2286.270 14.320 2286.590 14.380 ;
      LAYER via ;
        RECT 1766.960 1686.780 1767.220 1687.040 ;
        RECT 1772.940 1686.780 1773.200 1687.040 ;
        RECT 1772.940 14.320 1773.200 14.580 ;
        RECT 2286.300 14.320 2286.560 14.580 ;
      LAYER met2 ;
        RECT 1766.950 1700.000 1767.230 1704.000 ;
        RECT 1767.020 1687.070 1767.160 1700.000 ;
        RECT 1766.960 1686.750 1767.220 1687.070 ;
        RECT 1772.940 1686.750 1773.200 1687.070 ;
        RECT 1773.000 14.610 1773.140 1686.750 ;
        RECT 1772.940 14.290 1773.200 14.610 ;
        RECT 2286.300 14.290 2286.560 14.610 ;
        RECT 2286.360 2.400 2286.500 14.290 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1772.450 1688.000 1772.770 1688.060 ;
        RECT 2266.490 1688.000 2266.810 1688.060 ;
        RECT 1772.450 1687.860 2266.810 1688.000 ;
        RECT 1772.450 1687.800 1772.770 1687.860 ;
        RECT 2266.490 1687.800 2266.810 1687.860 ;
        RECT 2268.880 14.040 2300.300 14.180 ;
        RECT 2266.490 13.840 2266.810 13.900 ;
        RECT 2268.880 13.840 2269.020 14.040 ;
        RECT 2266.490 13.700 2269.020 13.840 ;
        RECT 2266.490 13.640 2266.810 13.700 ;
        RECT 2300.160 13.500 2300.300 14.040 ;
        RECT 2304.210 13.500 2304.530 13.560 ;
        RECT 2300.160 13.360 2304.530 13.500 ;
        RECT 2304.210 13.300 2304.530 13.360 ;
      LAYER via ;
        RECT 1772.480 1687.800 1772.740 1688.060 ;
        RECT 2266.520 1687.800 2266.780 1688.060 ;
        RECT 2266.520 13.640 2266.780 13.900 ;
        RECT 2304.240 13.300 2304.500 13.560 ;
      LAYER met2 ;
        RECT 1772.010 1700.410 1772.290 1704.000 ;
        RECT 1772.010 1700.270 1772.680 1700.410 ;
        RECT 1772.010 1700.000 1772.290 1700.270 ;
        RECT 1772.540 1688.090 1772.680 1700.270 ;
        RECT 1772.480 1687.770 1772.740 1688.090 ;
        RECT 2266.520 1687.770 2266.780 1688.090 ;
        RECT 2266.580 13.930 2266.720 1687.770 ;
        RECT 2266.520 13.610 2266.780 13.930 ;
        RECT 2304.240 13.270 2304.500 13.590 ;
        RECT 2304.300 2.400 2304.440 13.270 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1776.590 1687.320 1776.910 1687.380 ;
        RECT 1779.810 1687.320 1780.130 1687.380 ;
        RECT 1776.590 1687.180 1780.130 1687.320 ;
        RECT 1776.590 1687.120 1776.910 1687.180 ;
        RECT 1779.810 1687.120 1780.130 1687.180 ;
        RECT 1779.810 14.860 1780.130 14.920 ;
        RECT 2322.150 14.860 2322.470 14.920 ;
        RECT 1779.810 14.720 2322.470 14.860 ;
        RECT 1779.810 14.660 1780.130 14.720 ;
        RECT 2322.150 14.660 2322.470 14.720 ;
      LAYER via ;
        RECT 1776.620 1687.120 1776.880 1687.380 ;
        RECT 1779.840 1687.120 1780.100 1687.380 ;
        RECT 1779.840 14.660 1780.100 14.920 ;
        RECT 2322.180 14.660 2322.440 14.920 ;
      LAYER met2 ;
        RECT 1776.610 1700.000 1776.890 1704.000 ;
        RECT 1776.680 1687.410 1776.820 1700.000 ;
        RECT 1776.620 1687.090 1776.880 1687.410 ;
        RECT 1779.840 1687.090 1780.100 1687.410 ;
        RECT 1779.900 14.950 1780.040 1687.090 ;
        RECT 1779.840 14.630 1780.100 14.950 ;
        RECT 2322.180 14.630 2322.440 14.950 ;
        RECT 2322.240 2.400 2322.380 14.630 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 0.300 ;
=======
      LAYER li1 ;
        RECT 1824.965 1685.465 1825.135 1687.675 ;
      LAYER mcon ;
        RECT 1824.965 1687.505 1825.135 1687.675 ;
      LAYER met1 ;
        RECT 1824.905 1687.660 1825.195 1687.705 ;
        RECT 2287.190 1687.660 2287.510 1687.720 ;
        RECT 1824.905 1687.520 2287.510 1687.660 ;
        RECT 1824.905 1687.475 1825.195 1687.520 ;
        RECT 2287.190 1687.460 2287.510 1687.520 ;
        RECT 1781.650 1685.620 1781.970 1685.680 ;
        RECT 1824.905 1685.620 1825.195 1685.665 ;
        RECT 1781.650 1685.480 1825.195 1685.620 ;
        RECT 1781.650 1685.420 1781.970 1685.480 ;
        RECT 1824.905 1685.435 1825.195 1685.480 ;
        RECT 2287.190 14.520 2287.510 14.580 ;
        RECT 2287.190 14.380 2300.760 14.520 ;
        RECT 2287.190 14.320 2287.510 14.380 ;
        RECT 2300.620 13.840 2300.760 14.380 ;
        RECT 2339.630 14.180 2339.950 14.240 ;
        RECT 2304.760 14.040 2339.950 14.180 ;
        RECT 2304.760 13.840 2304.900 14.040 ;
        RECT 2339.630 13.980 2339.950 14.040 ;
        RECT 2300.620 13.700 2304.900 13.840 ;
      LAYER via ;
        RECT 2287.220 1687.460 2287.480 1687.720 ;
        RECT 1781.680 1685.420 1781.940 1685.680 ;
        RECT 2287.220 14.320 2287.480 14.580 ;
        RECT 2339.660 13.980 2339.920 14.240 ;
      LAYER met2 ;
        RECT 1781.670 1700.000 1781.950 1704.000 ;
        RECT 1781.740 1685.710 1781.880 1700.000 ;
        RECT 2287.220 1687.430 2287.480 1687.750 ;
        RECT 1781.680 1685.390 1781.940 1685.710 ;
        RECT 2287.280 14.610 2287.420 1687.430 ;
        RECT 2287.220 14.290 2287.480 14.610 ;
        RECT 2339.660 13.950 2339.920 14.270 ;
        RECT 2339.720 2.400 2339.860 13.950 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1786.250 15.880 1786.570 15.940 ;
        RECT 2357.570 15.880 2357.890 15.940 ;
        RECT 1786.250 15.740 2357.890 15.880 ;
        RECT 1786.250 15.680 1786.570 15.740 ;
        RECT 2357.570 15.680 2357.890 15.740 ;
      LAYER via ;
        RECT 1786.280 15.680 1786.540 15.940 ;
        RECT 2357.600 15.680 2357.860 15.940 ;
      LAYER met2 ;
        RECT 1786.270 1700.410 1786.550 1704.000 ;
        RECT 1786.270 1700.270 1786.940 1700.410 ;
        RECT 1786.270 1700.000 1786.550 1700.270 ;
        RECT 1786.800 24.890 1786.940 1700.270 ;
        RECT 1786.340 24.750 1786.940 24.890 ;
        RECT 1786.340 15.970 1786.480 24.750 ;
        RECT 1786.280 15.650 1786.540 15.970 ;
        RECT 2357.600 15.650 2357.860 15.970 ;
        RECT 2357.660 2.400 2357.800 15.650 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 0.300 ;
=======
      LAYER li1 ;
        RECT 1816.685 1685.805 1816.855 1687.335 ;
      LAYER mcon ;
        RECT 1816.685 1687.165 1816.855 1687.335 ;
      LAYER met1 ;
        RECT 1816.625 1687.320 1816.915 1687.365 ;
        RECT 2300.990 1687.320 2301.310 1687.380 ;
        RECT 1816.625 1687.180 2301.310 1687.320 ;
        RECT 1816.625 1687.135 1816.915 1687.180 ;
        RECT 2300.990 1687.120 2301.310 1687.180 ;
        RECT 1791.310 1685.960 1791.630 1686.020 ;
        RECT 1816.625 1685.960 1816.915 1686.005 ;
        RECT 1791.310 1685.820 1816.915 1685.960 ;
        RECT 1791.310 1685.760 1791.630 1685.820 ;
        RECT 1816.625 1685.775 1816.915 1685.820 ;
        RECT 2300.990 14.520 2301.310 14.580 ;
        RECT 2375.510 14.520 2375.830 14.580 ;
        RECT 2300.990 14.380 2375.830 14.520 ;
        RECT 2300.990 14.320 2301.310 14.380 ;
        RECT 2375.510 14.320 2375.830 14.380 ;
      LAYER via ;
        RECT 2301.020 1687.120 2301.280 1687.380 ;
        RECT 1791.340 1685.760 1791.600 1686.020 ;
        RECT 2301.020 14.320 2301.280 14.580 ;
        RECT 2375.540 14.320 2375.800 14.580 ;
      LAYER met2 ;
        RECT 1791.330 1700.000 1791.610 1704.000 ;
        RECT 1791.400 1686.050 1791.540 1700.000 ;
        RECT 2301.020 1687.090 2301.280 1687.410 ;
        RECT 1791.340 1685.730 1791.600 1686.050 ;
        RECT 2301.080 14.610 2301.220 1687.090 ;
        RECT 2301.020 14.290 2301.280 14.610 ;
        RECT 2375.540 14.290 2375.800 14.610 ;
        RECT 2375.600 2.400 2375.740 14.290 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 0.300 ;
=======
      LAYER met1 ;
        RECT 1795.910 1687.320 1796.230 1687.380 ;
        RECT 1800.510 1687.320 1800.830 1687.380 ;
        RECT 1795.910 1687.180 1800.830 1687.320 ;
        RECT 1795.910 1687.120 1796.230 1687.180 ;
        RECT 1800.510 1687.120 1800.830 1687.180 ;
        RECT 1800.510 16.900 1800.830 16.960 ;
        RECT 2393.450 16.900 2393.770 16.960 ;
        RECT 1800.510 16.760 2393.770 16.900 ;
        RECT 1800.510 16.700 1800.830 16.760 ;
        RECT 2393.450 16.700 2393.770 16.760 ;
      LAYER via ;
        RECT 1795.940 1687.120 1796.200 1687.380 ;
        RECT 1800.540 1687.120 1800.800 1687.380 ;
        RECT 1800.540 16.700 1800.800 16.960 ;
        RECT 2393.480 16.700 2393.740 16.960 ;
      LAYER met2 ;
        RECT 1795.930 1700.000 1796.210 1704.000 ;
        RECT 1796.000 1687.410 1796.140 1700.000 ;
        RECT 1795.940 1687.090 1796.200 1687.410 ;
        RECT 1800.540 1687.090 1800.800 1687.410 ;
        RECT 1800.600 16.990 1800.740 1687.090 ;
        RECT 1800.540 16.670 1800.800 16.990 ;
        RECT 2393.480 16.670 2393.740 16.990 ;
        RECT 2393.540 2.400 2393.680 16.670 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 0.300 ;
=======
      LAYER met1 ;
        RECT 2321.690 1686.980 2322.010 1687.040 ;
        RECT 1824.980 1686.840 2322.010 1686.980 ;
        RECT 1800.970 1686.640 1801.290 1686.700 ;
        RECT 1824.980 1686.640 1825.120 1686.840 ;
        RECT 2321.690 1686.780 2322.010 1686.840 ;
        RECT 1800.970 1686.500 1825.120 1686.640 ;
        RECT 1800.970 1686.440 1801.290 1686.500 ;
        RECT 2322.610 14.860 2322.930 14.920 ;
        RECT 2411.390 14.860 2411.710 14.920 ;
        RECT 2322.610 14.720 2411.710 14.860 ;
        RECT 2322.610 14.660 2322.930 14.720 ;
        RECT 2411.390 14.660 2411.710 14.720 ;
      LAYER via ;
        RECT 1801.000 1686.440 1801.260 1686.700 ;
        RECT 2321.720 1686.780 2321.980 1687.040 ;
        RECT 2322.640 14.660 2322.900 14.920 ;
        RECT 2411.420 14.660 2411.680 14.920 ;
      LAYER met2 ;
        RECT 1800.990 1700.000 1801.270 1704.000 ;
        RECT 1801.060 1686.730 1801.200 1700.000 ;
        RECT 2321.720 1686.750 2321.980 1687.070 ;
        RECT 1801.000 1686.410 1801.260 1686.730 ;
        RECT 2321.780 24.890 2321.920 1686.750 ;
        RECT 2321.780 24.750 2322.840 24.890 ;
        RECT 2322.700 14.950 2322.840 24.750 ;
        RECT 2322.640 14.630 2322.900 14.950 ;
        RECT 2411.420 14.630 2411.680 14.950 ;
        RECT 2411.480 2.400 2411.620 14.630 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 0.300 ;
=======
      LAYER met1 ;
        RECT 805.530 44.100 805.850 44.160 ;
        RECT 1367.190 44.100 1367.510 44.160 ;
        RECT 805.530 43.960 1367.510 44.100 ;
        RECT 805.530 43.900 805.850 43.960 ;
        RECT 1367.190 43.900 1367.510 43.960 ;
      LAYER via ;
        RECT 805.560 43.900 805.820 44.160 ;
        RECT 1367.220 43.900 1367.480 44.160 ;
      LAYER met2 ;
        RECT 1367.210 1700.000 1367.490 1704.000 ;
        RECT 1367.280 44.190 1367.420 1700.000 ;
        RECT 805.560 43.870 805.820 44.190 ;
        RECT 1367.220 43.870 1367.480 44.190 ;
        RECT 805.620 2.400 805.760 43.870 ;
        RECT 805.410 -4.800 805.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 0.300 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 0.300 ;
=======
      LAYER met1 ;
        RECT 2.830 24.040 3.150 24.100 ;
        RECT 1145.470 24.040 1145.790 24.100 ;
        RECT 2.830 23.900 1145.790 24.040 ;
        RECT 2.830 23.840 3.150 23.900 ;
        RECT 1145.470 23.840 1145.790 23.900 ;
      LAYER via ;
        RECT 2.860 23.840 3.120 24.100 ;
        RECT 1145.500 23.840 1145.760 24.100 ;
      LAYER met2 ;
        RECT 1150.550 1700.410 1150.830 1704.000 ;
        RECT 1145.560 1700.270 1150.830 1700.410 ;
        RECT 1145.560 24.130 1145.700 1700.270 ;
        RECT 1150.550 1700.000 1150.830 1700.270 ;
        RECT 2.860 23.810 3.120 24.130 ;
        RECT 1145.500 23.810 1145.760 24.130 ;
        RECT 2.920 2.400 3.060 23.810 ;
        RECT 2.710 -4.800 3.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 0.300 ;
=======
      LAYER li1 ;
        RECT 1147.385 1510.365 1147.555 1579.895 ;
        RECT 1146.465 1400.885 1146.635 1463.615 ;
        RECT 1147.385 1352.605 1147.555 1376.915 ;
        RECT 1146.925 1268.965 1147.095 1304.155 ;
        RECT 1146.465 917.745 1146.635 961.775 ;
        RECT 1146.465 531.505 1146.635 579.615 ;
        RECT 1146.465 434.945 1146.635 483.055 ;
        RECT 1146.465 338.045 1146.635 386.155 ;
        RECT 1146.465 241.485 1146.635 289.255 ;
        RECT 1146.925 193.205 1147.095 207.655 ;
        RECT 1146.005 138.125 1146.175 162.095 ;
      LAYER mcon ;
        RECT 1147.385 1579.725 1147.555 1579.895 ;
        RECT 1146.465 1463.445 1146.635 1463.615 ;
        RECT 1147.385 1376.745 1147.555 1376.915 ;
        RECT 1146.925 1303.985 1147.095 1304.155 ;
        RECT 1146.465 961.605 1146.635 961.775 ;
        RECT 1146.465 579.445 1146.635 579.615 ;
        RECT 1146.465 482.885 1146.635 483.055 ;
        RECT 1146.465 385.985 1146.635 386.155 ;
        RECT 1146.465 289.085 1146.635 289.255 ;
        RECT 1146.925 207.485 1147.095 207.655 ;
        RECT 1146.005 161.925 1146.175 162.095 ;
      LAYER met1 ;
        RECT 1147.310 1676.780 1147.630 1676.840 ;
        RECT 1151.910 1676.780 1152.230 1676.840 ;
        RECT 1147.310 1676.640 1152.230 1676.780 ;
        RECT 1147.310 1676.580 1147.630 1676.640 ;
        RECT 1151.910 1676.580 1152.230 1676.640 ;
        RECT 1146.390 1580.560 1146.710 1580.620 ;
        RECT 1147.310 1580.560 1147.630 1580.620 ;
        RECT 1146.390 1580.420 1147.630 1580.560 ;
        RECT 1146.390 1580.360 1146.710 1580.420 ;
        RECT 1147.310 1580.360 1147.630 1580.420 ;
        RECT 1147.310 1579.880 1147.630 1579.940 ;
        RECT 1147.115 1579.740 1147.630 1579.880 ;
        RECT 1147.310 1579.680 1147.630 1579.740 ;
        RECT 1147.310 1510.520 1147.630 1510.580 ;
        RECT 1147.115 1510.380 1147.630 1510.520 ;
        RECT 1147.310 1510.320 1147.630 1510.380 ;
        RECT 1146.405 1463.600 1146.695 1463.645 ;
        RECT 1147.310 1463.600 1147.630 1463.660 ;
        RECT 1146.405 1463.460 1147.630 1463.600 ;
        RECT 1146.405 1463.415 1146.695 1463.460 ;
        RECT 1147.310 1463.400 1147.630 1463.460 ;
        RECT 1146.405 1401.040 1146.695 1401.085 ;
        RECT 1147.310 1401.040 1147.630 1401.100 ;
        RECT 1146.405 1400.900 1147.630 1401.040 ;
        RECT 1146.405 1400.855 1146.695 1400.900 ;
        RECT 1147.310 1400.840 1147.630 1400.900 ;
        RECT 1147.310 1376.900 1147.630 1376.960 ;
        RECT 1147.115 1376.760 1147.630 1376.900 ;
        RECT 1147.310 1376.700 1147.630 1376.760 ;
        RECT 1146.390 1352.760 1146.710 1352.820 ;
        RECT 1147.325 1352.760 1147.615 1352.805 ;
        RECT 1146.390 1352.620 1147.615 1352.760 ;
        RECT 1146.390 1352.560 1146.710 1352.620 ;
        RECT 1147.325 1352.575 1147.615 1352.620 ;
        RECT 1146.390 1317.880 1146.710 1318.140 ;
        RECT 1146.480 1317.740 1146.620 1317.880 ;
        RECT 1146.850 1317.740 1147.170 1317.800 ;
        RECT 1146.480 1317.600 1147.170 1317.740 ;
        RECT 1146.850 1317.540 1147.170 1317.600 ;
        RECT 1146.850 1304.140 1147.170 1304.200 ;
        RECT 1146.655 1304.000 1147.170 1304.140 ;
        RECT 1146.850 1303.940 1147.170 1304.000 ;
        RECT 1146.850 1269.120 1147.170 1269.180 ;
        RECT 1146.655 1268.980 1147.170 1269.120 ;
        RECT 1146.850 1268.920 1147.170 1268.980 ;
        RECT 1146.850 1221.860 1147.170 1221.920 ;
        RECT 1146.480 1221.720 1147.170 1221.860 ;
        RECT 1146.480 1221.240 1146.620 1221.720 ;
        RECT 1146.850 1221.660 1147.170 1221.720 ;
        RECT 1146.390 1220.980 1146.710 1221.240 ;
        RECT 1146.850 1152.500 1147.170 1152.560 ;
        RECT 1147.770 1152.500 1148.090 1152.560 ;
        RECT 1146.850 1152.360 1148.090 1152.500 ;
        RECT 1146.850 1152.300 1147.170 1152.360 ;
        RECT 1147.770 1152.300 1148.090 1152.360 ;
        RECT 1146.850 1125.300 1147.170 1125.360 ;
        RECT 1146.480 1125.160 1147.170 1125.300 ;
        RECT 1146.480 1124.680 1146.620 1125.160 ;
        RECT 1146.850 1125.100 1147.170 1125.160 ;
        RECT 1146.390 1124.420 1146.710 1124.680 ;
        RECT 1147.310 1027.720 1147.630 1027.780 ;
        RECT 1148.230 1027.720 1148.550 1027.780 ;
        RECT 1147.310 1027.580 1148.550 1027.720 ;
        RECT 1147.310 1027.520 1147.630 1027.580 ;
        RECT 1148.230 1027.520 1148.550 1027.580 ;
        RECT 1146.390 980.120 1146.710 980.180 ;
        RECT 1147.310 980.120 1147.630 980.180 ;
        RECT 1146.390 979.980 1147.630 980.120 ;
        RECT 1146.390 979.920 1146.710 979.980 ;
        RECT 1147.310 979.920 1147.630 979.980 ;
        RECT 1146.390 961.760 1146.710 961.820 ;
        RECT 1146.195 961.620 1146.710 961.760 ;
        RECT 1146.390 961.560 1146.710 961.620 ;
        RECT 1146.405 917.900 1146.695 917.945 ;
        RECT 1146.850 917.900 1147.170 917.960 ;
        RECT 1146.405 917.760 1147.170 917.900 ;
        RECT 1146.405 917.715 1146.695 917.760 ;
        RECT 1146.850 917.700 1147.170 917.760 ;
        RECT 1146.850 883.700 1147.170 883.960 ;
        RECT 1146.940 882.940 1147.080 883.700 ;
        RECT 1146.850 882.680 1147.170 882.940 ;
        RECT 1146.390 786.800 1146.710 787.060 ;
        RECT 1146.480 786.660 1146.620 786.800 ;
        RECT 1146.850 786.660 1147.170 786.720 ;
        RECT 1146.480 786.520 1147.170 786.660 ;
        RECT 1146.850 786.460 1147.170 786.520 ;
        RECT 1146.850 772.720 1147.170 772.780 ;
        RECT 1147.770 772.720 1148.090 772.780 ;
        RECT 1146.850 772.580 1148.090 772.720 ;
        RECT 1146.850 772.520 1147.170 772.580 ;
        RECT 1147.770 772.520 1148.090 772.580 ;
        RECT 1146.390 689.900 1146.710 690.160 ;
        RECT 1146.480 689.760 1146.620 689.900 ;
        RECT 1146.850 689.760 1147.170 689.820 ;
        RECT 1146.480 689.620 1147.170 689.760 ;
        RECT 1146.850 689.560 1147.170 689.620 ;
        RECT 1146.850 676.160 1147.170 676.220 ;
        RECT 1147.770 676.160 1148.090 676.220 ;
        RECT 1146.850 676.020 1148.090 676.160 ;
        RECT 1146.850 675.960 1147.170 676.020 ;
        RECT 1147.770 675.960 1148.090 676.020 ;
        RECT 1146.390 593.340 1146.710 593.600 ;
        RECT 1146.480 593.200 1146.620 593.340 ;
        RECT 1146.850 593.200 1147.170 593.260 ;
        RECT 1146.480 593.060 1147.170 593.200 ;
        RECT 1146.850 593.000 1147.170 593.060 ;
        RECT 1146.405 579.600 1146.695 579.645 ;
        RECT 1146.850 579.600 1147.170 579.660 ;
        RECT 1146.405 579.460 1147.170 579.600 ;
        RECT 1146.405 579.415 1146.695 579.460 ;
        RECT 1146.850 579.400 1147.170 579.460 ;
        RECT 1146.390 531.660 1146.710 531.720 ;
        RECT 1146.195 531.520 1146.710 531.660 ;
        RECT 1146.390 531.460 1146.710 531.520 ;
        RECT 1146.390 496.780 1146.710 497.040 ;
        RECT 1146.480 496.640 1146.620 496.780 ;
        RECT 1146.850 496.640 1147.170 496.700 ;
        RECT 1146.480 496.500 1147.170 496.640 ;
        RECT 1146.850 496.440 1147.170 496.500 ;
        RECT 1146.405 483.040 1146.695 483.085 ;
        RECT 1146.850 483.040 1147.170 483.100 ;
        RECT 1146.405 482.900 1147.170 483.040 ;
        RECT 1146.405 482.855 1146.695 482.900 ;
        RECT 1146.850 482.840 1147.170 482.900 ;
        RECT 1146.390 435.100 1146.710 435.160 ;
        RECT 1146.195 434.960 1146.710 435.100 ;
        RECT 1146.390 434.900 1146.710 434.960 ;
        RECT 1146.390 400.220 1146.710 400.480 ;
        RECT 1146.480 399.740 1146.620 400.220 ;
        RECT 1146.850 399.740 1147.170 399.800 ;
        RECT 1146.480 399.600 1147.170 399.740 ;
        RECT 1146.850 399.540 1147.170 399.600 ;
        RECT 1146.405 386.140 1146.695 386.185 ;
        RECT 1146.850 386.140 1147.170 386.200 ;
        RECT 1146.405 386.000 1147.170 386.140 ;
        RECT 1146.405 385.955 1146.695 386.000 ;
        RECT 1146.850 385.940 1147.170 386.000 ;
        RECT 1146.390 338.200 1146.710 338.260 ;
        RECT 1146.195 338.060 1146.710 338.200 ;
        RECT 1146.390 338.000 1146.710 338.060 ;
        RECT 1146.390 289.920 1146.710 289.980 ;
        RECT 1146.850 289.920 1147.170 289.980 ;
        RECT 1146.390 289.780 1147.170 289.920 ;
        RECT 1146.390 289.720 1146.710 289.780 ;
        RECT 1146.850 289.720 1147.170 289.780 ;
        RECT 1146.390 289.240 1146.710 289.300 ;
        RECT 1146.195 289.100 1146.710 289.240 ;
        RECT 1146.390 289.040 1146.710 289.100 ;
        RECT 1146.405 241.640 1146.695 241.685 ;
        RECT 1146.850 241.640 1147.170 241.700 ;
        RECT 1146.405 241.500 1147.170 241.640 ;
        RECT 1146.405 241.455 1146.695 241.500 ;
        RECT 1146.850 241.440 1147.170 241.500 ;
        RECT 1146.850 207.640 1147.170 207.700 ;
        RECT 1146.655 207.500 1147.170 207.640 ;
        RECT 1146.850 207.440 1147.170 207.500 ;
        RECT 1145.930 193.360 1146.250 193.420 ;
        RECT 1146.865 193.360 1147.155 193.405 ;
        RECT 1145.930 193.220 1147.155 193.360 ;
        RECT 1145.930 193.160 1146.250 193.220 ;
        RECT 1146.865 193.175 1147.155 193.220 ;
        RECT 1145.930 162.080 1146.250 162.140 ;
        RECT 1145.735 161.940 1146.250 162.080 ;
        RECT 1145.930 161.880 1146.250 161.940 ;
        RECT 1145.945 138.280 1146.235 138.325 ;
        RECT 1146.850 138.280 1147.170 138.340 ;
        RECT 1145.945 138.140 1147.170 138.280 ;
        RECT 1145.945 138.095 1146.235 138.140 ;
        RECT 1146.850 138.080 1147.170 138.140 ;
        RECT 1146.850 110.740 1147.170 110.800 ;
        RECT 1146.480 110.600 1147.170 110.740 ;
        RECT 1146.480 110.460 1146.620 110.600 ;
        RECT 1146.850 110.540 1147.170 110.600 ;
        RECT 1146.390 110.200 1146.710 110.460 ;
        RECT 8.350 24.720 8.670 24.780 ;
        RECT 1145.930 24.720 1146.250 24.780 ;
        RECT 8.350 24.580 1146.250 24.720 ;
        RECT 8.350 24.520 8.670 24.580 ;
        RECT 1145.930 24.520 1146.250 24.580 ;
      LAYER via ;
        RECT 1147.340 1676.580 1147.600 1676.840 ;
        RECT 1151.940 1676.580 1152.200 1676.840 ;
        RECT 1146.420 1580.360 1146.680 1580.620 ;
        RECT 1147.340 1580.360 1147.600 1580.620 ;
        RECT 1147.340 1579.680 1147.600 1579.940 ;
        RECT 1147.340 1510.320 1147.600 1510.580 ;
        RECT 1147.340 1463.400 1147.600 1463.660 ;
        RECT 1147.340 1400.840 1147.600 1401.100 ;
        RECT 1147.340 1376.700 1147.600 1376.960 ;
        RECT 1146.420 1352.560 1146.680 1352.820 ;
        RECT 1146.420 1317.880 1146.680 1318.140 ;
        RECT 1146.880 1317.540 1147.140 1317.800 ;
        RECT 1146.880 1303.940 1147.140 1304.200 ;
        RECT 1146.880 1268.920 1147.140 1269.180 ;
        RECT 1146.880 1221.660 1147.140 1221.920 ;
        RECT 1146.420 1220.980 1146.680 1221.240 ;
        RECT 1146.880 1152.300 1147.140 1152.560 ;
        RECT 1147.800 1152.300 1148.060 1152.560 ;
        RECT 1146.880 1125.100 1147.140 1125.360 ;
        RECT 1146.420 1124.420 1146.680 1124.680 ;
        RECT 1147.340 1027.520 1147.600 1027.780 ;
        RECT 1148.260 1027.520 1148.520 1027.780 ;
        RECT 1146.420 979.920 1146.680 980.180 ;
        RECT 1147.340 979.920 1147.600 980.180 ;
        RECT 1146.420 961.560 1146.680 961.820 ;
        RECT 1146.880 917.700 1147.140 917.960 ;
        RECT 1146.880 883.700 1147.140 883.960 ;
        RECT 1146.880 882.680 1147.140 882.940 ;
        RECT 1146.420 786.800 1146.680 787.060 ;
        RECT 1146.880 786.460 1147.140 786.720 ;
        RECT 1146.880 772.520 1147.140 772.780 ;
        RECT 1147.800 772.520 1148.060 772.780 ;
        RECT 1146.420 689.900 1146.680 690.160 ;
        RECT 1146.880 689.560 1147.140 689.820 ;
        RECT 1146.880 675.960 1147.140 676.220 ;
        RECT 1147.800 675.960 1148.060 676.220 ;
        RECT 1146.420 593.340 1146.680 593.600 ;
        RECT 1146.880 593.000 1147.140 593.260 ;
        RECT 1146.880 579.400 1147.140 579.660 ;
        RECT 1146.420 531.460 1146.680 531.720 ;
        RECT 1146.420 496.780 1146.680 497.040 ;
        RECT 1146.880 496.440 1147.140 496.700 ;
        RECT 1146.880 482.840 1147.140 483.100 ;
        RECT 1146.420 434.900 1146.680 435.160 ;
        RECT 1146.420 400.220 1146.680 400.480 ;
        RECT 1146.880 399.540 1147.140 399.800 ;
        RECT 1146.880 385.940 1147.140 386.200 ;
        RECT 1146.420 338.000 1146.680 338.260 ;
        RECT 1146.420 289.720 1146.680 289.980 ;
        RECT 1146.880 289.720 1147.140 289.980 ;
        RECT 1146.420 289.040 1146.680 289.300 ;
        RECT 1146.880 241.440 1147.140 241.700 ;
        RECT 1146.880 207.440 1147.140 207.700 ;
        RECT 1145.960 193.160 1146.220 193.420 ;
        RECT 1145.960 161.880 1146.220 162.140 ;
        RECT 1146.880 138.080 1147.140 138.340 ;
        RECT 1146.880 110.540 1147.140 110.800 ;
        RECT 1146.420 110.200 1146.680 110.460 ;
        RECT 8.380 24.520 8.640 24.780 ;
        RECT 1145.960 24.520 1146.220 24.780 ;
      LAYER met2 ;
        RECT 1151.930 1700.000 1152.210 1704.000 ;
        RECT 1152.000 1676.870 1152.140 1700.000 ;
        RECT 1147.340 1676.550 1147.600 1676.870 ;
        RECT 1151.940 1676.550 1152.200 1676.870 ;
        RECT 1147.400 1628.445 1147.540 1676.550 ;
        RECT 1146.410 1628.075 1146.690 1628.445 ;
        RECT 1147.330 1628.075 1147.610 1628.445 ;
        RECT 1146.480 1580.650 1146.620 1628.075 ;
        RECT 1146.420 1580.330 1146.680 1580.650 ;
        RECT 1147.340 1580.330 1147.600 1580.650 ;
        RECT 1147.400 1579.970 1147.540 1580.330 ;
        RECT 1147.340 1579.650 1147.600 1579.970 ;
        RECT 1147.340 1510.290 1147.600 1510.610 ;
        RECT 1147.400 1463.690 1147.540 1510.290 ;
        RECT 1147.340 1463.370 1147.600 1463.690 ;
        RECT 1147.340 1400.810 1147.600 1401.130 ;
        RECT 1147.400 1376.990 1147.540 1400.810 ;
        RECT 1147.340 1376.670 1147.600 1376.990 ;
        RECT 1146.420 1352.530 1146.680 1352.850 ;
        RECT 1146.480 1318.170 1146.620 1352.530 ;
        RECT 1146.420 1317.850 1146.680 1318.170 ;
        RECT 1146.880 1317.510 1147.140 1317.830 ;
        RECT 1146.940 1304.230 1147.080 1317.510 ;
        RECT 1146.880 1303.910 1147.140 1304.230 ;
        RECT 1146.880 1268.890 1147.140 1269.210 ;
        RECT 1146.940 1221.950 1147.080 1268.890 ;
        RECT 1146.880 1221.630 1147.140 1221.950 ;
        RECT 1146.420 1220.950 1146.680 1221.270 ;
        RECT 1146.480 1200.725 1146.620 1220.950 ;
        RECT 1146.410 1200.355 1146.690 1200.725 ;
        RECT 1147.790 1200.355 1148.070 1200.725 ;
        RECT 1147.860 1152.590 1148.000 1200.355 ;
        RECT 1146.880 1152.270 1147.140 1152.590 ;
        RECT 1147.800 1152.270 1148.060 1152.590 ;
        RECT 1146.940 1125.390 1147.080 1152.270 ;
        RECT 1146.880 1125.070 1147.140 1125.390 ;
        RECT 1146.420 1124.390 1146.680 1124.710 ;
        RECT 1146.480 1104.165 1146.620 1124.390 ;
        RECT 1146.410 1103.795 1146.690 1104.165 ;
        RECT 1148.250 1103.795 1148.530 1104.165 ;
        RECT 1148.320 1027.810 1148.460 1103.795 ;
        RECT 1147.340 1027.490 1147.600 1027.810 ;
        RECT 1148.260 1027.490 1148.520 1027.810 ;
        RECT 1147.400 980.210 1147.540 1027.490 ;
        RECT 1146.420 979.890 1146.680 980.210 ;
        RECT 1147.340 979.890 1147.600 980.210 ;
        RECT 1146.480 961.850 1146.620 979.890 ;
        RECT 1146.420 961.530 1146.680 961.850 ;
        RECT 1146.880 917.670 1147.140 917.990 ;
        RECT 1146.940 883.990 1147.080 917.670 ;
        RECT 1146.880 883.670 1147.140 883.990 ;
        RECT 1146.880 882.650 1147.140 882.970 ;
        RECT 1146.940 834.770 1147.080 882.650 ;
        RECT 1146.480 834.630 1147.080 834.770 ;
        RECT 1146.480 787.090 1146.620 834.630 ;
        RECT 1146.420 786.770 1146.680 787.090 ;
        RECT 1146.880 786.430 1147.140 786.750 ;
        RECT 1146.940 772.810 1147.080 786.430 ;
        RECT 1146.880 772.490 1147.140 772.810 ;
        RECT 1147.800 772.490 1148.060 772.810 ;
        RECT 1147.860 724.725 1148.000 772.490 ;
        RECT 1146.410 724.355 1146.690 724.725 ;
        RECT 1147.790 724.355 1148.070 724.725 ;
        RECT 1146.480 690.190 1146.620 724.355 ;
        RECT 1146.420 689.870 1146.680 690.190 ;
        RECT 1146.880 689.530 1147.140 689.850 ;
        RECT 1146.940 676.250 1147.080 689.530 ;
        RECT 1146.880 675.930 1147.140 676.250 ;
        RECT 1147.800 675.930 1148.060 676.250 ;
        RECT 1147.860 628.165 1148.000 675.930 ;
        RECT 1146.410 627.795 1146.690 628.165 ;
        RECT 1147.790 627.795 1148.070 628.165 ;
        RECT 1146.480 593.630 1146.620 627.795 ;
        RECT 1146.420 593.310 1146.680 593.630 ;
        RECT 1146.880 592.970 1147.140 593.290 ;
        RECT 1146.940 579.690 1147.080 592.970 ;
        RECT 1146.880 579.370 1147.140 579.690 ;
        RECT 1146.420 531.430 1146.680 531.750 ;
        RECT 1146.480 497.070 1146.620 531.430 ;
        RECT 1146.420 496.750 1146.680 497.070 ;
        RECT 1146.880 496.410 1147.140 496.730 ;
        RECT 1146.940 483.130 1147.080 496.410 ;
        RECT 1146.880 482.810 1147.140 483.130 ;
        RECT 1146.420 434.870 1146.680 435.190 ;
        RECT 1146.480 400.510 1146.620 434.870 ;
        RECT 1146.420 400.190 1146.680 400.510 ;
        RECT 1146.880 399.510 1147.140 399.830 ;
        RECT 1146.940 386.230 1147.080 399.510 ;
        RECT 1146.880 385.910 1147.140 386.230 ;
        RECT 1146.420 337.970 1146.680 338.290 ;
        RECT 1146.480 304.370 1146.620 337.970 ;
        RECT 1146.480 304.230 1147.080 304.370 ;
        RECT 1146.940 290.010 1147.080 304.230 ;
        RECT 1146.420 289.690 1146.680 290.010 ;
        RECT 1146.880 289.690 1147.140 290.010 ;
        RECT 1146.480 289.330 1146.620 289.690 ;
        RECT 1146.420 289.010 1146.680 289.330 ;
        RECT 1146.880 241.410 1147.140 241.730 ;
        RECT 1146.940 207.730 1147.080 241.410 ;
        RECT 1146.880 207.410 1147.140 207.730 ;
        RECT 1145.960 193.130 1146.220 193.450 ;
        RECT 1146.020 162.170 1146.160 193.130 ;
        RECT 1145.960 161.850 1146.220 162.170 ;
        RECT 1146.880 138.050 1147.140 138.370 ;
        RECT 1146.940 110.830 1147.080 138.050 ;
        RECT 1146.880 110.510 1147.140 110.830 ;
        RECT 1146.420 110.170 1146.680 110.490 ;
        RECT 1146.480 72.490 1146.620 110.170 ;
        RECT 1146.020 72.350 1146.620 72.490 ;
        RECT 1146.020 24.810 1146.160 72.350 ;
        RECT 8.380 24.490 8.640 24.810 ;
        RECT 1145.960 24.490 1146.220 24.810 ;
        RECT 8.440 2.400 8.580 24.490 ;
        RECT 8.230 -4.800 8.790 2.400 ;
      LAYER via2 ;
        RECT 1146.410 1628.120 1146.690 1628.400 ;
        RECT 1147.330 1628.120 1147.610 1628.400 ;
        RECT 1146.410 1200.400 1146.690 1200.680 ;
        RECT 1147.790 1200.400 1148.070 1200.680 ;
        RECT 1146.410 1103.840 1146.690 1104.120 ;
        RECT 1148.250 1103.840 1148.530 1104.120 ;
        RECT 1146.410 724.400 1146.690 724.680 ;
        RECT 1147.790 724.400 1148.070 724.680 ;
        RECT 1146.410 627.840 1146.690 628.120 ;
        RECT 1147.790 627.840 1148.070 628.120 ;
      LAYER met3 ;
        RECT 1146.385 1628.410 1146.715 1628.425 ;
        RECT 1147.305 1628.410 1147.635 1628.425 ;
        RECT 1146.385 1628.110 1147.635 1628.410 ;
        RECT 1146.385 1628.095 1146.715 1628.110 ;
        RECT 1147.305 1628.095 1147.635 1628.110 ;
        RECT 1146.385 1200.690 1146.715 1200.705 ;
        RECT 1147.765 1200.690 1148.095 1200.705 ;
        RECT 1146.385 1200.390 1148.095 1200.690 ;
        RECT 1146.385 1200.375 1146.715 1200.390 ;
        RECT 1147.765 1200.375 1148.095 1200.390 ;
        RECT 1146.385 1104.130 1146.715 1104.145 ;
        RECT 1148.225 1104.130 1148.555 1104.145 ;
        RECT 1146.385 1103.830 1148.555 1104.130 ;
        RECT 1146.385 1103.815 1146.715 1103.830 ;
        RECT 1148.225 1103.815 1148.555 1103.830 ;
        RECT 1146.385 724.690 1146.715 724.705 ;
        RECT 1147.765 724.690 1148.095 724.705 ;
        RECT 1146.385 724.390 1148.095 724.690 ;
        RECT 1146.385 724.375 1146.715 724.390 ;
        RECT 1147.765 724.375 1148.095 724.390 ;
        RECT 1146.385 628.130 1146.715 628.145 ;
        RECT 1147.765 628.130 1148.095 628.145 ;
        RECT 1146.385 627.830 1148.095 628.130 ;
        RECT 1146.385 627.815 1146.715 627.830 ;
        RECT 1147.765 627.815 1148.095 627.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 0.300 ;
=======
      LAYER met1 ;
        RECT 14.330 24.380 14.650 24.440 ;
        RECT 1152.830 24.380 1153.150 24.440 ;
        RECT 14.330 24.240 1153.150 24.380 ;
        RECT 14.330 24.180 14.650 24.240 ;
        RECT 1152.830 24.180 1153.150 24.240 ;
      LAYER via ;
        RECT 14.360 24.180 14.620 24.440 ;
        RECT 1152.860 24.180 1153.120 24.440 ;
      LAYER met2 ;
        RECT 1153.310 1700.410 1153.590 1704.000 ;
        RECT 1152.920 1700.270 1153.590 1700.410 ;
        RECT 1152.920 24.470 1153.060 1700.270 ;
        RECT 1153.310 1700.000 1153.590 1700.270 ;
        RECT 14.360 24.150 14.620 24.470 ;
        RECT 1152.860 24.150 1153.120 24.470 ;
        RECT 14.420 2.400 14.560 24.150 ;
        RECT 14.210 -4.800 14.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 0.300 ;
=======
      LAYER met1 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 1160.190 25.060 1160.510 25.120 ;
        RECT 38.250 24.920 1160.510 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 1160.190 24.860 1160.510 24.920 ;
      LAYER via ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 1160.220 24.860 1160.480 25.120 ;
      LAYER met2 ;
        RECT 1159.750 1700.410 1160.030 1704.000 ;
        RECT 1159.750 1700.270 1160.420 1700.410 ;
        RECT 1159.750 1700.000 1160.030 1700.270 ;
        RECT 1160.280 25.150 1160.420 1700.270 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 1160.220 24.830 1160.480 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 38.130 -4.800 38.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 240.530 -4.800 241.090 0.300 ;
=======
        RECT 1214.490 1700.000 1214.770 1704.000 ;
        RECT 1214.560 24.325 1214.700 1700.000 ;
        RECT 240.670 23.955 240.950 24.325 ;
        RECT 1214.490 23.955 1214.770 24.325 ;
        RECT 240.740 2.400 240.880 23.955 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 240.670 24.000 240.950 24.280 ;
        RECT 1214.490 24.000 1214.770 24.280 ;
      LAYER met3 ;
        RECT 240.645 24.290 240.975 24.305 ;
        RECT 1214.465 24.290 1214.795 24.305 ;
        RECT 240.645 23.990 1214.795 24.290 ;
        RECT 240.645 23.975 240.975 23.990 ;
        RECT 1214.465 23.975 1214.795 23.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1214.930 1678.140 1215.250 1678.200 ;
        RECT 1218.150 1678.140 1218.470 1678.200 ;
        RECT 1214.930 1678.000 1218.470 1678.140 ;
        RECT 1214.930 1677.940 1215.250 1678.000 ;
        RECT 1218.150 1677.940 1218.470 1678.000 ;
      LAYER via ;
        RECT 1214.960 1677.940 1215.220 1678.200 ;
        RECT 1218.180 1677.940 1218.440 1678.200 ;
      LAYER met2 ;
        RECT 1219.550 1700.410 1219.830 1704.000 ;
        RECT 1218.240 1700.270 1219.830 1700.410 ;
        RECT 1218.240 1678.230 1218.380 1700.270 ;
        RECT 1219.550 1700.000 1219.830 1700.270 ;
        RECT 1214.960 1677.910 1215.220 1678.230 ;
        RECT 1218.180 1677.910 1218.440 1678.230 ;
        RECT 1215.020 25.005 1215.160 1677.910 ;
        RECT 258.150 24.635 258.430 25.005 ;
        RECT 1214.950 24.635 1215.230 25.005 ;
        RECT 258.220 2.400 258.360 24.635 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 258.150 24.680 258.430 24.960 ;
        RECT 1214.950 24.680 1215.230 24.960 ;
      LAYER met3 ;
        RECT 258.125 24.970 258.455 24.985 ;
        RECT 1214.925 24.970 1215.255 24.985 ;
        RECT 258.125 24.670 1215.255 24.970 ;
        RECT 258.125 24.655 258.455 24.670 ;
        RECT 1214.925 24.655 1215.255 24.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 0.300 ;
=======
      LAYER met1 ;
        RECT 1221.830 1695.480 1222.150 1695.540 ;
        RECT 1224.130 1695.480 1224.450 1695.540 ;
        RECT 1221.830 1695.340 1224.450 1695.480 ;
        RECT 1221.830 1695.280 1222.150 1695.340 ;
        RECT 1224.130 1695.280 1224.450 1695.340 ;
        RECT 276.070 25.400 276.390 25.460 ;
        RECT 1221.830 25.400 1222.150 25.460 ;
        RECT 276.070 25.260 1222.150 25.400 ;
        RECT 276.070 25.200 276.390 25.260 ;
        RECT 1221.830 25.200 1222.150 25.260 ;
      LAYER via ;
        RECT 1221.860 1695.280 1222.120 1695.540 ;
        RECT 1224.160 1695.280 1224.420 1695.540 ;
        RECT 276.100 25.200 276.360 25.460 ;
        RECT 1221.860 25.200 1222.120 25.460 ;
      LAYER met2 ;
        RECT 1224.150 1700.000 1224.430 1704.000 ;
        RECT 1224.220 1695.570 1224.360 1700.000 ;
        RECT 1221.860 1695.250 1222.120 1695.570 ;
        RECT 1224.160 1695.250 1224.420 1695.570 ;
        RECT 1221.920 25.490 1222.060 1695.250 ;
        RECT 276.100 25.170 276.360 25.490 ;
        RECT 1221.860 25.170 1222.120 25.490 ;
        RECT 276.160 2.400 276.300 25.170 ;
        RECT 275.950 -4.800 276.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 293.890 -4.800 294.450 0.300 ;
=======
        RECT 1229.210 1700.410 1229.490 1704.000 ;
        RECT 1229.210 1700.270 1229.880 1700.410 ;
        RECT 1229.210 1700.000 1229.490 1700.270 ;
        RECT 1229.740 31.125 1229.880 1700.270 ;
        RECT 294.030 30.755 294.310 31.125 ;
        RECT 1229.670 30.755 1229.950 31.125 ;
        RECT 294.100 2.400 294.240 30.755 ;
        RECT 293.890 -4.800 294.450 2.400 ;
      LAYER via2 ;
        RECT 294.030 30.800 294.310 31.080 ;
        RECT 1229.670 30.800 1229.950 31.080 ;
      LAYER met3 ;
        RECT 294.005 31.090 294.335 31.105 ;
        RECT 1229.645 31.090 1229.975 31.105 ;
        RECT 294.005 30.790 1229.975 31.090 ;
        RECT 294.005 30.775 294.335 30.790 ;
        RECT 1229.645 30.775 1229.975 30.790 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1228.730 1678.140 1229.050 1678.200 ;
        RECT 1232.870 1678.140 1233.190 1678.200 ;
        RECT 1228.730 1678.000 1233.190 1678.140 ;
        RECT 1228.730 1677.940 1229.050 1678.000 ;
        RECT 1232.870 1677.940 1233.190 1678.000 ;
      LAYER via ;
        RECT 1228.760 1677.940 1229.020 1678.200 ;
        RECT 1232.900 1677.940 1233.160 1678.200 ;
      LAYER met2 ;
        RECT 1233.810 1700.410 1234.090 1704.000 ;
        RECT 1232.960 1700.270 1234.090 1700.410 ;
        RECT 1232.960 1678.230 1233.100 1700.270 ;
        RECT 1233.810 1700.000 1234.090 1700.270 ;
        RECT 1228.760 1677.910 1229.020 1678.230 ;
        RECT 1232.900 1677.910 1233.160 1678.230 ;
        RECT 1228.820 31.805 1228.960 1677.910 ;
        RECT 311.970 31.435 312.250 31.805 ;
        RECT 1228.750 31.435 1229.030 31.805 ;
        RECT 312.040 2.400 312.180 31.435 ;
        RECT 311.830 -4.800 312.390 2.400 ;
      LAYER via2 ;
        RECT 311.970 31.480 312.250 31.760 ;
        RECT 1228.750 31.480 1229.030 31.760 ;
      LAYER met3 ;
        RECT 311.945 31.770 312.275 31.785 ;
        RECT 1228.725 31.770 1229.055 31.785 ;
        RECT 311.945 31.470 1229.055 31.770 ;
        RECT 311.945 31.455 312.275 31.470 ;
        RECT 1228.725 31.455 1229.055 31.470 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 329.770 -4.800 330.330 0.300 ;
=======
        RECT 1238.870 1700.410 1239.150 1704.000 ;
        RECT 1238.020 1700.270 1239.150 1700.410 ;
        RECT 1238.020 1678.650 1238.160 1700.270 ;
        RECT 1238.870 1700.000 1239.150 1700.270 ;
        RECT 1236.640 1678.510 1238.160 1678.650 ;
        RECT 1236.640 32.485 1236.780 1678.510 ;
        RECT 329.910 32.115 330.190 32.485 ;
        RECT 1236.570 32.115 1236.850 32.485 ;
        RECT 329.980 2.400 330.120 32.115 ;
        RECT 329.770 -4.800 330.330 2.400 ;
      LAYER via2 ;
        RECT 329.910 32.160 330.190 32.440 ;
        RECT 1236.570 32.160 1236.850 32.440 ;
      LAYER met3 ;
        RECT 329.885 32.450 330.215 32.465 ;
        RECT 1236.545 32.450 1236.875 32.465 ;
        RECT 329.885 32.150 1236.875 32.450 ;
        RECT 329.885 32.135 330.215 32.150 ;
        RECT 1236.545 32.135 1236.875 32.150 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 0.300 ;
=======
      LAYER met1 ;
        RECT 347.370 37.980 347.690 38.040 ;
        RECT 1242.530 37.980 1242.850 38.040 ;
        RECT 347.370 37.840 1242.850 37.980 ;
        RECT 347.370 37.780 347.690 37.840 ;
        RECT 1242.530 37.780 1242.850 37.840 ;
      LAYER via ;
        RECT 347.400 37.780 347.660 38.040 ;
        RECT 1242.560 37.780 1242.820 38.040 ;
      LAYER met2 ;
        RECT 1243.470 1700.410 1243.750 1704.000 ;
        RECT 1242.620 1700.270 1243.750 1700.410 ;
        RECT 1242.620 38.070 1242.760 1700.270 ;
        RECT 1243.470 1700.000 1243.750 1700.270 ;
        RECT 347.400 37.750 347.660 38.070 ;
        RECT 1242.560 37.750 1242.820 38.070 ;
        RECT 347.460 2.400 347.600 37.750 ;
        RECT 347.250 -4.800 347.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1242.990 1678.140 1243.310 1678.200 ;
        RECT 1247.130 1678.140 1247.450 1678.200 ;
        RECT 1242.990 1678.000 1247.450 1678.140 ;
        RECT 1242.990 1677.940 1243.310 1678.000 ;
        RECT 1247.130 1677.940 1247.450 1678.000 ;
        RECT 364.850 38.320 365.170 38.380 ;
        RECT 1242.990 38.320 1243.310 38.380 ;
        RECT 364.850 38.180 1243.310 38.320 ;
        RECT 364.850 38.120 365.170 38.180 ;
        RECT 1242.990 38.120 1243.310 38.180 ;
      LAYER via ;
        RECT 1243.020 1677.940 1243.280 1678.200 ;
        RECT 1247.160 1677.940 1247.420 1678.200 ;
        RECT 364.880 38.120 365.140 38.380 ;
        RECT 1243.020 38.120 1243.280 38.380 ;
      LAYER met2 ;
        RECT 1248.530 1700.410 1248.810 1704.000 ;
        RECT 1247.220 1700.270 1248.810 1700.410 ;
        RECT 1247.220 1678.230 1247.360 1700.270 ;
        RECT 1248.530 1700.000 1248.810 1700.270 ;
        RECT 1243.020 1677.910 1243.280 1678.230 ;
        RECT 1247.160 1677.910 1247.420 1678.230 ;
        RECT 1243.080 38.410 1243.220 1677.910 ;
        RECT 364.880 38.090 365.140 38.410 ;
        RECT 1243.020 38.090 1243.280 38.410 ;
        RECT 364.940 7.890 365.080 38.090 ;
        RECT 364.940 7.750 365.540 7.890 ;
        RECT 365.400 2.400 365.540 7.750 ;
        RECT 365.190 -4.800 365.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1249.430 1678.140 1249.750 1678.200 ;
        RECT 1251.730 1678.140 1252.050 1678.200 ;
        RECT 1249.430 1678.000 1252.050 1678.140 ;
        RECT 1249.430 1677.940 1249.750 1678.000 ;
        RECT 1251.730 1677.940 1252.050 1678.000 ;
        RECT 1249.430 1435.520 1249.750 1435.780 ;
        RECT 1249.520 1435.100 1249.660 1435.520 ;
        RECT 1249.430 1434.840 1249.750 1435.100 ;
        RECT 383.250 38.660 383.570 38.720 ;
        RECT 1249.430 38.660 1249.750 38.720 ;
        RECT 383.250 38.520 1249.750 38.660 ;
        RECT 383.250 38.460 383.570 38.520 ;
        RECT 1249.430 38.460 1249.750 38.520 ;
      LAYER via ;
        RECT 1249.460 1677.940 1249.720 1678.200 ;
        RECT 1251.760 1677.940 1252.020 1678.200 ;
        RECT 1249.460 1435.520 1249.720 1435.780 ;
        RECT 1249.460 1434.840 1249.720 1435.100 ;
        RECT 383.280 38.460 383.540 38.720 ;
        RECT 1249.460 38.460 1249.720 38.720 ;
      LAYER met2 ;
        RECT 1253.130 1700.410 1253.410 1704.000 ;
        RECT 1251.820 1700.270 1253.410 1700.410 ;
        RECT 1251.820 1678.230 1251.960 1700.270 ;
        RECT 1253.130 1700.000 1253.410 1700.270 ;
        RECT 1249.460 1677.910 1249.720 1678.230 ;
        RECT 1251.760 1677.910 1252.020 1678.230 ;
        RECT 1249.520 1435.810 1249.660 1677.910 ;
        RECT 1249.460 1435.490 1249.720 1435.810 ;
        RECT 1249.460 1434.810 1249.720 1435.130 ;
        RECT 1249.520 38.750 1249.660 1434.810 ;
        RECT 383.280 38.430 383.540 38.750 ;
        RECT 1249.460 38.430 1249.720 38.750 ;
        RECT 383.340 2.400 383.480 38.430 ;
        RECT 383.130 -4.800 383.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 0.300 ;
=======
      LAYER li1 ;
        RECT 1257.785 1594.005 1257.955 1680.535 ;
        RECT 1257.785 386.325 1257.955 434.775 ;
      LAYER mcon ;
        RECT 1257.785 1680.365 1257.955 1680.535 ;
        RECT 1257.785 434.605 1257.955 434.775 ;
      LAYER met1 ;
        RECT 1257.710 1680.520 1258.030 1680.580 ;
        RECT 1257.515 1680.380 1258.030 1680.520 ;
        RECT 1257.710 1680.320 1258.030 1680.380 ;
        RECT 1257.710 1594.160 1258.030 1594.220 ;
        RECT 1257.515 1594.020 1258.030 1594.160 ;
        RECT 1257.710 1593.960 1258.030 1594.020 ;
        RECT 1258.170 1546.220 1258.490 1546.280 ;
        RECT 1257.800 1546.080 1258.490 1546.220 ;
        RECT 1257.800 1545.940 1257.940 1546.080 ;
        RECT 1258.170 1546.020 1258.490 1546.080 ;
        RECT 1257.710 1545.680 1258.030 1545.940 ;
        RECT 1257.710 966.180 1258.030 966.240 ;
        RECT 1258.630 966.180 1258.950 966.240 ;
        RECT 1257.710 966.040 1258.950 966.180 ;
        RECT 1257.710 965.980 1258.030 966.040 ;
        RECT 1258.630 965.980 1258.950 966.040 ;
        RECT 1257.710 434.760 1258.030 434.820 ;
        RECT 1257.515 434.620 1258.030 434.760 ;
        RECT 1257.710 434.560 1258.030 434.620 ;
        RECT 1257.710 386.480 1258.030 386.540 ;
        RECT 1257.515 386.340 1258.030 386.480 ;
        RECT 1257.710 386.280 1258.030 386.340 ;
      LAYER via ;
        RECT 1257.740 1680.320 1258.000 1680.580 ;
        RECT 1257.740 1593.960 1258.000 1594.220 ;
        RECT 1258.200 1546.020 1258.460 1546.280 ;
        RECT 1257.740 1545.680 1258.000 1545.940 ;
        RECT 1257.740 965.980 1258.000 966.240 ;
        RECT 1258.660 965.980 1258.920 966.240 ;
        RECT 1257.740 434.560 1258.000 434.820 ;
        RECT 1257.740 386.280 1258.000 386.540 ;
      LAYER met2 ;
        RECT 1257.730 1700.000 1258.010 1704.000 ;
        RECT 1257.800 1680.610 1257.940 1700.000 ;
        RECT 1257.740 1680.290 1258.000 1680.610 ;
        RECT 1257.740 1593.930 1258.000 1594.250 ;
        RECT 1257.800 1593.650 1257.940 1593.930 ;
        RECT 1257.800 1593.510 1258.400 1593.650 ;
        RECT 1258.260 1546.310 1258.400 1593.510 ;
        RECT 1258.200 1545.990 1258.460 1546.310 ;
        RECT 1257.740 1545.650 1258.000 1545.970 ;
        RECT 1257.800 1014.405 1257.940 1545.650 ;
        RECT 1257.730 1014.035 1258.010 1014.405 ;
        RECT 1258.650 1014.035 1258.930 1014.405 ;
        RECT 1258.720 966.270 1258.860 1014.035 ;
        RECT 1257.740 965.950 1258.000 966.270 ;
        RECT 1258.660 965.950 1258.920 966.270 ;
        RECT 1257.800 434.850 1257.940 965.950 ;
        RECT 1257.740 434.530 1258.000 434.850 ;
        RECT 1257.740 386.250 1258.000 386.570 ;
        RECT 1257.800 46.765 1257.940 386.250 ;
        RECT 401.210 46.395 401.490 46.765 ;
        RECT 1257.730 46.395 1258.010 46.765 ;
        RECT 401.280 2.400 401.420 46.395 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 1257.730 1014.080 1258.010 1014.360 ;
        RECT 1258.650 1014.080 1258.930 1014.360 ;
        RECT 401.210 46.440 401.490 46.720 ;
        RECT 1257.730 46.440 1258.010 46.720 ;
      LAYER met3 ;
        RECT 1257.705 1014.370 1258.035 1014.385 ;
        RECT 1258.625 1014.370 1258.955 1014.385 ;
        RECT 1257.705 1014.070 1258.955 1014.370 ;
        RECT 1257.705 1014.055 1258.035 1014.070 ;
        RECT 1258.625 1014.055 1258.955 1014.070 ;
        RECT 401.185 46.730 401.515 46.745 ;
        RECT 1257.705 46.730 1258.035 46.745 ;
        RECT 401.185 46.430 1258.035 46.730 ;
        RECT 401.185 46.415 401.515 46.430 ;
        RECT 1257.705 46.415 1258.035 46.430 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 62.050 -4.800 62.610 0.300 ;
=======
        RECT 1166.190 1700.410 1166.470 1704.000 ;
        RECT 1166.190 1700.270 1167.320 1700.410 ;
        RECT 1166.190 1700.000 1166.470 1700.270 ;
        RECT 1167.180 38.605 1167.320 1700.270 ;
        RECT 62.190 38.235 62.470 38.605 ;
        RECT 1167.110 38.235 1167.390 38.605 ;
        RECT 62.260 2.400 62.400 38.235 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 62.190 38.280 62.470 38.560 ;
        RECT 1167.110 38.280 1167.390 38.560 ;
      LAYER met3 ;
        RECT 62.165 38.570 62.495 38.585 ;
        RECT 1167.085 38.570 1167.415 38.585 ;
        RECT 62.165 38.270 1167.415 38.570 ;
        RECT 62.165 38.255 62.495 38.270 ;
        RECT 1167.085 38.255 1167.415 38.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 419.010 -4.800 419.570 0.300 ;
=======
        RECT 1262.790 1700.000 1263.070 1704.000 ;
        RECT 1262.860 47.445 1263.000 1700.000 ;
        RECT 419.150 47.075 419.430 47.445 ;
        RECT 1262.790 47.075 1263.070 47.445 ;
        RECT 419.220 2.400 419.360 47.075 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 419.150 47.120 419.430 47.400 ;
        RECT 1262.790 47.120 1263.070 47.400 ;
      LAYER met3 ;
        RECT 419.125 47.410 419.455 47.425 ;
        RECT 1262.765 47.410 1263.095 47.425 ;
        RECT 419.125 47.110 1263.095 47.410 ;
        RECT 419.125 47.095 419.455 47.110 ;
        RECT 1262.765 47.095 1263.095 47.110 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1263.230 1665.560 1263.550 1665.620 ;
        RECT 1266.450 1665.560 1266.770 1665.620 ;
        RECT 1263.230 1665.420 1266.770 1665.560 ;
        RECT 1263.230 1665.360 1263.550 1665.420 ;
        RECT 1266.450 1665.360 1266.770 1665.420 ;
      LAYER via ;
        RECT 1263.260 1665.360 1263.520 1665.620 ;
        RECT 1266.480 1665.360 1266.740 1665.620 ;
      LAYER met2 ;
        RECT 1267.390 1700.410 1267.670 1704.000 ;
        RECT 1266.540 1700.270 1267.670 1700.410 ;
        RECT 1266.540 1665.650 1266.680 1700.270 ;
        RECT 1267.390 1700.000 1267.670 1700.270 ;
        RECT 1263.260 1665.330 1263.520 1665.650 ;
        RECT 1266.480 1665.330 1266.740 1665.650 ;
        RECT 1263.320 48.125 1263.460 1665.330 ;
        RECT 436.630 47.755 436.910 48.125 ;
        RECT 1263.250 47.755 1263.530 48.125 ;
        RECT 436.700 2.400 436.840 47.755 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 436.630 47.800 436.910 48.080 ;
        RECT 1263.250 47.800 1263.530 48.080 ;
      LAYER met3 ;
        RECT 436.605 48.090 436.935 48.105 ;
        RECT 1263.225 48.090 1263.555 48.105 ;
        RECT 436.605 47.790 1263.555 48.090 ;
        RECT 436.605 47.775 436.935 47.790 ;
        RECT 1263.225 47.775 1263.555 47.790 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 0.300 ;
=======
      LAYER met1 ;
        RECT 454.550 44.780 454.870 44.840 ;
        RECT 1270.130 44.780 1270.450 44.840 ;
        RECT 454.550 44.640 1270.450 44.780 ;
        RECT 454.550 44.580 454.870 44.640 ;
        RECT 1270.130 44.580 1270.450 44.640 ;
      LAYER via ;
        RECT 454.580 44.580 454.840 44.840 ;
        RECT 1270.160 44.580 1270.420 44.840 ;
      LAYER met2 ;
        RECT 1272.450 1700.410 1272.730 1704.000 ;
        RECT 1271.140 1700.270 1272.730 1700.410 ;
        RECT 1271.140 1678.140 1271.280 1700.270 ;
        RECT 1272.450 1700.000 1272.730 1700.270 ;
        RECT 1270.220 1678.000 1271.280 1678.140 ;
        RECT 1270.220 44.870 1270.360 1678.000 ;
        RECT 454.580 44.550 454.840 44.870 ;
        RECT 1270.160 44.550 1270.420 44.870 ;
        RECT 454.640 2.400 454.780 44.550 ;
        RECT 454.430 -4.800 454.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 0.300 ;
=======
      LAYER met1 ;
        RECT 472.490 45.120 472.810 45.180 ;
        RECT 1277.030 45.120 1277.350 45.180 ;
        RECT 472.490 44.980 1277.350 45.120 ;
        RECT 472.490 44.920 472.810 44.980 ;
        RECT 1277.030 44.920 1277.350 44.980 ;
      LAYER via ;
        RECT 472.520 44.920 472.780 45.180 ;
        RECT 1277.060 44.920 1277.320 45.180 ;
      LAYER met2 ;
        RECT 1277.050 1700.000 1277.330 1704.000 ;
        RECT 1277.120 45.210 1277.260 1700.000 ;
        RECT 472.520 44.890 472.780 45.210 ;
        RECT 1277.060 44.890 1277.320 45.210 ;
        RECT 472.580 2.400 472.720 44.890 ;
        RECT 472.370 -4.800 472.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 0.300 ;
=======
      LAYER li1 ;
        RECT 1278.485 1490.645 1278.655 1538.755 ;
        RECT 1278.025 1401.225 1278.195 1448.995 ;
        RECT 1278.485 45.305 1278.655 131.155 ;
      LAYER mcon ;
        RECT 1278.485 1538.585 1278.655 1538.755 ;
        RECT 1278.025 1448.825 1278.195 1448.995 ;
        RECT 1278.485 130.985 1278.655 131.155 ;
      LAYER met1 ;
        RECT 1278.410 1539.420 1278.730 1539.480 ;
        RECT 1279.330 1539.420 1279.650 1539.480 ;
        RECT 1278.410 1539.280 1279.650 1539.420 ;
        RECT 1278.410 1539.220 1278.730 1539.280 ;
        RECT 1279.330 1539.220 1279.650 1539.280 ;
        RECT 1278.425 1538.740 1278.715 1538.785 ;
        RECT 1279.330 1538.740 1279.650 1538.800 ;
        RECT 1278.425 1538.600 1279.650 1538.740 ;
        RECT 1278.425 1538.555 1278.715 1538.600 ;
        RECT 1279.330 1538.540 1279.650 1538.600 ;
        RECT 1278.410 1490.800 1278.730 1490.860 ;
        RECT 1278.215 1490.660 1278.730 1490.800 ;
        RECT 1278.410 1490.600 1278.730 1490.660 ;
        RECT 1277.965 1448.980 1278.255 1449.025 ;
        RECT 1278.410 1448.980 1278.730 1449.040 ;
        RECT 1277.965 1448.840 1278.730 1448.980 ;
        RECT 1277.965 1448.795 1278.255 1448.840 ;
        RECT 1278.410 1448.780 1278.730 1448.840 ;
        RECT 1277.950 1401.380 1278.270 1401.440 ;
        RECT 1277.755 1401.240 1278.270 1401.380 ;
        RECT 1277.950 1401.180 1278.270 1401.240 ;
        RECT 1277.950 1269.600 1278.270 1269.860 ;
        RECT 1278.040 1269.120 1278.180 1269.600 ;
        RECT 1278.410 1269.120 1278.730 1269.180 ;
        RECT 1278.040 1268.980 1278.730 1269.120 ;
        RECT 1278.410 1268.920 1278.730 1268.980 ;
        RECT 1278.410 1207.920 1278.730 1207.980 ;
        RECT 1278.040 1207.780 1278.730 1207.920 ;
        RECT 1278.040 1207.640 1278.180 1207.780 ;
        RECT 1278.410 1207.720 1278.730 1207.780 ;
        RECT 1277.950 1207.380 1278.270 1207.640 ;
        RECT 1278.410 959.040 1278.730 959.100 ;
        RECT 1279.330 959.040 1279.650 959.100 ;
        RECT 1278.410 958.900 1279.650 959.040 ;
        RECT 1278.410 958.840 1278.730 958.900 ;
        RECT 1279.330 958.840 1279.650 958.900 ;
        RECT 1277.950 910.760 1278.270 910.820 ;
        RECT 1278.870 910.760 1279.190 910.820 ;
        RECT 1277.950 910.620 1279.190 910.760 ;
        RECT 1277.950 910.560 1278.270 910.620 ;
        RECT 1278.870 910.560 1279.190 910.620 ;
        RECT 1277.950 759.120 1278.270 759.180 ;
        RECT 1278.410 759.120 1278.730 759.180 ;
        RECT 1277.950 758.980 1278.730 759.120 ;
        RECT 1277.950 758.920 1278.270 758.980 ;
        RECT 1278.410 758.920 1278.730 758.980 ;
        RECT 1277.950 572.940 1278.270 573.200 ;
        RECT 1278.040 572.800 1278.180 572.940 ;
        RECT 1278.410 572.800 1278.730 572.860 ;
        RECT 1278.040 572.660 1278.730 572.800 ;
        RECT 1278.410 572.600 1278.730 572.660 ;
        RECT 1277.950 476.240 1278.270 476.300 ;
        RECT 1278.410 476.240 1278.730 476.300 ;
        RECT 1277.950 476.100 1278.730 476.240 ;
        RECT 1277.950 476.040 1278.270 476.100 ;
        RECT 1278.410 476.040 1278.730 476.100 ;
        RECT 1277.950 434.560 1278.270 434.820 ;
        RECT 1278.040 434.420 1278.180 434.560 ;
        RECT 1278.410 434.420 1278.730 434.480 ;
        RECT 1278.040 434.280 1278.730 434.420 ;
        RECT 1278.410 434.220 1278.730 434.280 ;
        RECT 1277.950 186.560 1278.270 186.620 ;
        RECT 1278.410 186.560 1278.730 186.620 ;
        RECT 1277.950 186.420 1278.730 186.560 ;
        RECT 1277.950 186.360 1278.270 186.420 ;
        RECT 1278.410 186.360 1278.730 186.420 ;
        RECT 1277.950 137.740 1278.270 138.000 ;
        RECT 1278.040 137.600 1278.180 137.740 ;
        RECT 1278.410 137.600 1278.730 137.660 ;
        RECT 1278.040 137.460 1278.730 137.600 ;
        RECT 1278.410 137.400 1278.730 137.460 ;
        RECT 1278.410 131.140 1278.730 131.200 ;
        RECT 1278.215 131.000 1278.730 131.140 ;
        RECT 1278.410 130.940 1278.730 131.000 ;
        RECT 490.430 45.460 490.750 45.520 ;
        RECT 1278.425 45.460 1278.715 45.505 ;
        RECT 490.430 45.320 1278.715 45.460 ;
        RECT 490.430 45.260 490.750 45.320 ;
        RECT 1278.425 45.275 1278.715 45.320 ;
      LAYER via ;
        RECT 1278.440 1539.220 1278.700 1539.480 ;
        RECT 1279.360 1539.220 1279.620 1539.480 ;
        RECT 1279.360 1538.540 1279.620 1538.800 ;
        RECT 1278.440 1490.600 1278.700 1490.860 ;
        RECT 1278.440 1448.780 1278.700 1449.040 ;
        RECT 1277.980 1401.180 1278.240 1401.440 ;
        RECT 1277.980 1269.600 1278.240 1269.860 ;
        RECT 1278.440 1268.920 1278.700 1269.180 ;
        RECT 1278.440 1207.720 1278.700 1207.980 ;
        RECT 1277.980 1207.380 1278.240 1207.640 ;
        RECT 1278.440 958.840 1278.700 959.100 ;
        RECT 1279.360 958.840 1279.620 959.100 ;
        RECT 1277.980 910.560 1278.240 910.820 ;
        RECT 1278.900 910.560 1279.160 910.820 ;
        RECT 1277.980 758.920 1278.240 759.180 ;
        RECT 1278.440 758.920 1278.700 759.180 ;
        RECT 1277.980 572.940 1278.240 573.200 ;
        RECT 1278.440 572.600 1278.700 572.860 ;
        RECT 1277.980 476.040 1278.240 476.300 ;
        RECT 1278.440 476.040 1278.700 476.300 ;
        RECT 1277.980 434.560 1278.240 434.820 ;
        RECT 1278.440 434.220 1278.700 434.480 ;
        RECT 1277.980 186.360 1278.240 186.620 ;
        RECT 1278.440 186.360 1278.700 186.620 ;
        RECT 1277.980 137.740 1278.240 138.000 ;
        RECT 1278.440 137.400 1278.700 137.660 ;
        RECT 1278.440 130.940 1278.700 131.200 ;
        RECT 490.460 45.260 490.720 45.520 ;
      LAYER met2 ;
        RECT 1282.110 1700.410 1282.390 1704.000 ;
        RECT 1281.260 1700.270 1282.390 1700.410 ;
        RECT 1281.260 1656.210 1281.400 1700.270 ;
        RECT 1282.110 1700.000 1282.390 1700.270 ;
        RECT 1278.500 1656.070 1281.400 1656.210 ;
        RECT 1278.500 1605.210 1278.640 1656.070 ;
        RECT 1278.040 1605.070 1278.640 1605.210 ;
        RECT 1278.040 1603.850 1278.180 1605.070 ;
        RECT 1278.040 1603.710 1278.640 1603.850 ;
        RECT 1278.500 1539.510 1278.640 1603.710 ;
        RECT 1278.440 1539.190 1278.700 1539.510 ;
        RECT 1279.360 1539.190 1279.620 1539.510 ;
        RECT 1279.420 1538.830 1279.560 1539.190 ;
        RECT 1279.360 1538.510 1279.620 1538.830 ;
        RECT 1278.440 1490.570 1278.700 1490.890 ;
        RECT 1278.500 1449.070 1278.640 1490.570 ;
        RECT 1278.440 1448.750 1278.700 1449.070 ;
        RECT 1277.980 1401.150 1278.240 1401.470 ;
        RECT 1278.040 1269.890 1278.180 1401.150 ;
        RECT 1277.980 1269.570 1278.240 1269.890 ;
        RECT 1278.440 1268.890 1278.700 1269.210 ;
        RECT 1278.500 1208.010 1278.640 1268.890 ;
        RECT 1278.440 1207.690 1278.700 1208.010 ;
        RECT 1277.980 1207.350 1278.240 1207.670 ;
        RECT 1278.040 1200.725 1278.180 1207.350 ;
        RECT 1277.970 1200.355 1278.250 1200.725 ;
        RECT 1278.890 1200.355 1279.170 1200.725 ;
        RECT 1278.960 1176.130 1279.100 1200.355 ;
        RECT 1278.500 1175.990 1279.100 1176.130 ;
        RECT 1278.500 1056.565 1278.640 1175.990 ;
        RECT 1278.430 1056.195 1278.710 1056.565 ;
        RECT 1278.430 1055.515 1278.710 1055.885 ;
        RECT 1278.500 959.130 1278.640 1055.515 ;
        RECT 1278.440 958.810 1278.700 959.130 ;
        RECT 1279.360 958.810 1279.620 959.130 ;
        RECT 1279.420 911.045 1279.560 958.810 ;
        RECT 1277.970 910.675 1278.250 911.045 ;
        RECT 1277.980 910.530 1278.240 910.675 ;
        RECT 1278.900 910.530 1279.160 910.850 ;
        RECT 1279.350 910.675 1279.630 911.045 ;
        RECT 1278.960 821.285 1279.100 910.530 ;
        RECT 1277.970 820.915 1278.250 821.285 ;
        RECT 1278.890 820.915 1279.170 821.285 ;
        RECT 1278.040 759.210 1278.180 820.915 ;
        RECT 1277.980 758.890 1278.240 759.210 ;
        RECT 1278.440 758.890 1278.700 759.210 ;
        RECT 1278.500 758.610 1278.640 758.890 ;
        RECT 1278.500 758.470 1279.100 758.610 ;
        RECT 1278.960 688.570 1279.100 758.470 ;
        RECT 1278.500 688.430 1279.100 688.570 ;
        RECT 1278.500 628.845 1278.640 688.430 ;
        RECT 1278.430 628.475 1278.710 628.845 ;
        RECT 1277.970 627.795 1278.250 628.165 ;
        RECT 1278.040 573.230 1278.180 627.795 ;
        RECT 1277.980 572.910 1278.240 573.230 ;
        RECT 1278.440 572.570 1278.700 572.890 ;
        RECT 1278.500 476.330 1278.640 572.570 ;
        RECT 1277.980 476.010 1278.240 476.330 ;
        RECT 1278.440 476.010 1278.700 476.330 ;
        RECT 1278.040 434.850 1278.180 476.010 ;
        RECT 1277.980 434.530 1278.240 434.850 ;
        RECT 1278.440 434.190 1278.700 434.510 ;
        RECT 1278.500 338.370 1278.640 434.190 ;
        RECT 1278.040 338.230 1278.640 338.370 ;
        RECT 1278.040 186.650 1278.180 338.230 ;
        RECT 1277.980 186.330 1278.240 186.650 ;
        RECT 1278.440 186.330 1278.700 186.650 ;
        RECT 1278.500 162.250 1278.640 186.330 ;
        RECT 1278.040 162.110 1278.640 162.250 ;
        RECT 1278.040 138.030 1278.180 162.110 ;
        RECT 1277.980 137.710 1278.240 138.030 ;
        RECT 1278.440 137.370 1278.700 137.690 ;
        RECT 1278.500 131.230 1278.640 137.370 ;
        RECT 1278.440 130.910 1278.700 131.230 ;
        RECT 490.460 45.230 490.720 45.550 ;
        RECT 490.520 2.400 490.660 45.230 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 1277.970 1200.400 1278.250 1200.680 ;
        RECT 1278.890 1200.400 1279.170 1200.680 ;
        RECT 1278.430 1056.240 1278.710 1056.520 ;
        RECT 1278.430 1055.560 1278.710 1055.840 ;
        RECT 1277.970 910.720 1278.250 911.000 ;
        RECT 1279.350 910.720 1279.630 911.000 ;
        RECT 1277.970 820.960 1278.250 821.240 ;
        RECT 1278.890 820.960 1279.170 821.240 ;
        RECT 1278.430 628.520 1278.710 628.800 ;
        RECT 1277.970 627.840 1278.250 628.120 ;
      LAYER met3 ;
        RECT 1277.945 1200.690 1278.275 1200.705 ;
        RECT 1278.865 1200.690 1279.195 1200.705 ;
        RECT 1277.945 1200.390 1279.195 1200.690 ;
        RECT 1277.945 1200.375 1278.275 1200.390 ;
        RECT 1278.865 1200.375 1279.195 1200.390 ;
        RECT 1278.405 1056.530 1278.735 1056.545 ;
        RECT 1278.190 1056.215 1278.735 1056.530 ;
        RECT 1278.190 1055.865 1278.490 1056.215 ;
        RECT 1278.190 1055.550 1278.735 1055.865 ;
        RECT 1278.405 1055.535 1278.735 1055.550 ;
        RECT 1277.945 911.010 1278.275 911.025 ;
        RECT 1279.325 911.010 1279.655 911.025 ;
        RECT 1277.945 910.710 1279.655 911.010 ;
        RECT 1277.945 910.695 1278.275 910.710 ;
        RECT 1279.325 910.695 1279.655 910.710 ;
        RECT 1277.945 821.250 1278.275 821.265 ;
        RECT 1278.865 821.250 1279.195 821.265 ;
        RECT 1277.945 820.950 1279.195 821.250 ;
        RECT 1277.945 820.935 1278.275 820.950 ;
        RECT 1278.865 820.935 1279.195 820.950 ;
        RECT 1278.405 628.810 1278.735 628.825 ;
        RECT 1278.190 628.495 1278.735 628.810 ;
        RECT 1278.190 628.145 1278.490 628.495 ;
        RECT 1277.945 627.830 1278.490 628.145 ;
        RECT 1277.945 627.815 1278.275 627.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1283.930 1678.140 1284.250 1678.200 ;
        RECT 1285.770 1678.140 1286.090 1678.200 ;
        RECT 1283.930 1678.000 1286.090 1678.140 ;
        RECT 1283.930 1677.940 1284.250 1678.000 ;
        RECT 1285.770 1677.940 1286.090 1678.000 ;
        RECT 507.910 45.800 508.230 45.860 ;
        RECT 1283.930 45.800 1284.250 45.860 ;
        RECT 507.910 45.660 1284.250 45.800 ;
        RECT 507.910 45.600 508.230 45.660 ;
        RECT 1283.930 45.600 1284.250 45.660 ;
      LAYER via ;
        RECT 1283.960 1677.940 1284.220 1678.200 ;
        RECT 1285.800 1677.940 1286.060 1678.200 ;
        RECT 507.940 45.600 508.200 45.860 ;
        RECT 1283.960 45.600 1284.220 45.860 ;
      LAYER met2 ;
        RECT 1286.710 1700.410 1286.990 1704.000 ;
        RECT 1285.860 1700.270 1286.990 1700.410 ;
        RECT 1285.860 1678.230 1286.000 1700.270 ;
        RECT 1286.710 1700.000 1286.990 1700.270 ;
        RECT 1283.960 1677.910 1284.220 1678.230 ;
        RECT 1285.800 1677.910 1286.060 1678.230 ;
        RECT 1284.020 45.890 1284.160 1677.910 ;
        RECT 507.940 45.570 508.200 45.890 ;
        RECT 1283.960 45.570 1284.220 45.890 ;
        RECT 508.000 2.400 508.140 45.570 ;
        RECT 507.790 -4.800 508.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 0.300 ;
=======
      LAYER met1 ;
        RECT 525.850 46.140 526.170 46.200 ;
        RECT 1290.830 46.140 1291.150 46.200 ;
        RECT 525.850 46.000 1291.150 46.140 ;
        RECT 525.850 45.940 526.170 46.000 ;
        RECT 1290.830 45.940 1291.150 46.000 ;
      LAYER via ;
        RECT 525.880 45.940 526.140 46.200 ;
        RECT 1290.860 45.940 1291.120 46.200 ;
      LAYER met2 ;
        RECT 1291.770 1700.410 1292.050 1704.000 ;
        RECT 1290.920 1700.270 1292.050 1700.410 ;
        RECT 1290.920 46.230 1291.060 1700.270 ;
        RECT 1291.770 1700.000 1292.050 1700.270 ;
        RECT 525.880 45.910 526.140 46.230 ;
        RECT 1290.860 45.910 1291.120 46.230 ;
        RECT 525.940 2.400 526.080 45.910 ;
        RECT 525.730 -4.800 526.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 0.300 ;
=======
      LAYER met1 ;
        RECT 1291.290 1678.140 1291.610 1678.200 ;
        RECT 1295.430 1678.140 1295.750 1678.200 ;
        RECT 1291.290 1678.000 1295.750 1678.140 ;
        RECT 1291.290 1677.940 1291.610 1678.000 ;
        RECT 1295.430 1677.940 1295.750 1678.000 ;
        RECT 544.710 52.600 545.030 52.660 ;
        RECT 1291.290 52.600 1291.610 52.660 ;
        RECT 544.710 52.460 1291.610 52.600 ;
        RECT 544.710 52.400 545.030 52.460 ;
        RECT 1291.290 52.400 1291.610 52.460 ;
      LAYER via ;
        RECT 1291.320 1677.940 1291.580 1678.200 ;
        RECT 1295.460 1677.940 1295.720 1678.200 ;
        RECT 544.740 52.400 545.000 52.660 ;
        RECT 1291.320 52.400 1291.580 52.660 ;
      LAYER met2 ;
        RECT 1296.370 1700.410 1296.650 1704.000 ;
        RECT 1295.520 1700.270 1296.650 1700.410 ;
        RECT 1295.520 1678.230 1295.660 1700.270 ;
        RECT 1296.370 1700.000 1296.650 1700.270 ;
        RECT 1291.320 1677.910 1291.580 1678.230 ;
        RECT 1295.460 1677.910 1295.720 1678.230 ;
        RECT 1291.380 52.690 1291.520 1677.910 ;
        RECT 544.740 52.370 545.000 52.690 ;
        RECT 1291.320 52.370 1291.580 52.690 ;
        RECT 544.800 17.410 544.940 52.370 ;
        RECT 543.880 17.270 544.940 17.410 ;
        RECT 543.880 2.400 544.020 17.270 ;
        RECT 543.670 -4.800 544.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 0.300 ;
=======
      LAYER met1 ;
        RECT 565.410 52.940 565.730 53.000 ;
        RECT 1297.730 52.940 1298.050 53.000 ;
        RECT 565.410 52.800 1298.050 52.940 ;
        RECT 565.410 52.740 565.730 52.800 ;
        RECT 1297.730 52.740 1298.050 52.800 ;
        RECT 561.730 15.200 562.050 15.260 ;
        RECT 565.410 15.200 565.730 15.260 ;
        RECT 561.730 15.060 565.730 15.200 ;
        RECT 561.730 15.000 562.050 15.060 ;
        RECT 565.410 15.000 565.730 15.060 ;
      LAYER via ;
        RECT 565.440 52.740 565.700 53.000 ;
        RECT 1297.760 52.740 1298.020 53.000 ;
        RECT 561.760 15.000 562.020 15.260 ;
        RECT 565.440 15.000 565.700 15.260 ;
      LAYER met2 ;
        RECT 1301.430 1700.410 1301.710 1704.000 ;
        RECT 1300.120 1700.270 1301.710 1700.410 ;
        RECT 1300.120 1678.140 1300.260 1700.270 ;
        RECT 1301.430 1700.000 1301.710 1700.270 ;
        RECT 1297.820 1678.000 1300.260 1678.140 ;
        RECT 1297.820 53.030 1297.960 1678.000 ;
        RECT 565.440 52.710 565.700 53.030 ;
        RECT 1297.760 52.710 1298.020 53.030 ;
        RECT 565.500 15.290 565.640 52.710 ;
        RECT 561.760 14.970 562.020 15.290 ;
        RECT 565.440 14.970 565.700 15.290 ;
        RECT 561.820 2.400 561.960 14.970 ;
        RECT 561.610 -4.800 562.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 0.300 ;
=======
      LAYER met1 ;
        RECT 585.650 53.280 585.970 53.340 ;
        RECT 1306.010 53.280 1306.330 53.340 ;
        RECT 585.650 53.140 1306.330 53.280 ;
        RECT 585.650 53.080 585.970 53.140 ;
        RECT 1306.010 53.080 1306.330 53.140 ;
        RECT 579.670 15.540 579.990 15.600 ;
        RECT 585.650 15.540 585.970 15.600 ;
        RECT 579.670 15.400 585.970 15.540 ;
        RECT 579.670 15.340 579.990 15.400 ;
        RECT 585.650 15.340 585.970 15.400 ;
      LAYER via ;
        RECT 585.680 53.080 585.940 53.340 ;
        RECT 1306.040 53.080 1306.300 53.340 ;
        RECT 579.700 15.340 579.960 15.600 ;
        RECT 585.680 15.340 585.940 15.600 ;
      LAYER met2 ;
        RECT 1306.030 1700.000 1306.310 1704.000 ;
        RECT 1306.100 53.370 1306.240 1700.000 ;
        RECT 585.680 53.050 585.940 53.370 ;
        RECT 1306.040 53.050 1306.300 53.370 ;
        RECT 585.740 15.630 585.880 53.050 ;
        RECT 579.700 15.310 579.960 15.630 ;
        RECT 585.680 15.310 585.940 15.630 ;
        RECT 579.760 2.400 579.900 15.310 ;
        RECT 579.550 -4.800 580.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1166.630 1690.720 1166.950 1690.780 ;
        RECT 1171.690 1690.720 1172.010 1690.780 ;
        RECT 1166.630 1690.580 1172.010 1690.720 ;
        RECT 1166.630 1690.520 1166.950 1690.580 ;
        RECT 1171.690 1690.520 1172.010 1690.580 ;
      LAYER via ;
        RECT 1166.660 1690.520 1166.920 1690.780 ;
        RECT 1171.720 1690.520 1171.980 1690.780 ;
      LAYER met2 ;
        RECT 1172.630 1700.410 1172.910 1704.000 ;
        RECT 1171.780 1700.270 1172.910 1700.410 ;
        RECT 1171.780 1690.810 1171.920 1700.270 ;
        RECT 1172.630 1700.000 1172.910 1700.270 ;
        RECT 1166.660 1690.490 1166.920 1690.810 ;
        RECT 1171.720 1690.490 1171.980 1690.810 ;
        RECT 1166.720 39.285 1166.860 1690.490 ;
        RECT 86.110 38.915 86.390 39.285 ;
        RECT 1166.650 38.915 1166.930 39.285 ;
        RECT 86.180 2.400 86.320 38.915 ;
        RECT 85.970 -4.800 86.530 2.400 ;
      LAYER via2 ;
        RECT 86.110 38.960 86.390 39.240 ;
        RECT 1166.650 38.960 1166.930 39.240 ;
      LAYER met3 ;
        RECT 86.085 39.250 86.415 39.265 ;
        RECT 1166.625 39.250 1166.955 39.265 ;
        RECT 86.085 38.950 1166.955 39.250 ;
        RECT 86.085 38.935 86.415 38.950 ;
        RECT 1166.625 38.935 1166.955 38.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 0.300 ;
=======
      LAYER met1 ;
        RECT 599.910 53.620 600.230 53.680 ;
        RECT 1311.990 53.620 1312.310 53.680 ;
        RECT 599.910 53.480 1312.310 53.620 ;
        RECT 599.910 53.420 600.230 53.480 ;
        RECT 1311.990 53.420 1312.310 53.480 ;
        RECT 597.150 15.540 597.470 15.600 ;
        RECT 599.910 15.540 600.230 15.600 ;
        RECT 597.150 15.400 600.230 15.540 ;
        RECT 597.150 15.340 597.470 15.400 ;
        RECT 599.910 15.340 600.230 15.400 ;
      LAYER via ;
        RECT 599.940 53.420 600.200 53.680 ;
        RECT 1312.020 53.420 1312.280 53.680 ;
        RECT 597.180 15.340 597.440 15.600 ;
        RECT 599.940 15.340 600.200 15.600 ;
      LAYER met2 ;
        RECT 1311.090 1700.410 1311.370 1704.000 ;
        RECT 1311.090 1700.270 1312.220 1700.410 ;
        RECT 1311.090 1700.000 1311.370 1700.270 ;
        RECT 1312.080 53.710 1312.220 1700.270 ;
        RECT 599.940 53.390 600.200 53.710 ;
        RECT 1312.020 53.390 1312.280 53.710 ;
        RECT 600.000 15.630 600.140 53.390 ;
        RECT 597.180 15.310 597.440 15.630 ;
        RECT 599.940 15.310 600.200 15.630 ;
        RECT 597.240 2.400 597.380 15.310 ;
        RECT 597.030 -4.800 597.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1311.530 1678.140 1311.850 1678.200 ;
        RECT 1314.750 1678.140 1315.070 1678.200 ;
        RECT 1311.530 1678.000 1315.070 1678.140 ;
        RECT 1311.530 1677.940 1311.850 1678.000 ;
        RECT 1314.750 1677.940 1315.070 1678.000 ;
        RECT 620.610 53.960 620.930 54.020 ;
        RECT 1311.530 53.960 1311.850 54.020 ;
        RECT 620.610 53.820 1311.850 53.960 ;
        RECT 620.610 53.760 620.930 53.820 ;
        RECT 1311.530 53.760 1311.850 53.820 ;
        RECT 615.090 14.860 615.410 14.920 ;
        RECT 620.610 14.860 620.930 14.920 ;
        RECT 615.090 14.720 620.930 14.860 ;
        RECT 615.090 14.660 615.410 14.720 ;
        RECT 620.610 14.660 620.930 14.720 ;
      LAYER via ;
        RECT 1311.560 1677.940 1311.820 1678.200 ;
        RECT 1314.780 1677.940 1315.040 1678.200 ;
        RECT 620.640 53.760 620.900 54.020 ;
        RECT 1311.560 53.760 1311.820 54.020 ;
        RECT 615.120 14.660 615.380 14.920 ;
        RECT 620.640 14.660 620.900 14.920 ;
      LAYER met2 ;
        RECT 1315.690 1700.410 1315.970 1704.000 ;
        RECT 1314.840 1700.270 1315.970 1700.410 ;
        RECT 1314.840 1678.230 1314.980 1700.270 ;
        RECT 1315.690 1700.000 1315.970 1700.270 ;
        RECT 1311.560 1677.910 1311.820 1678.230 ;
        RECT 1314.780 1677.910 1315.040 1678.230 ;
        RECT 1311.620 54.050 1311.760 1677.910 ;
        RECT 620.640 53.730 620.900 54.050 ;
        RECT 1311.560 53.730 1311.820 54.050 ;
        RECT 620.700 14.950 620.840 53.730 ;
        RECT 615.120 14.630 615.380 14.950 ;
        RECT 620.640 14.630 620.900 14.950 ;
        RECT 615.180 2.400 615.320 14.630 ;
        RECT 614.970 -4.800 615.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 0.300 ;
=======
      LAYER li1 ;
        RECT 1175.445 1449.165 1175.615 1497.275 ;
        RECT 1175.445 1256.045 1175.615 1304.155 ;
        RECT 1174.985 765.765 1175.155 807.075 ;
        RECT 1174.985 613.785 1175.155 620.755 ;
        RECT 1175.445 524.365 1175.615 566.015 ;
      LAYER mcon ;
        RECT 1175.445 1497.105 1175.615 1497.275 ;
        RECT 1175.445 1303.985 1175.615 1304.155 ;
        RECT 1174.985 806.905 1175.155 807.075 ;
        RECT 1174.985 620.585 1175.155 620.755 ;
        RECT 1175.445 565.845 1175.615 566.015 ;
      LAYER met1 ;
        RECT 1175.370 1558.940 1175.690 1559.200 ;
        RECT 1175.460 1558.520 1175.600 1558.940 ;
        RECT 1175.370 1558.260 1175.690 1558.520 ;
        RECT 1175.370 1497.260 1175.690 1497.320 ;
        RECT 1175.175 1497.120 1175.690 1497.260 ;
        RECT 1175.370 1497.060 1175.690 1497.120 ;
        RECT 1175.370 1449.320 1175.690 1449.380 ;
        RECT 1175.175 1449.180 1175.690 1449.320 ;
        RECT 1175.370 1449.120 1175.690 1449.180 ;
        RECT 1175.370 1365.820 1175.690 1366.080 ;
        RECT 1175.460 1365.400 1175.600 1365.820 ;
        RECT 1175.370 1365.140 1175.690 1365.400 ;
        RECT 1175.370 1304.140 1175.690 1304.200 ;
        RECT 1175.175 1304.000 1175.690 1304.140 ;
        RECT 1175.370 1303.940 1175.690 1304.000 ;
        RECT 1175.370 1256.200 1175.690 1256.260 ;
        RECT 1175.175 1256.060 1175.690 1256.200 ;
        RECT 1175.370 1256.000 1175.690 1256.060 ;
        RECT 1174.450 1159.300 1174.770 1159.360 ;
        RECT 1175.370 1159.300 1175.690 1159.360 ;
        RECT 1174.450 1159.160 1175.690 1159.300 ;
        RECT 1174.450 1159.100 1174.770 1159.160 ;
        RECT 1175.370 1159.100 1175.690 1159.160 ;
        RECT 1174.450 1062.740 1174.770 1062.800 ;
        RECT 1175.370 1062.740 1175.690 1062.800 ;
        RECT 1174.450 1062.600 1175.690 1062.740 ;
        RECT 1174.450 1062.540 1174.770 1062.600 ;
        RECT 1175.370 1062.540 1175.690 1062.600 ;
        RECT 1175.830 980.120 1176.150 980.180 ;
        RECT 1175.460 979.980 1176.150 980.120 ;
        RECT 1175.460 979.840 1175.600 979.980 ;
        RECT 1175.830 979.920 1176.150 979.980 ;
        RECT 1175.370 979.580 1175.690 979.840 ;
        RECT 1175.370 917.900 1175.690 917.960 ;
        RECT 1175.830 917.900 1176.150 917.960 ;
        RECT 1175.370 917.760 1176.150 917.900 ;
        RECT 1175.370 917.700 1175.690 917.760 ;
        RECT 1175.830 917.700 1176.150 917.760 ;
        RECT 1175.370 869.620 1175.690 869.680 ;
        RECT 1175.830 869.620 1176.150 869.680 ;
        RECT 1175.370 869.480 1176.150 869.620 ;
        RECT 1175.370 869.420 1175.690 869.480 ;
        RECT 1175.830 869.420 1176.150 869.480 ;
        RECT 1174.910 807.060 1175.230 807.120 ;
        RECT 1174.715 806.920 1175.230 807.060 ;
        RECT 1174.910 806.860 1175.230 806.920 ;
        RECT 1174.910 765.920 1175.230 765.980 ;
        RECT 1174.715 765.780 1175.230 765.920 ;
        RECT 1174.910 765.720 1175.230 765.780 ;
        RECT 1174.910 724.580 1175.230 724.840 ;
        RECT 1175.000 724.440 1175.140 724.580 ;
        RECT 1175.370 724.440 1175.690 724.500 ;
        RECT 1175.000 724.300 1175.690 724.440 ;
        RECT 1175.370 724.240 1175.690 724.300 ;
        RECT 1174.910 669.700 1175.230 669.760 ;
        RECT 1175.370 669.700 1175.690 669.760 ;
        RECT 1174.910 669.560 1175.690 669.700 ;
        RECT 1174.910 669.500 1175.230 669.560 ;
        RECT 1175.370 669.500 1175.690 669.560 ;
        RECT 1174.910 620.740 1175.230 620.800 ;
        RECT 1174.715 620.600 1175.230 620.740 ;
        RECT 1174.910 620.540 1175.230 620.600 ;
        RECT 1174.910 613.940 1175.230 614.000 ;
        RECT 1174.715 613.800 1175.230 613.940 ;
        RECT 1174.910 613.740 1175.230 613.800 ;
        RECT 1174.910 566.340 1175.230 566.400 ;
        RECT 1174.910 566.200 1175.600 566.340 ;
        RECT 1174.910 566.140 1175.230 566.200 ;
        RECT 1175.460 566.045 1175.600 566.200 ;
        RECT 1175.385 565.815 1175.675 566.045 ;
        RECT 1175.370 524.520 1175.690 524.580 ;
        RECT 1175.175 524.380 1175.690 524.520 ;
        RECT 1175.370 524.320 1175.690 524.380 ;
        RECT 1175.370 497.120 1175.690 497.380 ;
        RECT 1175.460 496.700 1175.600 497.120 ;
        RECT 1175.370 496.440 1175.690 496.700 ;
        RECT 1175.830 290.060 1176.150 290.320 ;
        RECT 1175.920 289.640 1176.060 290.060 ;
        RECT 1175.830 289.380 1176.150 289.640 ;
        RECT 1174.910 241.640 1175.230 241.700 ;
        RECT 1175.830 241.640 1176.150 241.700 ;
        RECT 1174.910 241.500 1176.150 241.640 ;
        RECT 1174.910 241.440 1175.230 241.500 ;
        RECT 1175.830 241.440 1176.150 241.500 ;
        RECT 1174.910 186.700 1175.230 186.960 ;
        RECT 1175.000 186.560 1175.140 186.700 ;
        RECT 1175.370 186.560 1175.690 186.620 ;
        RECT 1175.000 186.420 1175.690 186.560 ;
        RECT 1175.370 186.360 1175.690 186.420 ;
        RECT 1174.450 73.340 1174.770 73.400 ;
        RECT 1175.370 73.340 1175.690 73.400 ;
        RECT 1174.450 73.200 1175.690 73.340 ;
        RECT 1174.450 73.140 1174.770 73.200 ;
        RECT 1175.370 73.140 1175.690 73.200 ;
      LAYER via ;
        RECT 1175.400 1558.940 1175.660 1559.200 ;
        RECT 1175.400 1558.260 1175.660 1558.520 ;
        RECT 1175.400 1497.060 1175.660 1497.320 ;
        RECT 1175.400 1449.120 1175.660 1449.380 ;
        RECT 1175.400 1365.820 1175.660 1366.080 ;
        RECT 1175.400 1365.140 1175.660 1365.400 ;
        RECT 1175.400 1303.940 1175.660 1304.200 ;
        RECT 1175.400 1256.000 1175.660 1256.260 ;
        RECT 1174.480 1159.100 1174.740 1159.360 ;
        RECT 1175.400 1159.100 1175.660 1159.360 ;
        RECT 1174.480 1062.540 1174.740 1062.800 ;
        RECT 1175.400 1062.540 1175.660 1062.800 ;
        RECT 1175.860 979.920 1176.120 980.180 ;
        RECT 1175.400 979.580 1175.660 979.840 ;
        RECT 1175.400 917.700 1175.660 917.960 ;
        RECT 1175.860 917.700 1176.120 917.960 ;
        RECT 1175.400 869.420 1175.660 869.680 ;
        RECT 1175.860 869.420 1176.120 869.680 ;
        RECT 1174.940 806.860 1175.200 807.120 ;
        RECT 1174.940 765.720 1175.200 765.980 ;
        RECT 1174.940 724.580 1175.200 724.840 ;
        RECT 1175.400 724.240 1175.660 724.500 ;
        RECT 1174.940 669.500 1175.200 669.760 ;
        RECT 1175.400 669.500 1175.660 669.760 ;
        RECT 1174.940 620.540 1175.200 620.800 ;
        RECT 1174.940 613.740 1175.200 614.000 ;
        RECT 1174.940 566.140 1175.200 566.400 ;
        RECT 1175.400 524.320 1175.660 524.580 ;
        RECT 1175.400 497.120 1175.660 497.380 ;
        RECT 1175.400 496.440 1175.660 496.700 ;
        RECT 1175.860 290.060 1176.120 290.320 ;
        RECT 1175.860 289.380 1176.120 289.640 ;
        RECT 1174.940 241.440 1175.200 241.700 ;
        RECT 1175.860 241.440 1176.120 241.700 ;
        RECT 1174.940 186.700 1175.200 186.960 ;
        RECT 1175.400 186.360 1175.660 186.620 ;
        RECT 1174.480 73.140 1174.740 73.400 ;
        RECT 1175.400 73.140 1175.660 73.400 ;
      LAYER met2 ;
        RECT 1179.070 1700.410 1179.350 1704.000 ;
        RECT 1178.220 1700.270 1179.350 1700.410 ;
        RECT 1178.220 1676.610 1178.360 1700.270 ;
        RECT 1179.070 1700.000 1179.350 1700.270 ;
        RECT 1175.460 1676.470 1178.360 1676.610 ;
        RECT 1175.460 1559.230 1175.600 1676.470 ;
        RECT 1175.400 1558.910 1175.660 1559.230 ;
        RECT 1175.400 1558.230 1175.660 1558.550 ;
        RECT 1175.460 1497.350 1175.600 1558.230 ;
        RECT 1175.400 1497.030 1175.660 1497.350 ;
        RECT 1175.400 1449.090 1175.660 1449.410 ;
        RECT 1175.460 1366.110 1175.600 1449.090 ;
        RECT 1175.400 1365.790 1175.660 1366.110 ;
        RECT 1175.400 1365.110 1175.660 1365.430 ;
        RECT 1175.460 1304.230 1175.600 1365.110 ;
        RECT 1175.400 1303.910 1175.660 1304.230 ;
        RECT 1175.400 1255.970 1175.660 1256.290 ;
        RECT 1175.460 1207.525 1175.600 1255.970 ;
        RECT 1174.470 1207.155 1174.750 1207.525 ;
        RECT 1175.390 1207.155 1175.670 1207.525 ;
        RECT 1174.540 1159.390 1174.680 1207.155 ;
        RECT 1174.480 1159.070 1174.740 1159.390 ;
        RECT 1175.400 1159.070 1175.660 1159.390 ;
        RECT 1175.460 1110.965 1175.600 1159.070 ;
        RECT 1174.470 1110.595 1174.750 1110.965 ;
        RECT 1175.390 1110.595 1175.670 1110.965 ;
        RECT 1174.540 1062.830 1174.680 1110.595 ;
        RECT 1174.480 1062.510 1174.740 1062.830 ;
        RECT 1175.400 1062.510 1175.660 1062.830 ;
        RECT 1175.460 1014.290 1175.600 1062.510 ;
        RECT 1175.460 1014.150 1176.060 1014.290 ;
        RECT 1175.920 980.210 1176.060 1014.150 ;
        RECT 1175.860 979.890 1176.120 980.210 ;
        RECT 1175.400 979.550 1175.660 979.870 ;
        RECT 1175.460 917.990 1175.600 979.550 ;
        RECT 1175.400 917.670 1175.660 917.990 ;
        RECT 1175.860 917.670 1176.120 917.990 ;
        RECT 1175.920 869.710 1176.060 917.670 ;
        RECT 1175.400 869.390 1175.660 869.710 ;
        RECT 1175.860 869.390 1176.120 869.710 ;
        RECT 1175.460 815.165 1175.600 869.390 ;
        RECT 1175.390 814.795 1175.670 815.165 ;
        RECT 1174.930 814.115 1175.210 814.485 ;
        RECT 1175.000 807.150 1175.140 814.115 ;
        RECT 1174.940 806.830 1175.200 807.150 ;
        RECT 1174.940 765.690 1175.200 766.010 ;
        RECT 1175.000 724.870 1175.140 765.690 ;
        RECT 1174.940 724.550 1175.200 724.870 ;
        RECT 1175.400 724.210 1175.660 724.530 ;
        RECT 1175.460 669.790 1175.600 724.210 ;
        RECT 1174.940 669.470 1175.200 669.790 ;
        RECT 1175.400 669.470 1175.660 669.790 ;
        RECT 1175.000 620.830 1175.140 669.470 ;
        RECT 1174.940 620.510 1175.200 620.830 ;
        RECT 1174.940 613.710 1175.200 614.030 ;
        RECT 1175.000 566.430 1175.140 613.710 ;
        RECT 1174.940 566.110 1175.200 566.430 ;
        RECT 1175.400 524.290 1175.660 524.610 ;
        RECT 1175.460 497.410 1175.600 524.290 ;
        RECT 1175.400 497.090 1175.660 497.410 ;
        RECT 1175.400 496.410 1175.660 496.730 ;
        RECT 1175.460 435.725 1175.600 496.410 ;
        RECT 1175.390 435.355 1175.670 435.725 ;
        RECT 1174.930 434.675 1175.210 435.045 ;
        RECT 1175.000 409.090 1175.140 434.675 ;
        RECT 1175.000 408.950 1176.060 409.090 ;
        RECT 1175.920 290.350 1176.060 408.950 ;
        RECT 1175.860 290.030 1176.120 290.350 ;
        RECT 1175.860 289.350 1176.120 289.670 ;
        RECT 1175.920 241.730 1176.060 289.350 ;
        RECT 1174.940 241.410 1175.200 241.730 ;
        RECT 1175.860 241.410 1176.120 241.730 ;
        RECT 1175.000 186.990 1175.140 241.410 ;
        RECT 1174.940 186.670 1175.200 186.990 ;
        RECT 1175.400 186.330 1175.660 186.650 ;
        RECT 1175.460 73.430 1175.600 186.330 ;
        RECT 1174.480 73.110 1174.740 73.430 ;
        RECT 1175.400 73.110 1175.660 73.430 ;
        RECT 1174.540 39.965 1174.680 73.110 ;
        RECT 109.570 39.595 109.850 39.965 ;
        RECT 1174.470 39.595 1174.750 39.965 ;
        RECT 109.640 2.400 109.780 39.595 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 1174.470 1207.200 1174.750 1207.480 ;
        RECT 1175.390 1207.200 1175.670 1207.480 ;
        RECT 1174.470 1110.640 1174.750 1110.920 ;
        RECT 1175.390 1110.640 1175.670 1110.920 ;
        RECT 1175.390 814.840 1175.670 815.120 ;
        RECT 1174.930 814.160 1175.210 814.440 ;
        RECT 1175.390 435.400 1175.670 435.680 ;
        RECT 1174.930 434.720 1175.210 435.000 ;
        RECT 109.570 39.640 109.850 39.920 ;
        RECT 1174.470 39.640 1174.750 39.920 ;
      LAYER met3 ;
        RECT 1174.445 1207.490 1174.775 1207.505 ;
        RECT 1175.365 1207.490 1175.695 1207.505 ;
        RECT 1174.445 1207.190 1175.695 1207.490 ;
        RECT 1174.445 1207.175 1174.775 1207.190 ;
        RECT 1175.365 1207.175 1175.695 1207.190 ;
        RECT 1174.445 1110.930 1174.775 1110.945 ;
        RECT 1175.365 1110.930 1175.695 1110.945 ;
        RECT 1174.445 1110.630 1175.695 1110.930 ;
        RECT 1174.445 1110.615 1174.775 1110.630 ;
        RECT 1175.365 1110.615 1175.695 1110.630 ;
        RECT 1175.365 815.130 1175.695 815.145 ;
        RECT 1175.150 814.815 1175.695 815.130 ;
        RECT 1175.150 814.465 1175.450 814.815 ;
        RECT 1174.905 814.150 1175.450 814.465 ;
        RECT 1174.905 814.135 1175.235 814.150 ;
        RECT 1175.365 435.690 1175.695 435.705 ;
        RECT 1175.150 435.375 1175.695 435.690 ;
        RECT 1175.150 435.025 1175.450 435.375 ;
        RECT 1174.905 434.710 1175.450 435.025 ;
        RECT 1174.905 434.695 1175.235 434.710 ;
        RECT 109.545 39.930 109.875 39.945 ;
        RECT 1174.445 39.930 1174.775 39.945 ;
        RECT 109.545 39.630 1174.775 39.930 ;
        RECT 109.545 39.615 109.875 39.630 ;
        RECT 1174.445 39.615 1174.775 39.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 0.300 ;
=======
      LAYER li1 ;
        RECT 1181.885 814.385 1182.055 821.355 ;
        RECT 1181.425 572.645 1181.595 620.755 ;
        RECT 1181.885 324.445 1182.055 372.215 ;
        RECT 1181.425 131.325 1181.595 138.635 ;
      LAYER mcon ;
        RECT 1181.885 821.185 1182.055 821.355 ;
        RECT 1181.425 620.585 1181.595 620.755 ;
        RECT 1181.885 372.045 1182.055 372.215 ;
        RECT 1181.425 138.465 1181.595 138.635 ;
      LAYER met1 ;
        RECT 1181.810 821.340 1182.130 821.400 ;
        RECT 1181.615 821.200 1182.130 821.340 ;
        RECT 1181.810 821.140 1182.130 821.200 ;
        RECT 1181.810 814.540 1182.130 814.600 ;
        RECT 1181.615 814.400 1182.130 814.540 ;
        RECT 1181.810 814.340 1182.130 814.400 ;
        RECT 1181.810 813.860 1182.130 813.920 ;
        RECT 1182.270 813.860 1182.590 813.920 ;
        RECT 1181.810 813.720 1182.590 813.860 ;
        RECT 1181.810 813.660 1182.130 813.720 ;
        RECT 1182.270 813.660 1182.590 813.720 ;
        RECT 1181.350 620.740 1181.670 620.800 ;
        RECT 1181.155 620.600 1181.670 620.740 ;
        RECT 1181.350 620.540 1181.670 620.600 ;
        RECT 1181.365 572.800 1181.655 572.845 ;
        RECT 1181.810 572.800 1182.130 572.860 ;
        RECT 1181.365 572.660 1182.130 572.800 ;
        RECT 1181.365 572.615 1181.655 572.660 ;
        RECT 1181.810 572.600 1182.130 572.660 ;
        RECT 1180.890 421.160 1181.210 421.220 ;
        RECT 1182.730 421.160 1183.050 421.220 ;
        RECT 1180.890 421.020 1183.050 421.160 ;
        RECT 1180.890 420.960 1181.210 421.020 ;
        RECT 1182.730 420.960 1183.050 421.020 ;
        RECT 1182.270 372.340 1182.590 372.600 ;
        RECT 1181.825 372.200 1182.115 372.245 ;
        RECT 1182.360 372.200 1182.500 372.340 ;
        RECT 1181.825 372.060 1182.500 372.200 ;
        RECT 1181.825 372.015 1182.115 372.060 ;
        RECT 1181.810 324.600 1182.130 324.660 ;
        RECT 1181.615 324.460 1182.130 324.600 ;
        RECT 1181.810 324.400 1182.130 324.460 ;
        RECT 1181.365 138.620 1181.655 138.665 ;
        RECT 1181.810 138.620 1182.130 138.680 ;
        RECT 1181.365 138.480 1182.130 138.620 ;
        RECT 1181.365 138.435 1181.655 138.480 ;
        RECT 1181.810 138.420 1182.130 138.480 ;
        RECT 1181.350 131.480 1181.670 131.540 ;
        RECT 1181.155 131.340 1181.670 131.480 ;
        RECT 1181.350 131.280 1181.670 131.340 ;
      LAYER via ;
        RECT 1181.840 821.140 1182.100 821.400 ;
        RECT 1181.840 814.340 1182.100 814.600 ;
        RECT 1181.840 813.660 1182.100 813.920 ;
        RECT 1182.300 813.660 1182.560 813.920 ;
        RECT 1181.380 620.540 1181.640 620.800 ;
        RECT 1181.840 572.600 1182.100 572.860 ;
        RECT 1180.920 420.960 1181.180 421.220 ;
        RECT 1182.760 420.960 1183.020 421.220 ;
        RECT 1182.300 372.340 1182.560 372.600 ;
        RECT 1181.840 324.400 1182.100 324.660 ;
        RECT 1181.840 138.420 1182.100 138.680 ;
        RECT 1181.380 131.280 1181.640 131.540 ;
      LAYER met2 ;
        RECT 1185.510 1700.410 1185.790 1704.000 ;
        RECT 1185.120 1700.270 1185.790 1700.410 ;
        RECT 1185.120 1676.610 1185.260 1700.270 ;
        RECT 1185.510 1700.000 1185.790 1700.270 ;
        RECT 1181.440 1676.470 1185.260 1676.610 ;
        RECT 1181.440 1655.530 1181.580 1676.470 ;
        RECT 1181.440 1655.390 1182.040 1655.530 ;
        RECT 1181.900 1511.370 1182.040 1655.390 ;
        RECT 1181.440 1511.230 1182.040 1511.370 ;
        RECT 1181.440 1510.690 1181.580 1511.230 ;
        RECT 1181.440 1510.550 1182.040 1510.690 ;
        RECT 1181.900 1414.810 1182.040 1510.550 ;
        RECT 1181.440 1414.670 1182.040 1414.810 ;
        RECT 1181.440 1414.130 1181.580 1414.670 ;
        RECT 1181.440 1413.990 1182.040 1414.130 ;
        RECT 1181.900 1318.250 1182.040 1413.990 ;
        RECT 1181.440 1318.110 1182.040 1318.250 ;
        RECT 1181.440 1317.570 1181.580 1318.110 ;
        RECT 1181.440 1317.430 1182.040 1317.570 ;
        RECT 1181.900 1221.690 1182.040 1317.430 ;
        RECT 1181.440 1221.550 1182.040 1221.690 ;
        RECT 1181.440 1221.010 1181.580 1221.550 ;
        RECT 1181.440 1220.870 1182.040 1221.010 ;
        RECT 1181.900 1125.130 1182.040 1220.870 ;
        RECT 1181.440 1124.990 1182.040 1125.130 ;
        RECT 1181.440 1124.450 1181.580 1124.990 ;
        RECT 1181.440 1124.310 1182.040 1124.450 ;
        RECT 1181.900 1028.570 1182.040 1124.310 ;
        RECT 1181.440 1028.430 1182.040 1028.570 ;
        RECT 1181.440 1027.890 1181.580 1028.430 ;
        RECT 1181.440 1027.750 1182.040 1027.890 ;
        RECT 1181.900 932.010 1182.040 1027.750 ;
        RECT 1181.440 931.870 1182.040 932.010 ;
        RECT 1181.440 931.330 1181.580 931.870 ;
        RECT 1181.440 931.190 1182.040 931.330 ;
        RECT 1181.900 821.430 1182.040 931.190 ;
        RECT 1181.840 821.110 1182.100 821.430 ;
        RECT 1181.840 814.310 1182.100 814.630 ;
        RECT 1181.900 813.950 1182.040 814.310 ;
        RECT 1181.840 813.630 1182.100 813.950 ;
        RECT 1182.300 813.630 1182.560 813.950 ;
        RECT 1182.360 724.725 1182.500 813.630 ;
        RECT 1181.370 724.355 1181.650 724.725 ;
        RECT 1182.290 724.355 1182.570 724.725 ;
        RECT 1181.440 628.845 1181.580 724.355 ;
        RECT 1181.370 628.475 1181.650 628.845 ;
        RECT 1181.370 627.795 1181.650 628.165 ;
        RECT 1181.440 620.830 1181.580 627.795 ;
        RECT 1181.380 620.510 1181.640 620.830 ;
        RECT 1181.840 572.570 1182.100 572.890 ;
        RECT 1181.900 524.690 1182.040 572.570 ;
        RECT 1181.440 524.550 1182.040 524.690 ;
        RECT 1181.440 496.980 1181.580 524.550 ;
        RECT 1180.980 496.840 1181.580 496.980 ;
        RECT 1180.980 470.405 1181.120 496.840 ;
        RECT 1180.910 470.035 1181.190 470.405 ;
        RECT 1180.910 468.675 1181.190 469.045 ;
        RECT 1180.980 421.250 1181.120 468.675 ;
        RECT 1180.920 420.930 1181.180 421.250 ;
        RECT 1182.760 420.930 1183.020 421.250 ;
        RECT 1182.820 379.170 1182.960 420.930 ;
        RECT 1182.360 379.030 1182.960 379.170 ;
        RECT 1182.360 372.630 1182.500 379.030 ;
        RECT 1182.300 372.310 1182.560 372.630 ;
        RECT 1181.840 324.370 1182.100 324.690 ;
        RECT 1181.900 138.710 1182.040 324.370 ;
        RECT 1181.840 138.390 1182.100 138.710 ;
        RECT 1181.380 131.250 1181.640 131.570 ;
        RECT 1181.440 40.645 1181.580 131.250 ;
        RECT 133.490 40.275 133.770 40.645 ;
        RECT 1181.370 40.275 1181.650 40.645 ;
        RECT 133.560 2.400 133.700 40.275 ;
        RECT 133.350 -4.800 133.910 2.400 ;
      LAYER via2 ;
        RECT 1181.370 724.400 1181.650 724.680 ;
        RECT 1182.290 724.400 1182.570 724.680 ;
        RECT 1181.370 628.520 1181.650 628.800 ;
        RECT 1181.370 627.840 1181.650 628.120 ;
        RECT 1180.910 470.080 1181.190 470.360 ;
        RECT 1180.910 468.720 1181.190 469.000 ;
        RECT 133.490 40.320 133.770 40.600 ;
        RECT 1181.370 40.320 1181.650 40.600 ;
      LAYER met3 ;
        RECT 1181.345 724.690 1181.675 724.705 ;
        RECT 1182.265 724.690 1182.595 724.705 ;
        RECT 1181.345 724.390 1182.595 724.690 ;
        RECT 1181.345 724.375 1181.675 724.390 ;
        RECT 1182.265 724.375 1182.595 724.390 ;
        RECT 1181.345 628.810 1181.675 628.825 ;
        RECT 1181.345 628.495 1181.890 628.810 ;
        RECT 1181.590 628.145 1181.890 628.495 ;
        RECT 1181.345 627.830 1181.890 628.145 ;
        RECT 1181.345 627.815 1181.675 627.830 ;
        RECT 1180.885 470.370 1181.215 470.385 ;
        RECT 1180.885 470.070 1181.890 470.370 ;
        RECT 1180.885 470.055 1181.215 470.070 ;
        RECT 1180.885 469.010 1181.215 469.025 ;
        RECT 1181.590 469.010 1181.890 470.070 ;
        RECT 1180.885 468.710 1181.890 469.010 ;
        RECT 1180.885 468.695 1181.215 468.710 ;
        RECT 133.465 40.610 133.795 40.625 ;
        RECT 1181.345 40.610 1181.675 40.625 ;
        RECT 133.465 40.310 1181.675 40.610 ;
        RECT 133.465 40.295 133.795 40.310 ;
        RECT 1181.345 40.295 1181.675 40.310 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1187.790 1694.120 1188.110 1694.180 ;
        RECT 1190.550 1694.120 1190.870 1694.180 ;
        RECT 1187.790 1693.980 1190.870 1694.120 ;
        RECT 1187.790 1693.920 1188.110 1693.980 ;
        RECT 1190.550 1693.920 1190.870 1693.980 ;
      LAYER via ;
        RECT 1187.820 1693.920 1188.080 1694.180 ;
        RECT 1190.580 1693.920 1190.840 1694.180 ;
      LAYER met2 ;
        RECT 1190.570 1700.000 1190.850 1704.000 ;
        RECT 1190.640 1694.210 1190.780 1700.000 ;
        RECT 1187.820 1693.890 1188.080 1694.210 ;
        RECT 1190.580 1693.890 1190.840 1694.210 ;
        RECT 1187.880 45.405 1188.020 1693.890 ;
        RECT 151.430 45.035 151.710 45.405 ;
        RECT 1187.810 45.035 1188.090 45.405 ;
        RECT 151.500 2.400 151.640 45.035 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 151.430 45.080 151.710 45.360 ;
        RECT 1187.810 45.080 1188.090 45.360 ;
      LAYER met3 ;
        RECT 151.405 45.370 151.735 45.385 ;
        RECT 1187.785 45.370 1188.115 45.385 ;
        RECT 151.405 45.070 1188.115 45.370 ;
        RECT 151.405 45.055 151.735 45.070 ;
        RECT 1187.785 45.055 1188.115 45.070 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 169.230 -4.800 169.790 0.300 ;
=======
        RECT 1195.170 1700.410 1195.450 1704.000 ;
        RECT 1194.780 1700.270 1195.450 1700.410 ;
        RECT 1194.780 46.085 1194.920 1700.270 ;
        RECT 1195.170 1700.000 1195.450 1700.270 ;
        RECT 169.370 45.715 169.650 46.085 ;
        RECT 1194.710 45.715 1194.990 46.085 ;
        RECT 169.440 2.400 169.580 45.715 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 169.370 45.760 169.650 46.040 ;
        RECT 1194.710 45.760 1194.990 46.040 ;
      LAYER met3 ;
        RECT 169.345 46.050 169.675 46.065 ;
        RECT 1194.685 46.050 1195.015 46.065 ;
        RECT 169.345 45.750 1195.015 46.050 ;
        RECT 169.345 45.735 169.675 45.750 ;
        RECT 1194.685 45.735 1195.015 45.750 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 0.300 ;
=======
      LAYER li1 ;
        RECT 1196.145 675.665 1196.315 717.655 ;
        RECT 1196.605 469.285 1196.775 517.395 ;
        RECT 1196.145 385.645 1196.315 427.635 ;
      LAYER mcon ;
        RECT 1196.145 717.485 1196.315 717.655 ;
        RECT 1196.605 517.225 1196.775 517.395 ;
        RECT 1196.145 427.465 1196.315 427.635 ;
      LAYER met1 ;
        RECT 1196.530 1558.940 1196.850 1559.200 ;
        RECT 1196.620 1558.520 1196.760 1558.940 ;
        RECT 1196.530 1558.260 1196.850 1558.520 ;
        RECT 1196.530 1462.380 1196.850 1462.640 ;
        RECT 1196.620 1461.960 1196.760 1462.380 ;
        RECT 1196.530 1461.700 1196.850 1461.960 ;
        RECT 1196.530 1365.820 1196.850 1366.080 ;
        RECT 1196.620 1365.400 1196.760 1365.820 ;
        RECT 1196.530 1365.140 1196.850 1365.400 ;
        RECT 1196.530 1269.260 1196.850 1269.520 ;
        RECT 1196.620 1268.840 1196.760 1269.260 ;
        RECT 1196.530 1268.580 1196.850 1268.840 ;
        RECT 1196.530 1172.700 1196.850 1172.960 ;
        RECT 1196.620 1172.280 1196.760 1172.700 ;
        RECT 1196.530 1172.020 1196.850 1172.280 ;
        RECT 1196.530 1076.140 1196.850 1076.400 ;
        RECT 1196.620 1075.720 1196.760 1076.140 ;
        RECT 1196.530 1075.460 1196.850 1075.720 ;
        RECT 1196.070 772.720 1196.390 772.780 ;
        RECT 1196.530 772.720 1196.850 772.780 ;
        RECT 1196.070 772.580 1196.850 772.720 ;
        RECT 1196.070 772.520 1196.390 772.580 ;
        RECT 1196.530 772.520 1196.850 772.580 ;
        RECT 1196.070 717.640 1196.390 717.700 ;
        RECT 1195.875 717.500 1196.390 717.640 ;
        RECT 1196.070 717.440 1196.390 717.500 ;
        RECT 1196.085 675.820 1196.375 675.865 ;
        RECT 1196.990 675.820 1197.310 675.880 ;
        RECT 1196.085 675.680 1197.310 675.820 ;
        RECT 1196.085 675.635 1196.375 675.680 ;
        RECT 1196.990 675.620 1197.310 675.680 ;
        RECT 1196.530 628.220 1196.850 628.280 ;
        RECT 1196.990 628.220 1197.310 628.280 ;
        RECT 1196.530 628.080 1197.310 628.220 ;
        RECT 1196.530 628.020 1196.850 628.080 ;
        RECT 1196.990 628.020 1197.310 628.080 ;
        RECT 1196.070 572.460 1196.390 572.520 ;
        RECT 1196.990 572.460 1197.310 572.520 ;
        RECT 1196.070 572.320 1197.310 572.460 ;
        RECT 1196.070 572.260 1196.390 572.320 ;
        RECT 1196.990 572.260 1197.310 572.320 ;
        RECT 1196.530 517.380 1196.850 517.440 ;
        RECT 1196.335 517.240 1196.850 517.380 ;
        RECT 1196.530 517.180 1196.850 517.240 ;
        RECT 1196.530 469.440 1196.850 469.500 ;
        RECT 1196.335 469.300 1196.850 469.440 ;
        RECT 1196.530 469.240 1196.850 469.300 ;
        RECT 1196.070 427.620 1196.390 427.680 ;
        RECT 1195.875 427.480 1196.390 427.620 ;
        RECT 1196.070 427.420 1196.390 427.480 ;
        RECT 1196.085 385.800 1196.375 385.845 ;
        RECT 1196.990 385.800 1197.310 385.860 ;
        RECT 1196.085 385.660 1197.310 385.800 ;
        RECT 1196.085 385.615 1196.375 385.660 ;
        RECT 1196.990 385.600 1197.310 385.660 ;
        RECT 1196.530 338.200 1196.850 338.260 ;
        RECT 1196.990 338.200 1197.310 338.260 ;
        RECT 1196.530 338.060 1197.310 338.200 ;
        RECT 1196.530 338.000 1196.850 338.060 ;
        RECT 1196.990 338.000 1197.310 338.060 ;
        RECT 1196.070 158.820 1196.390 159.080 ;
        RECT 1196.160 158.000 1196.300 158.820 ;
        RECT 1196.530 158.000 1196.850 158.060 ;
        RECT 1196.160 157.860 1196.850 158.000 ;
        RECT 1196.530 157.800 1196.850 157.860 ;
        RECT 1196.530 137.740 1196.850 138.000 ;
        RECT 1196.620 137.320 1196.760 137.740 ;
        RECT 1196.530 137.060 1196.850 137.320 ;
      LAYER via ;
        RECT 1196.560 1558.940 1196.820 1559.200 ;
        RECT 1196.560 1558.260 1196.820 1558.520 ;
        RECT 1196.560 1462.380 1196.820 1462.640 ;
        RECT 1196.560 1461.700 1196.820 1461.960 ;
        RECT 1196.560 1365.820 1196.820 1366.080 ;
        RECT 1196.560 1365.140 1196.820 1365.400 ;
        RECT 1196.560 1269.260 1196.820 1269.520 ;
        RECT 1196.560 1268.580 1196.820 1268.840 ;
        RECT 1196.560 1172.700 1196.820 1172.960 ;
        RECT 1196.560 1172.020 1196.820 1172.280 ;
        RECT 1196.560 1076.140 1196.820 1076.400 ;
        RECT 1196.560 1075.460 1196.820 1075.720 ;
        RECT 1196.100 772.520 1196.360 772.780 ;
        RECT 1196.560 772.520 1196.820 772.780 ;
        RECT 1196.100 717.440 1196.360 717.700 ;
        RECT 1197.020 675.620 1197.280 675.880 ;
        RECT 1196.560 628.020 1196.820 628.280 ;
        RECT 1197.020 628.020 1197.280 628.280 ;
        RECT 1196.100 572.260 1196.360 572.520 ;
        RECT 1197.020 572.260 1197.280 572.520 ;
        RECT 1196.560 517.180 1196.820 517.440 ;
        RECT 1196.560 469.240 1196.820 469.500 ;
        RECT 1196.100 427.420 1196.360 427.680 ;
        RECT 1197.020 385.600 1197.280 385.860 ;
        RECT 1196.560 338.000 1196.820 338.260 ;
        RECT 1197.020 338.000 1197.280 338.260 ;
        RECT 1196.100 158.820 1196.360 159.080 ;
        RECT 1196.560 157.800 1196.820 158.060 ;
        RECT 1196.560 137.740 1196.820 138.000 ;
        RECT 1196.560 137.060 1196.820 137.320 ;
      LAYER met2 ;
        RECT 1200.230 1700.410 1200.510 1704.000 ;
        RECT 1199.380 1700.270 1200.510 1700.410 ;
        RECT 1199.380 1677.290 1199.520 1700.270 ;
        RECT 1200.230 1700.000 1200.510 1700.270 ;
        RECT 1196.620 1677.150 1199.520 1677.290 ;
        RECT 1196.620 1559.230 1196.760 1677.150 ;
        RECT 1196.560 1558.910 1196.820 1559.230 ;
        RECT 1196.560 1558.230 1196.820 1558.550 ;
        RECT 1196.620 1462.670 1196.760 1558.230 ;
        RECT 1196.560 1462.350 1196.820 1462.670 ;
        RECT 1196.560 1461.670 1196.820 1461.990 ;
        RECT 1196.620 1366.110 1196.760 1461.670 ;
        RECT 1196.560 1365.790 1196.820 1366.110 ;
        RECT 1196.560 1365.110 1196.820 1365.430 ;
        RECT 1196.620 1269.550 1196.760 1365.110 ;
        RECT 1196.560 1269.230 1196.820 1269.550 ;
        RECT 1196.560 1268.550 1196.820 1268.870 ;
        RECT 1196.620 1172.990 1196.760 1268.550 ;
        RECT 1196.560 1172.670 1196.820 1172.990 ;
        RECT 1196.560 1171.990 1196.820 1172.310 ;
        RECT 1196.620 1076.430 1196.760 1171.990 ;
        RECT 1196.560 1076.110 1196.820 1076.430 ;
        RECT 1196.560 1075.430 1196.820 1075.750 ;
        RECT 1196.620 772.810 1196.760 1075.430 ;
        RECT 1196.100 772.490 1196.360 772.810 ;
        RECT 1196.560 772.490 1196.820 772.810 ;
        RECT 1196.160 717.730 1196.300 772.490 ;
        RECT 1196.100 717.410 1196.360 717.730 ;
        RECT 1197.020 675.590 1197.280 675.910 ;
        RECT 1197.080 628.310 1197.220 675.590 ;
        RECT 1196.560 627.990 1196.820 628.310 ;
        RECT 1197.020 627.990 1197.280 628.310 ;
        RECT 1196.620 572.970 1196.760 627.990 ;
        RECT 1196.160 572.830 1196.760 572.970 ;
        RECT 1196.160 572.550 1196.300 572.830 ;
        RECT 1196.100 572.230 1196.360 572.550 ;
        RECT 1197.020 572.230 1197.280 572.550 ;
        RECT 1197.080 547.810 1197.220 572.230 ;
        RECT 1196.620 547.670 1197.220 547.810 ;
        RECT 1196.620 517.470 1196.760 547.670 ;
        RECT 1196.560 517.150 1196.820 517.470 ;
        RECT 1196.560 469.210 1196.820 469.530 ;
        RECT 1196.620 435.725 1196.760 469.210 ;
        RECT 1196.550 435.355 1196.830 435.725 ;
        RECT 1196.090 434.675 1196.370 435.045 ;
        RECT 1196.160 427.710 1196.300 434.675 ;
        RECT 1196.100 427.390 1196.360 427.710 ;
        RECT 1197.020 385.570 1197.280 385.890 ;
        RECT 1197.080 338.290 1197.220 385.570 ;
        RECT 1196.560 337.970 1196.820 338.290 ;
        RECT 1197.020 337.970 1197.280 338.290 ;
        RECT 1196.620 186.730 1196.760 337.970 ;
        RECT 1196.160 186.590 1196.760 186.730 ;
        RECT 1196.160 159.110 1196.300 186.590 ;
        RECT 1196.100 158.790 1196.360 159.110 ;
        RECT 1196.560 157.770 1196.820 158.090 ;
        RECT 1196.620 138.030 1196.760 157.770 ;
        RECT 1196.560 137.710 1196.820 138.030 ;
        RECT 1196.560 137.030 1196.820 137.350 ;
        RECT 1196.620 51.525 1196.760 137.030 ;
        RECT 186.850 51.155 187.130 51.525 ;
        RECT 1196.550 51.155 1196.830 51.525 ;
        RECT 186.920 2.400 187.060 51.155 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 1196.550 435.400 1196.830 435.680 ;
        RECT 1196.090 434.720 1196.370 435.000 ;
        RECT 186.850 51.200 187.130 51.480 ;
        RECT 1196.550 51.200 1196.830 51.480 ;
      LAYER met3 ;
        RECT 1196.525 435.690 1196.855 435.705 ;
        RECT 1196.310 435.375 1196.855 435.690 ;
        RECT 1196.310 435.025 1196.610 435.375 ;
        RECT 1196.065 434.710 1196.610 435.025 ;
        RECT 1196.065 434.695 1196.395 434.710 ;
        RECT 186.825 51.490 187.155 51.505 ;
        RECT 1196.525 51.490 1196.855 51.505 ;
        RECT 186.825 51.190 1196.855 51.490 ;
        RECT 186.825 51.175 187.155 51.190 ;
        RECT 1196.525 51.175 1196.855 51.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 204.650 -4.800 205.210 0.300 ;
=======
        RECT 1204.830 1700.410 1205.110 1704.000 ;
        RECT 1203.980 1700.270 1205.110 1700.410 ;
        RECT 1203.980 1678.140 1204.120 1700.270 ;
        RECT 1204.830 1700.000 1205.110 1700.270 ;
        RECT 1201.220 1678.000 1204.120 1678.140 ;
        RECT 1201.220 52.205 1201.360 1678.000 ;
        RECT 204.790 51.835 205.070 52.205 ;
        RECT 1201.150 51.835 1201.430 52.205 ;
        RECT 204.860 2.400 205.000 51.835 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 204.790 51.880 205.070 52.160 ;
        RECT 1201.150 51.880 1201.430 52.160 ;
      LAYER met3 ;
        RECT 204.765 52.170 205.095 52.185 ;
        RECT 1201.125 52.170 1201.455 52.185 ;
        RECT 204.765 51.870 1201.455 52.170 ;
        RECT 204.765 51.855 205.095 51.870 ;
        RECT 1201.125 51.855 1201.455 51.870 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 0.300 ;
=======
      LAYER met1 ;
        RECT 222.710 20.640 223.030 20.700 ;
        RECT 227.310 20.640 227.630 20.700 ;
        RECT 222.710 20.500 227.630 20.640 ;
        RECT 222.710 20.440 223.030 20.500 ;
        RECT 227.310 20.440 227.630 20.500 ;
      LAYER via ;
        RECT 222.740 20.440 223.000 20.700 ;
        RECT 227.340 20.440 227.600 20.700 ;
      LAYER met2 ;
        RECT 1209.890 1700.410 1210.170 1704.000 ;
        RECT 1209.500 1700.270 1210.170 1700.410 ;
        RECT 1209.500 52.885 1209.640 1700.270 ;
        RECT 1209.890 1700.000 1210.170 1700.270 ;
        RECT 227.330 52.515 227.610 52.885 ;
        RECT 1209.430 52.515 1209.710 52.885 ;
        RECT 227.400 20.730 227.540 52.515 ;
        RECT 222.740 20.410 223.000 20.730 ;
        RECT 227.340 20.410 227.600 20.730 ;
        RECT 222.800 2.400 222.940 20.410 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 227.330 52.560 227.610 52.840 ;
        RECT 1209.430 52.560 1209.710 52.840 ;
      LAYER met3 ;
        RECT 227.305 52.850 227.635 52.865 ;
        RECT 1209.405 52.850 1209.735 52.865 ;
        RECT 227.305 52.550 1209.735 52.850 ;
        RECT 227.305 52.535 227.635 52.550 ;
        RECT 1209.405 52.535 1209.735 52.550 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 20.190 -4.800 20.750 0.300 ;
=======
        RECT 1155.150 1700.410 1155.430 1704.000 ;
        RECT 1154.300 1700.270 1155.430 1700.410 ;
        RECT 1154.300 37.925 1154.440 1700.270 ;
        RECT 1155.150 1700.000 1155.430 1700.270 ;
        RECT 20.330 37.555 20.610 37.925 ;
        RECT 1154.230 37.555 1154.510 37.925 ;
        RECT 20.400 2.400 20.540 37.555 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 20.330 37.600 20.610 37.880 ;
        RECT 1154.230 37.600 1154.510 37.880 ;
      LAYER met3 ;
        RECT 20.305 37.890 20.635 37.905 ;
        RECT 1154.205 37.890 1154.535 37.905 ;
        RECT 20.305 37.590 1154.535 37.890 ;
        RECT 20.305 37.575 20.635 37.590 ;
        RECT 1154.205 37.575 1154.535 37.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 44.110 -4.800 44.670 0.300 ;
=======
        RECT 1161.590 1700.410 1161.870 1704.000 ;
        RECT 1160.740 1700.270 1161.870 1700.410 ;
        RECT 1160.740 44.725 1160.880 1700.270 ;
        RECT 1161.590 1700.000 1161.870 1700.270 ;
        RECT 44.250 44.355 44.530 44.725 ;
        RECT 1160.670 44.355 1160.950 44.725 ;
        RECT 44.320 2.400 44.460 44.355 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 44.250 44.400 44.530 44.680 ;
        RECT 1160.670 44.400 1160.950 44.680 ;
      LAYER met3 ;
        RECT 44.225 44.690 44.555 44.705 ;
        RECT 1160.645 44.690 1160.975 44.705 ;
        RECT 44.225 44.390 1160.975 44.690 ;
        RECT 44.225 44.375 44.555 44.390 ;
        RECT 1160.645 44.375 1160.975 44.390 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 246.510 -4.800 247.070 0.300 ;
=======
        RECT 1216.330 1700.410 1216.610 1704.000 ;
        RECT 1215.940 1700.270 1216.610 1700.410 ;
        RECT 1215.940 53.565 1216.080 1700.270 ;
        RECT 1216.330 1700.000 1216.610 1700.270 ;
        RECT 248.030 53.195 248.310 53.565 ;
        RECT 1215.870 53.195 1216.150 53.565 ;
        RECT 248.100 16.730 248.240 53.195 ;
        RECT 246.720 16.590 248.240 16.730 ;
        RECT 246.720 2.400 246.860 16.590 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 248.030 53.240 248.310 53.520 ;
        RECT 1215.870 53.240 1216.150 53.520 ;
      LAYER met3 ;
        RECT 248.005 53.530 248.335 53.545 ;
        RECT 1215.845 53.530 1216.175 53.545 ;
        RECT 248.005 53.230 1216.175 53.530 ;
        RECT 248.005 53.215 248.335 53.230 ;
        RECT 1215.845 53.215 1216.175 53.230 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1215.390 1678.480 1215.710 1678.540 ;
        RECT 1219.990 1678.480 1220.310 1678.540 ;
        RECT 1215.390 1678.340 1220.310 1678.480 ;
        RECT 1215.390 1678.280 1215.710 1678.340 ;
        RECT 1219.990 1678.280 1220.310 1678.340 ;
        RECT 264.110 16.900 264.430 16.960 ;
        RECT 268.710 16.900 269.030 16.960 ;
        RECT 264.110 16.760 269.030 16.900 ;
        RECT 264.110 16.700 264.430 16.760 ;
        RECT 268.710 16.700 269.030 16.760 ;
      LAYER via ;
        RECT 1215.420 1678.280 1215.680 1678.540 ;
        RECT 1220.020 1678.280 1220.280 1678.540 ;
        RECT 264.140 16.700 264.400 16.960 ;
        RECT 268.740 16.700 269.000 16.960 ;
      LAYER met2 ;
        RECT 1220.930 1700.410 1221.210 1704.000 ;
        RECT 1220.080 1700.270 1221.210 1700.410 ;
        RECT 1220.080 1678.570 1220.220 1700.270 ;
        RECT 1220.930 1700.000 1221.210 1700.270 ;
        RECT 1215.420 1678.250 1215.680 1678.570 ;
        RECT 1220.020 1678.250 1220.280 1678.570 ;
        RECT 1215.480 54.245 1215.620 1678.250 ;
        RECT 268.730 53.875 269.010 54.245 ;
        RECT 1215.410 53.875 1215.690 54.245 ;
        RECT 268.800 16.990 268.940 53.875 ;
        RECT 264.140 16.670 264.400 16.990 ;
        RECT 268.740 16.670 269.000 16.990 ;
        RECT 264.200 2.400 264.340 16.670 ;
        RECT 263.990 -4.800 264.550 2.400 ;
      LAYER via2 ;
        RECT 268.730 53.920 269.010 54.200 ;
        RECT 1215.410 53.920 1215.690 54.200 ;
      LAYER met3 ;
        RECT 268.705 54.210 269.035 54.225 ;
        RECT 1215.385 54.210 1215.715 54.225 ;
        RECT 268.705 53.910 1215.715 54.210 ;
        RECT 268.705 53.895 269.035 53.910 ;
        RECT 1215.385 53.895 1215.715 53.910 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1222.290 1678.140 1222.610 1678.200 ;
        RECT 1224.590 1678.140 1224.910 1678.200 ;
        RECT 1222.290 1678.000 1224.910 1678.140 ;
        RECT 1222.290 1677.940 1222.610 1678.000 ;
        RECT 1224.590 1677.940 1224.910 1678.000 ;
      LAYER via ;
        RECT 1222.320 1677.940 1222.580 1678.200 ;
        RECT 1224.620 1677.940 1224.880 1678.200 ;
      LAYER met2 ;
        RECT 1225.990 1700.410 1226.270 1704.000 ;
        RECT 1224.680 1700.270 1226.270 1700.410 ;
        RECT 1224.680 1678.230 1224.820 1700.270 ;
        RECT 1225.990 1700.000 1226.270 1700.270 ;
        RECT 1222.320 1677.910 1222.580 1678.230 ;
        RECT 1224.620 1677.910 1224.880 1678.230 ;
        RECT 1222.380 54.925 1222.520 1677.910 ;
        RECT 282.070 54.555 282.350 54.925 ;
        RECT 1222.310 54.555 1222.590 54.925 ;
        RECT 282.140 2.400 282.280 54.555 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 282.070 54.600 282.350 54.880 ;
        RECT 1222.310 54.600 1222.590 54.880 ;
      LAYER met3 ;
        RECT 282.045 54.890 282.375 54.905 ;
        RECT 1222.285 54.890 1222.615 54.905 ;
        RECT 282.045 54.590 1222.615 54.890 ;
        RECT 282.045 54.575 282.375 54.590 ;
        RECT 1222.285 54.575 1222.615 54.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 0.300 ;
=======
      LAYER met1 ;
        RECT 303.210 51.580 303.530 51.640 ;
        RECT 1230.110 51.580 1230.430 51.640 ;
        RECT 303.210 51.440 1230.430 51.580 ;
        RECT 303.210 51.380 303.530 51.440 ;
        RECT 1230.110 51.380 1230.430 51.440 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 299.990 16.760 303.530 16.900 ;
        RECT 299.990 16.700 300.310 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 303.240 51.380 303.500 51.640 ;
        RECT 1230.140 51.380 1230.400 51.640 ;
        RECT 300.020 16.700 300.280 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 1230.590 1700.410 1230.870 1704.000 ;
        RECT 1230.200 1700.270 1230.870 1700.410 ;
        RECT 1230.200 51.670 1230.340 1700.270 ;
        RECT 1230.590 1700.000 1230.870 1700.270 ;
        RECT 303.240 51.350 303.500 51.670 ;
        RECT 1230.140 51.350 1230.400 51.670 ;
        RECT 303.300 16.990 303.440 51.350 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 0.300 ;
=======
      LAYER met1 ;
        RECT 323.450 51.920 323.770 51.980 ;
        RECT 1236.090 51.920 1236.410 51.980 ;
        RECT 323.450 51.780 1236.410 51.920 ;
        RECT 323.450 51.720 323.770 51.780 ;
        RECT 1236.090 51.720 1236.410 51.780 ;
        RECT 317.930 16.900 318.250 16.960 ;
        RECT 323.450 16.900 323.770 16.960 ;
        RECT 317.930 16.760 323.770 16.900 ;
        RECT 317.930 16.700 318.250 16.760 ;
        RECT 323.450 16.700 323.770 16.760 ;
      LAYER via ;
        RECT 323.480 51.720 323.740 51.980 ;
        RECT 1236.120 51.720 1236.380 51.980 ;
        RECT 317.960 16.700 318.220 16.960 ;
        RECT 323.480 16.700 323.740 16.960 ;
      LAYER met2 ;
        RECT 1235.650 1700.410 1235.930 1704.000 ;
        RECT 1235.650 1700.270 1236.320 1700.410 ;
        RECT 1235.650 1700.000 1235.930 1700.270 ;
        RECT 1236.180 52.010 1236.320 1700.270 ;
        RECT 323.480 51.690 323.740 52.010 ;
        RECT 1236.120 51.690 1236.380 52.010 ;
        RECT 323.540 16.990 323.680 51.690 ;
        RECT 317.960 16.670 318.220 16.990 ;
        RECT 323.480 16.670 323.740 16.990 ;
        RECT 318.020 2.400 318.160 16.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 0.300 ;
=======
      LAYER li1 ;
        RECT 1237.085 1400.205 1237.255 1414.655 ;
        RECT 1237.545 517.905 1237.715 545.955 ;
        RECT 1237.545 434.605 1237.715 469.115 ;
        RECT 1238.005 258.825 1238.175 305.575 ;
        RECT 1238.005 183.685 1238.175 227.715 ;
      LAYER mcon ;
        RECT 1237.085 1414.485 1237.255 1414.655 ;
        RECT 1237.545 545.785 1237.715 545.955 ;
        RECT 1237.545 468.945 1237.715 469.115 ;
        RECT 1238.005 305.405 1238.175 305.575 ;
        RECT 1238.005 227.545 1238.175 227.715 ;
      LAYER met1 ;
        RECT 1237.930 1559.620 1238.250 1559.880 ;
        RECT 1238.020 1559.200 1238.160 1559.620 ;
        RECT 1237.930 1558.940 1238.250 1559.200 ;
        RECT 1237.025 1414.640 1237.315 1414.685 ;
        RECT 1237.470 1414.640 1237.790 1414.700 ;
        RECT 1237.025 1414.500 1237.790 1414.640 ;
        RECT 1237.025 1414.455 1237.315 1414.500 ;
        RECT 1237.470 1414.440 1237.790 1414.500 ;
        RECT 1237.010 1400.360 1237.330 1400.420 ;
        RECT 1236.815 1400.220 1237.330 1400.360 ;
        RECT 1237.010 1400.160 1237.330 1400.220 ;
        RECT 1237.010 1345.620 1237.330 1345.680 ;
        RECT 1237.930 1345.620 1238.250 1345.680 ;
        RECT 1237.010 1345.480 1238.250 1345.620 ;
        RECT 1237.010 1345.420 1237.330 1345.480 ;
        RECT 1237.930 1345.420 1238.250 1345.480 ;
        RECT 1237.470 1283.400 1237.790 1283.460 ;
        RECT 1238.390 1283.400 1238.710 1283.460 ;
        RECT 1237.470 1283.260 1238.710 1283.400 ;
        RECT 1237.470 1283.200 1237.790 1283.260 ;
        RECT 1238.390 1283.200 1238.710 1283.260 ;
        RECT 1237.930 1159.300 1238.250 1159.360 ;
        RECT 1238.390 1159.300 1238.710 1159.360 ;
        RECT 1237.930 1159.160 1238.710 1159.300 ;
        RECT 1237.930 1159.100 1238.250 1159.160 ;
        RECT 1238.390 1159.100 1238.710 1159.160 ;
        RECT 1237.470 1076.680 1237.790 1076.740 ;
        RECT 1237.470 1076.540 1238.160 1076.680 ;
        RECT 1237.470 1076.480 1237.790 1076.540 ;
        RECT 1238.020 1076.400 1238.160 1076.540 ;
        RECT 1237.930 1076.140 1238.250 1076.400 ;
        RECT 1237.470 724.440 1237.790 724.500 ;
        RECT 1238.390 724.440 1238.710 724.500 ;
        RECT 1237.470 724.300 1238.710 724.440 ;
        RECT 1237.470 724.240 1237.790 724.300 ;
        RECT 1238.390 724.240 1238.710 724.300 ;
        RECT 1237.470 572.800 1237.790 572.860 ;
        RECT 1237.930 572.800 1238.250 572.860 ;
        RECT 1237.470 572.660 1238.250 572.800 ;
        RECT 1237.470 572.600 1237.790 572.660 ;
        RECT 1237.930 572.600 1238.250 572.660 ;
        RECT 1237.470 545.940 1237.790 546.000 ;
        RECT 1237.275 545.800 1237.790 545.940 ;
        RECT 1237.470 545.740 1237.790 545.800 ;
        RECT 1237.470 518.060 1237.790 518.120 ;
        RECT 1237.275 517.920 1237.790 518.060 ;
        RECT 1237.470 517.860 1237.790 517.920 ;
        RECT 1237.010 517.380 1237.330 517.440 ;
        RECT 1237.470 517.380 1237.790 517.440 ;
        RECT 1237.010 517.240 1237.790 517.380 ;
        RECT 1237.010 517.180 1237.330 517.240 ;
        RECT 1237.470 517.180 1237.790 517.240 ;
        RECT 1237.470 469.100 1237.790 469.160 ;
        RECT 1237.275 468.960 1237.790 469.100 ;
        RECT 1237.470 468.900 1237.790 468.960 ;
        RECT 1237.485 434.760 1237.775 434.805 ;
        RECT 1237.930 434.760 1238.250 434.820 ;
        RECT 1237.485 434.620 1238.250 434.760 ;
        RECT 1237.485 434.575 1237.775 434.620 ;
        RECT 1237.930 434.560 1238.250 434.620 ;
        RECT 1237.930 305.560 1238.250 305.620 ;
        RECT 1237.735 305.420 1238.250 305.560 ;
        RECT 1237.930 305.360 1238.250 305.420 ;
        RECT 1237.470 258.980 1237.790 259.040 ;
        RECT 1237.945 258.980 1238.235 259.025 ;
        RECT 1237.470 258.840 1238.235 258.980 ;
        RECT 1237.470 258.780 1237.790 258.840 ;
        RECT 1237.945 258.795 1238.235 258.840 ;
        RECT 1237.930 227.700 1238.250 227.760 ;
        RECT 1237.735 227.560 1238.250 227.700 ;
        RECT 1237.930 227.500 1238.250 227.560 ;
        RECT 1237.930 183.840 1238.250 183.900 ;
        RECT 1237.735 183.700 1238.250 183.840 ;
        RECT 1237.930 183.640 1238.250 183.700 ;
        RECT 1237.930 159.020 1238.250 159.080 ;
        RECT 1237.560 158.880 1238.250 159.020 ;
        RECT 1237.560 158.740 1237.700 158.880 ;
        RECT 1237.930 158.820 1238.250 158.880 ;
        RECT 1237.470 158.480 1237.790 158.740 ;
        RECT 337.710 52.260 338.030 52.320 ;
        RECT 1237.470 52.260 1237.790 52.320 ;
        RECT 337.710 52.120 1237.790 52.260 ;
        RECT 337.710 52.060 338.030 52.120 ;
        RECT 1237.470 52.060 1237.790 52.120 ;
      LAYER via ;
        RECT 1237.960 1559.620 1238.220 1559.880 ;
        RECT 1237.960 1558.940 1238.220 1559.200 ;
        RECT 1237.500 1414.440 1237.760 1414.700 ;
        RECT 1237.040 1400.160 1237.300 1400.420 ;
        RECT 1237.040 1345.420 1237.300 1345.680 ;
        RECT 1237.960 1345.420 1238.220 1345.680 ;
        RECT 1237.500 1283.200 1237.760 1283.460 ;
        RECT 1238.420 1283.200 1238.680 1283.460 ;
        RECT 1237.960 1159.100 1238.220 1159.360 ;
        RECT 1238.420 1159.100 1238.680 1159.360 ;
        RECT 1237.500 1076.480 1237.760 1076.740 ;
        RECT 1237.960 1076.140 1238.220 1076.400 ;
        RECT 1237.500 724.240 1237.760 724.500 ;
        RECT 1238.420 724.240 1238.680 724.500 ;
        RECT 1237.500 572.600 1237.760 572.860 ;
        RECT 1237.960 572.600 1238.220 572.860 ;
        RECT 1237.500 545.740 1237.760 546.000 ;
        RECT 1237.500 517.860 1237.760 518.120 ;
        RECT 1237.040 517.180 1237.300 517.440 ;
        RECT 1237.500 517.180 1237.760 517.440 ;
        RECT 1237.500 468.900 1237.760 469.160 ;
        RECT 1237.960 434.560 1238.220 434.820 ;
        RECT 1237.960 305.360 1238.220 305.620 ;
        RECT 1237.500 258.780 1237.760 259.040 ;
        RECT 1237.960 227.500 1238.220 227.760 ;
        RECT 1237.960 183.640 1238.220 183.900 ;
        RECT 1237.960 158.820 1238.220 159.080 ;
        RECT 1237.500 158.480 1237.760 158.740 ;
        RECT 337.740 52.060 338.000 52.320 ;
        RECT 1237.500 52.060 1237.760 52.320 ;
      LAYER met2 ;
        RECT 1240.250 1700.410 1240.530 1704.000 ;
        RECT 1239.860 1700.270 1240.530 1700.410 ;
        RECT 1239.860 1677.970 1240.000 1700.270 ;
        RECT 1240.250 1700.000 1240.530 1700.270 ;
        RECT 1238.020 1677.830 1240.000 1677.970 ;
        RECT 1238.020 1559.910 1238.160 1677.830 ;
        RECT 1237.960 1559.590 1238.220 1559.910 ;
        RECT 1237.960 1558.910 1238.220 1559.230 ;
        RECT 1238.020 1463.090 1238.160 1558.910 ;
        RECT 1237.560 1462.950 1238.160 1463.090 ;
        RECT 1237.560 1462.410 1237.700 1462.950 ;
        RECT 1237.560 1462.270 1238.160 1462.410 ;
        RECT 1238.020 1442.010 1238.160 1462.270 ;
        RECT 1237.560 1441.870 1238.160 1442.010 ;
        RECT 1237.560 1414.730 1237.700 1441.870 ;
        RECT 1237.500 1414.410 1237.760 1414.730 ;
        RECT 1237.040 1400.130 1237.300 1400.450 ;
        RECT 1237.100 1345.710 1237.240 1400.130 ;
        RECT 1237.040 1345.390 1237.300 1345.710 ;
        RECT 1237.960 1345.390 1238.220 1345.710 ;
        RECT 1238.020 1314.170 1238.160 1345.390 ;
        RECT 1237.560 1314.030 1238.160 1314.170 ;
        RECT 1237.560 1283.490 1237.700 1314.030 ;
        RECT 1237.500 1283.170 1237.760 1283.490 ;
        RECT 1238.420 1283.170 1238.680 1283.490 ;
        RECT 1238.480 1159.390 1238.620 1283.170 ;
        RECT 1237.960 1159.070 1238.220 1159.390 ;
        RECT 1238.420 1159.070 1238.680 1159.390 ;
        RECT 1238.020 1104.050 1238.160 1159.070 ;
        RECT 1237.560 1103.910 1238.160 1104.050 ;
        RECT 1237.560 1076.770 1237.700 1103.910 ;
        RECT 1237.500 1076.450 1237.760 1076.770 ;
        RECT 1237.960 1076.110 1238.220 1076.430 ;
        RECT 1238.020 835.450 1238.160 1076.110 ;
        RECT 1237.560 835.310 1238.160 835.450 ;
        RECT 1237.560 834.770 1237.700 835.310 ;
        RECT 1237.560 834.630 1238.160 834.770 ;
        RECT 1238.020 773.685 1238.160 834.630 ;
        RECT 1237.950 773.315 1238.230 773.685 ;
        RECT 1237.950 772.635 1238.230 773.005 ;
        RECT 1238.020 738.890 1238.160 772.635 ;
        RECT 1238.020 738.750 1238.620 738.890 ;
        RECT 1238.480 724.725 1238.620 738.750 ;
        RECT 1237.490 724.355 1237.770 724.725 ;
        RECT 1238.410 724.355 1238.690 724.725 ;
        RECT 1237.500 724.210 1237.760 724.355 ;
        RECT 1238.420 724.210 1238.680 724.355 ;
        RECT 1238.480 699.450 1238.620 724.210 ;
        RECT 1238.020 699.310 1238.620 699.450 ;
        RECT 1238.020 628.845 1238.160 699.310 ;
        RECT 1237.950 628.475 1238.230 628.845 ;
        RECT 1237.950 627.795 1238.230 628.165 ;
        RECT 1238.020 572.890 1238.160 627.795 ;
        RECT 1237.500 572.570 1237.760 572.890 ;
        RECT 1237.960 572.570 1238.220 572.890 ;
        RECT 1237.560 546.030 1237.700 572.570 ;
        RECT 1237.500 545.710 1237.760 546.030 ;
        RECT 1237.500 517.830 1237.760 518.150 ;
        RECT 1237.560 517.470 1237.700 517.830 ;
        RECT 1237.040 517.150 1237.300 517.470 ;
        RECT 1237.500 517.150 1237.760 517.470 ;
        RECT 1237.100 475.730 1237.240 517.150 ;
        RECT 1237.100 475.590 1237.700 475.730 ;
        RECT 1237.560 469.190 1237.700 475.590 ;
        RECT 1237.500 468.870 1237.760 469.190 ;
        RECT 1237.960 434.530 1238.220 434.850 ;
        RECT 1238.020 305.650 1238.160 434.530 ;
        RECT 1237.960 305.330 1238.220 305.650 ;
        RECT 1237.500 258.750 1237.760 259.070 ;
        RECT 1237.560 235.010 1237.700 258.750 ;
        RECT 1237.560 234.870 1238.160 235.010 ;
        RECT 1238.020 227.790 1238.160 234.870 ;
        RECT 1237.960 227.470 1238.220 227.790 ;
        RECT 1237.960 183.610 1238.220 183.930 ;
        RECT 1238.020 159.110 1238.160 183.610 ;
        RECT 1237.960 158.790 1238.220 159.110 ;
        RECT 1237.500 158.450 1237.760 158.770 ;
        RECT 1237.560 52.350 1237.700 158.450 ;
        RECT 337.740 52.030 338.000 52.350 ;
        RECT 1237.500 52.030 1237.760 52.350 ;
        RECT 337.800 17.410 337.940 52.030 ;
        RECT 335.960 17.270 337.940 17.410 ;
        RECT 335.960 2.400 336.100 17.270 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 1237.950 773.360 1238.230 773.640 ;
        RECT 1237.950 772.680 1238.230 772.960 ;
        RECT 1237.490 724.400 1237.770 724.680 ;
        RECT 1238.410 724.400 1238.690 724.680 ;
        RECT 1237.950 628.520 1238.230 628.800 ;
        RECT 1237.950 627.840 1238.230 628.120 ;
      LAYER met3 ;
        RECT 1237.925 773.650 1238.255 773.665 ;
        RECT 1237.710 773.335 1238.255 773.650 ;
        RECT 1237.710 772.985 1238.010 773.335 ;
        RECT 1237.710 772.670 1238.255 772.985 ;
        RECT 1237.925 772.655 1238.255 772.670 ;
        RECT 1237.465 724.690 1237.795 724.705 ;
        RECT 1238.385 724.690 1238.715 724.705 ;
        RECT 1237.465 724.390 1238.715 724.690 ;
        RECT 1237.465 724.375 1237.795 724.390 ;
        RECT 1238.385 724.375 1238.715 724.390 ;
        RECT 1237.925 628.810 1238.255 628.825 ;
        RECT 1237.710 628.495 1238.255 628.810 ;
        RECT 1237.710 628.145 1238.010 628.495 ;
        RECT 1237.710 627.830 1238.255 628.145 ;
        RECT 1237.925 627.815 1238.255 627.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 0.300 ;
=======
      LAYER met1 ;
        RECT 358.410 59.060 358.730 59.120 ;
        RECT 1244.370 59.060 1244.690 59.120 ;
        RECT 358.410 58.920 1244.690 59.060 ;
        RECT 358.410 58.860 358.730 58.920 ;
        RECT 1244.370 58.860 1244.690 58.920 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 358.410 16.900 358.730 16.960 ;
        RECT 353.350 16.760 358.730 16.900 ;
        RECT 353.350 16.700 353.670 16.760 ;
        RECT 358.410 16.700 358.730 16.760 ;
      LAYER via ;
        RECT 358.440 58.860 358.700 59.120 ;
        RECT 1244.400 58.860 1244.660 59.120 ;
        RECT 353.380 16.700 353.640 16.960 ;
        RECT 358.440 16.700 358.700 16.960 ;
      LAYER met2 ;
        RECT 1245.310 1700.410 1245.590 1704.000 ;
        RECT 1244.460 1700.270 1245.590 1700.410 ;
        RECT 1244.460 59.150 1244.600 1700.270 ;
        RECT 1245.310 1700.000 1245.590 1700.270 ;
        RECT 358.440 58.830 358.700 59.150 ;
        RECT 1244.400 58.830 1244.660 59.150 ;
        RECT 358.500 16.990 358.640 58.830 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 358.440 16.670 358.700 16.990 ;
        RECT 353.440 2.400 353.580 16.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 0.300 ;
=======
      LAYER li1 ;
        RECT 1249.965 1655.885 1250.135 1683.595 ;
        RECT 1249.965 1331.865 1250.135 1379.975 ;
        RECT 1249.965 1193.825 1250.135 1259.275 ;
        RECT 1250.425 1048.985 1250.595 1097.095 ;
        RECT 1249.965 869.465 1250.135 917.575 ;
        RECT 1250.425 620.925 1250.595 669.375 ;
        RECT 1249.965 476.085 1250.135 524.195 ;
        RECT 1249.965 379.525 1250.135 427.635 ;
        RECT 1249.965 59.245 1250.135 62.475 ;
      LAYER mcon ;
        RECT 1249.965 1683.425 1250.135 1683.595 ;
        RECT 1249.965 1379.805 1250.135 1379.975 ;
        RECT 1249.965 1259.105 1250.135 1259.275 ;
        RECT 1250.425 1096.925 1250.595 1097.095 ;
        RECT 1249.965 917.405 1250.135 917.575 ;
        RECT 1250.425 669.205 1250.595 669.375 ;
        RECT 1249.965 524.025 1250.135 524.195 ;
        RECT 1249.965 427.465 1250.135 427.635 ;
        RECT 1249.965 62.305 1250.135 62.475 ;
      LAYER met1 ;
        RECT 1249.890 1691.060 1250.210 1691.120 ;
        RECT 1250.350 1691.060 1250.670 1691.120 ;
        RECT 1249.890 1690.920 1250.670 1691.060 ;
        RECT 1249.890 1690.860 1250.210 1690.920 ;
        RECT 1250.350 1690.860 1250.670 1690.920 ;
        RECT 1249.905 1683.580 1250.195 1683.625 ;
        RECT 1250.350 1683.580 1250.670 1683.640 ;
        RECT 1249.905 1683.440 1250.670 1683.580 ;
        RECT 1249.905 1683.395 1250.195 1683.440 ;
        RECT 1250.350 1683.380 1250.670 1683.440 ;
        RECT 1249.905 1656.040 1250.195 1656.085 ;
        RECT 1250.350 1656.040 1250.670 1656.100 ;
        RECT 1249.905 1655.900 1250.670 1656.040 ;
        RECT 1249.905 1655.855 1250.195 1655.900 ;
        RECT 1250.350 1655.840 1250.670 1655.900 ;
        RECT 1249.890 1545.880 1250.210 1545.940 ;
        RECT 1250.810 1545.880 1251.130 1545.940 ;
        RECT 1249.890 1545.740 1251.130 1545.880 ;
        RECT 1249.890 1545.680 1250.210 1545.740 ;
        RECT 1250.810 1545.680 1251.130 1545.740 ;
        RECT 1248.050 1393.560 1248.370 1393.620 ;
        RECT 1249.890 1393.560 1250.210 1393.620 ;
        RECT 1248.050 1393.420 1250.210 1393.560 ;
        RECT 1248.050 1393.360 1248.370 1393.420 ;
        RECT 1249.890 1393.360 1250.210 1393.420 ;
        RECT 1249.890 1379.960 1250.210 1380.020 ;
        RECT 1249.695 1379.820 1250.210 1379.960 ;
        RECT 1249.890 1379.760 1250.210 1379.820 ;
        RECT 1249.905 1332.020 1250.195 1332.065 ;
        RECT 1250.350 1332.020 1250.670 1332.080 ;
        RECT 1249.905 1331.880 1250.670 1332.020 ;
        RECT 1249.905 1331.835 1250.195 1331.880 ;
        RECT 1250.350 1331.820 1250.670 1331.880 ;
        RECT 1249.905 1259.260 1250.195 1259.305 ;
        RECT 1251.270 1259.260 1251.590 1259.320 ;
        RECT 1249.905 1259.120 1251.590 1259.260 ;
        RECT 1249.905 1259.075 1250.195 1259.120 ;
        RECT 1251.270 1259.060 1251.590 1259.120 ;
        RECT 1249.905 1193.980 1250.195 1194.025 ;
        RECT 1250.350 1193.980 1250.670 1194.040 ;
        RECT 1249.905 1193.840 1250.670 1193.980 ;
        RECT 1249.905 1193.795 1250.195 1193.840 ;
        RECT 1250.350 1193.780 1250.670 1193.840 ;
        RECT 1249.890 1152.500 1250.210 1152.560 ;
        RECT 1250.350 1152.500 1250.670 1152.560 ;
        RECT 1249.890 1152.360 1250.670 1152.500 ;
        RECT 1249.890 1152.300 1250.210 1152.360 ;
        RECT 1250.350 1152.300 1250.670 1152.360 ;
        RECT 1249.890 1104.220 1250.210 1104.280 ;
        RECT 1250.810 1104.220 1251.130 1104.280 ;
        RECT 1249.890 1104.080 1251.130 1104.220 ;
        RECT 1249.890 1104.020 1250.210 1104.080 ;
        RECT 1250.810 1104.020 1251.130 1104.080 ;
        RECT 1250.365 1097.080 1250.655 1097.125 ;
        RECT 1250.810 1097.080 1251.130 1097.140 ;
        RECT 1250.365 1096.940 1251.130 1097.080 ;
        RECT 1250.365 1096.895 1250.655 1096.940 ;
        RECT 1250.810 1096.880 1251.130 1096.940 ;
        RECT 1250.350 1049.140 1250.670 1049.200 ;
        RECT 1250.155 1049.000 1250.670 1049.140 ;
        RECT 1250.350 1048.940 1250.670 1049.000 ;
        RECT 1249.890 979.440 1250.210 979.500 ;
        RECT 1250.810 979.440 1251.130 979.500 ;
        RECT 1249.890 979.300 1251.130 979.440 ;
        RECT 1249.890 979.240 1250.210 979.300 ;
        RECT 1250.810 979.240 1251.130 979.300 ;
        RECT 1249.890 931.640 1250.210 931.900 ;
        RECT 1249.980 931.160 1250.120 931.640 ;
        RECT 1250.350 931.160 1250.670 931.220 ;
        RECT 1249.980 931.020 1250.670 931.160 ;
        RECT 1250.350 930.960 1250.670 931.020 ;
        RECT 1249.905 917.560 1250.195 917.605 ;
        RECT 1250.350 917.560 1250.670 917.620 ;
        RECT 1249.905 917.420 1250.670 917.560 ;
        RECT 1249.905 917.375 1250.195 917.420 ;
        RECT 1250.350 917.360 1250.670 917.420 ;
        RECT 1249.890 869.620 1250.210 869.680 ;
        RECT 1249.695 869.480 1250.210 869.620 ;
        RECT 1249.890 869.420 1250.210 869.480 ;
        RECT 1250.350 669.360 1250.670 669.420 ;
        RECT 1250.155 669.220 1250.670 669.360 ;
        RECT 1250.350 669.160 1250.670 669.220 ;
        RECT 1250.350 621.080 1250.670 621.140 ;
        RECT 1250.155 620.940 1250.670 621.080 ;
        RECT 1250.350 620.880 1250.670 620.940 ;
        RECT 1249.890 572.800 1250.210 572.860 ;
        RECT 1250.350 572.800 1250.670 572.860 ;
        RECT 1249.890 572.660 1250.670 572.800 ;
        RECT 1249.890 572.600 1250.210 572.660 ;
        RECT 1250.350 572.600 1250.670 572.660 ;
        RECT 1249.890 531.320 1250.210 531.380 ;
        RECT 1250.350 531.320 1250.670 531.380 ;
        RECT 1249.890 531.180 1250.670 531.320 ;
        RECT 1249.890 531.120 1250.210 531.180 ;
        RECT 1250.350 531.120 1250.670 531.180 ;
        RECT 1249.890 524.180 1250.210 524.240 ;
        RECT 1249.695 524.040 1250.210 524.180 ;
        RECT 1249.890 523.980 1250.210 524.040 ;
        RECT 1249.890 476.240 1250.210 476.300 ;
        RECT 1249.695 476.100 1250.210 476.240 ;
        RECT 1249.890 476.040 1250.210 476.100 ;
        RECT 1249.890 427.620 1250.210 427.680 ;
        RECT 1249.695 427.480 1250.210 427.620 ;
        RECT 1249.890 427.420 1250.210 427.480 ;
        RECT 1249.890 379.680 1250.210 379.740 ;
        RECT 1249.695 379.540 1250.210 379.680 ;
        RECT 1249.890 379.480 1250.210 379.540 ;
        RECT 1250.350 331.060 1250.670 331.120 ;
        RECT 1249.980 330.920 1250.670 331.060 ;
        RECT 1249.980 330.780 1250.120 330.920 ;
        RECT 1250.350 330.860 1250.670 330.920 ;
        RECT 1249.890 330.520 1250.210 330.780 ;
        RECT 1249.890 241.640 1250.210 241.700 ;
        RECT 1250.350 241.640 1250.670 241.700 ;
        RECT 1249.890 241.500 1250.670 241.640 ;
        RECT 1249.890 241.440 1250.210 241.500 ;
        RECT 1250.350 241.440 1250.670 241.500 ;
        RECT 1250.350 137.940 1250.670 138.000 ;
        RECT 1249.980 137.800 1250.670 137.940 ;
        RECT 1249.980 137.660 1250.120 137.800 ;
        RECT 1250.350 137.740 1250.670 137.800 ;
        RECT 1249.890 137.400 1250.210 137.660 ;
        RECT 1249.890 62.460 1250.210 62.520 ;
        RECT 1249.695 62.320 1250.210 62.460 ;
        RECT 1249.890 62.260 1250.210 62.320 ;
        RECT 372.210 59.400 372.530 59.460 ;
        RECT 1249.905 59.400 1250.195 59.445 ;
        RECT 372.210 59.260 1250.195 59.400 ;
        RECT 372.210 59.200 372.530 59.260 ;
        RECT 1249.905 59.215 1250.195 59.260 ;
      LAYER via ;
        RECT 1249.920 1690.860 1250.180 1691.120 ;
        RECT 1250.380 1690.860 1250.640 1691.120 ;
        RECT 1250.380 1683.380 1250.640 1683.640 ;
        RECT 1250.380 1655.840 1250.640 1656.100 ;
        RECT 1249.920 1545.680 1250.180 1545.940 ;
        RECT 1250.840 1545.680 1251.100 1545.940 ;
        RECT 1248.080 1393.360 1248.340 1393.620 ;
        RECT 1249.920 1393.360 1250.180 1393.620 ;
        RECT 1249.920 1379.760 1250.180 1380.020 ;
        RECT 1250.380 1331.820 1250.640 1332.080 ;
        RECT 1251.300 1259.060 1251.560 1259.320 ;
        RECT 1250.380 1193.780 1250.640 1194.040 ;
        RECT 1249.920 1152.300 1250.180 1152.560 ;
        RECT 1250.380 1152.300 1250.640 1152.560 ;
        RECT 1249.920 1104.020 1250.180 1104.280 ;
        RECT 1250.840 1104.020 1251.100 1104.280 ;
        RECT 1250.840 1096.880 1251.100 1097.140 ;
        RECT 1250.380 1048.940 1250.640 1049.200 ;
        RECT 1249.920 979.240 1250.180 979.500 ;
        RECT 1250.840 979.240 1251.100 979.500 ;
        RECT 1249.920 931.640 1250.180 931.900 ;
        RECT 1250.380 930.960 1250.640 931.220 ;
        RECT 1250.380 917.360 1250.640 917.620 ;
        RECT 1249.920 869.420 1250.180 869.680 ;
        RECT 1250.380 669.160 1250.640 669.420 ;
        RECT 1250.380 620.880 1250.640 621.140 ;
        RECT 1249.920 572.600 1250.180 572.860 ;
        RECT 1250.380 572.600 1250.640 572.860 ;
        RECT 1249.920 531.120 1250.180 531.380 ;
        RECT 1250.380 531.120 1250.640 531.380 ;
        RECT 1249.920 523.980 1250.180 524.240 ;
        RECT 1249.920 476.040 1250.180 476.300 ;
        RECT 1249.920 427.420 1250.180 427.680 ;
        RECT 1249.920 379.480 1250.180 379.740 ;
        RECT 1250.380 330.860 1250.640 331.120 ;
        RECT 1249.920 330.520 1250.180 330.780 ;
        RECT 1249.920 241.440 1250.180 241.700 ;
        RECT 1250.380 241.440 1250.640 241.700 ;
        RECT 1250.380 137.740 1250.640 138.000 ;
        RECT 1249.920 137.400 1250.180 137.660 ;
        RECT 1249.920 62.260 1250.180 62.520 ;
        RECT 372.240 59.200 372.500 59.460 ;
      LAYER met2 ;
        RECT 1249.910 1700.000 1250.190 1704.000 ;
        RECT 1249.980 1691.150 1250.120 1700.000 ;
        RECT 1249.920 1690.830 1250.180 1691.150 ;
        RECT 1250.380 1690.830 1250.640 1691.150 ;
        RECT 1250.440 1683.670 1250.580 1690.830 ;
        RECT 1250.380 1683.350 1250.640 1683.670 ;
        RECT 1250.380 1655.810 1250.640 1656.130 ;
        RECT 1250.440 1593.650 1250.580 1655.810 ;
        RECT 1249.980 1593.510 1250.580 1593.650 ;
        RECT 1249.980 1545.970 1250.120 1593.510 ;
        RECT 1249.920 1545.650 1250.180 1545.970 ;
        RECT 1250.840 1545.650 1251.100 1545.970 ;
        RECT 1250.900 1428.525 1251.040 1545.650 ;
        RECT 1248.070 1428.155 1248.350 1428.525 ;
        RECT 1250.830 1428.155 1251.110 1428.525 ;
        RECT 1248.140 1393.650 1248.280 1428.155 ;
        RECT 1248.080 1393.330 1248.340 1393.650 ;
        RECT 1249.920 1393.330 1250.180 1393.650 ;
        RECT 1249.980 1380.050 1250.120 1393.330 ;
        RECT 1249.920 1379.730 1250.180 1380.050 ;
        RECT 1250.380 1331.790 1250.640 1332.110 ;
        RECT 1250.440 1307.370 1250.580 1331.790 ;
        RECT 1250.440 1307.230 1251.040 1307.370 ;
        RECT 1250.900 1283.570 1251.040 1307.230 ;
        RECT 1250.900 1283.430 1251.500 1283.570 ;
        RECT 1251.360 1259.350 1251.500 1283.430 ;
        RECT 1251.300 1259.030 1251.560 1259.350 ;
        RECT 1250.380 1193.750 1250.640 1194.070 ;
        RECT 1250.440 1152.590 1250.580 1193.750 ;
        RECT 1249.920 1152.270 1250.180 1152.590 ;
        RECT 1250.380 1152.270 1250.640 1152.590 ;
        RECT 1249.980 1104.310 1250.120 1152.270 ;
        RECT 1249.920 1103.990 1250.180 1104.310 ;
        RECT 1250.840 1103.990 1251.100 1104.310 ;
        RECT 1250.900 1097.170 1251.040 1103.990 ;
        RECT 1250.840 1096.850 1251.100 1097.170 ;
        RECT 1250.380 1048.910 1250.640 1049.230 ;
        RECT 1250.440 1014.405 1250.580 1048.910 ;
        RECT 1250.370 1014.035 1250.650 1014.405 ;
        RECT 1250.830 1013.355 1251.110 1013.725 ;
        RECT 1250.900 979.530 1251.040 1013.355 ;
        RECT 1249.920 979.210 1250.180 979.530 ;
        RECT 1250.840 979.210 1251.100 979.530 ;
        RECT 1249.980 931.930 1250.120 979.210 ;
        RECT 1249.920 931.610 1250.180 931.930 ;
        RECT 1250.380 930.930 1250.640 931.250 ;
        RECT 1250.440 917.650 1250.580 930.930 ;
        RECT 1250.380 917.330 1250.640 917.650 ;
        RECT 1249.920 869.390 1250.180 869.710 ;
        RECT 1249.980 845.650 1250.120 869.390 ;
        RECT 1249.980 845.510 1250.580 845.650 ;
        RECT 1250.440 773.685 1250.580 845.510 ;
        RECT 1250.370 773.315 1250.650 773.685 ;
        RECT 1249.910 772.635 1250.190 773.005 ;
        RECT 1249.980 748.410 1250.120 772.635 ;
        RECT 1249.980 748.270 1250.580 748.410 ;
        RECT 1250.440 669.450 1250.580 748.270 ;
        RECT 1250.380 669.130 1250.640 669.450 ;
        RECT 1250.380 620.850 1250.640 621.170 ;
        RECT 1250.440 572.890 1250.580 620.850 ;
        RECT 1249.920 572.570 1250.180 572.890 ;
        RECT 1250.380 572.570 1250.640 572.890 ;
        RECT 1249.980 555.970 1250.120 572.570 ;
        RECT 1249.980 555.830 1250.580 555.970 ;
        RECT 1250.440 531.410 1250.580 555.830 ;
        RECT 1249.920 531.090 1250.180 531.410 ;
        RECT 1250.380 531.090 1250.640 531.410 ;
        RECT 1249.980 524.270 1250.120 531.090 ;
        RECT 1249.920 523.950 1250.180 524.270 ;
        RECT 1249.920 476.010 1250.180 476.330 ;
        RECT 1249.980 435.725 1250.120 476.010 ;
        RECT 1249.910 435.355 1250.190 435.725 ;
        RECT 1249.910 434.675 1250.190 435.045 ;
        RECT 1249.980 427.710 1250.120 434.675 ;
        RECT 1249.920 427.390 1250.180 427.710 ;
        RECT 1249.920 379.450 1250.180 379.770 ;
        RECT 1249.980 355.370 1250.120 379.450 ;
        RECT 1249.980 355.230 1251.040 355.370 ;
        RECT 1250.900 351.800 1251.040 355.230 ;
        RECT 1250.440 351.660 1251.040 351.800 ;
        RECT 1250.440 331.150 1250.580 351.660 ;
        RECT 1250.380 330.830 1250.640 331.150 ;
        RECT 1249.920 330.490 1250.180 330.810 ;
        RECT 1249.980 241.730 1250.120 330.490 ;
        RECT 1249.920 241.410 1250.180 241.730 ;
        RECT 1250.380 241.410 1250.640 241.730 ;
        RECT 1250.440 186.730 1250.580 241.410 ;
        RECT 1249.980 186.590 1250.580 186.730 ;
        RECT 1249.980 162.930 1250.120 186.590 ;
        RECT 1249.980 162.790 1250.580 162.930 ;
        RECT 1250.440 138.030 1250.580 162.790 ;
        RECT 1250.380 137.710 1250.640 138.030 ;
        RECT 1249.920 137.370 1250.180 137.690 ;
        RECT 1249.980 62.550 1250.120 137.370 ;
        RECT 1249.920 62.230 1250.180 62.550 ;
        RECT 372.240 59.170 372.500 59.490 ;
        RECT 372.300 17.410 372.440 59.170 ;
        RECT 371.380 17.270 372.440 17.410 ;
        RECT 371.380 2.400 371.520 17.270 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 1248.070 1428.200 1248.350 1428.480 ;
        RECT 1250.830 1428.200 1251.110 1428.480 ;
        RECT 1250.370 1014.080 1250.650 1014.360 ;
        RECT 1250.830 1013.400 1251.110 1013.680 ;
        RECT 1250.370 773.360 1250.650 773.640 ;
        RECT 1249.910 772.680 1250.190 772.960 ;
        RECT 1249.910 435.400 1250.190 435.680 ;
        RECT 1249.910 434.720 1250.190 435.000 ;
      LAYER met3 ;
        RECT 1248.045 1428.490 1248.375 1428.505 ;
        RECT 1250.805 1428.490 1251.135 1428.505 ;
        RECT 1248.045 1428.190 1251.135 1428.490 ;
        RECT 1248.045 1428.175 1248.375 1428.190 ;
        RECT 1250.805 1428.175 1251.135 1428.190 ;
        RECT 1250.345 1014.370 1250.675 1014.385 ;
        RECT 1250.345 1014.055 1250.890 1014.370 ;
        RECT 1250.590 1013.705 1250.890 1014.055 ;
        RECT 1250.590 1013.390 1251.135 1013.705 ;
        RECT 1250.805 1013.375 1251.135 1013.390 ;
        RECT 1250.345 773.650 1250.675 773.665 ;
        RECT 1249.670 773.350 1250.675 773.650 ;
        RECT 1249.670 772.985 1249.970 773.350 ;
        RECT 1250.345 773.335 1250.675 773.350 ;
        RECT 1249.670 772.670 1250.215 772.985 ;
        RECT 1249.885 772.655 1250.215 772.670 ;
        RECT 1249.885 435.690 1250.215 435.705 ;
        RECT 1249.670 435.375 1250.215 435.690 ;
        RECT 1249.670 435.025 1249.970 435.375 ;
        RECT 1249.670 434.710 1250.215 435.025 ;
        RECT 1249.885 434.695 1250.215 434.710 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 0.300 ;
=======
      LAYER li1 ;
        RECT 1251.345 1538.925 1251.515 1587.035 ;
        RECT 1251.345 1386.945 1251.515 1414.995 ;
        RECT 1251.345 1297.185 1251.515 1345.295 ;
        RECT 1251.345 1104.065 1251.515 1140.955 ;
        RECT 1251.805 565.845 1251.975 590.155 ;
        RECT 1251.345 331.245 1251.515 379.355 ;
        RECT 1251.345 59.585 1251.515 96.475 ;
      LAYER mcon ;
        RECT 1251.345 1586.865 1251.515 1587.035 ;
        RECT 1251.345 1414.825 1251.515 1414.995 ;
        RECT 1251.345 1345.125 1251.515 1345.295 ;
        RECT 1251.345 1140.785 1251.515 1140.955 ;
        RECT 1251.805 589.985 1251.975 590.155 ;
        RECT 1251.345 379.185 1251.515 379.355 ;
        RECT 1251.345 96.305 1251.515 96.475 ;
      LAYER met1 ;
        RECT 1251.270 1587.020 1251.590 1587.080 ;
        RECT 1251.075 1586.880 1251.590 1587.020 ;
        RECT 1251.270 1586.820 1251.590 1586.880 ;
        RECT 1251.285 1539.080 1251.575 1539.125 ;
        RECT 1251.730 1539.080 1252.050 1539.140 ;
        RECT 1251.285 1538.940 1252.050 1539.080 ;
        RECT 1251.285 1538.895 1251.575 1538.940 ;
        RECT 1251.730 1538.880 1252.050 1538.940 ;
        RECT 1251.270 1414.980 1251.590 1415.040 ;
        RECT 1251.075 1414.840 1251.590 1414.980 ;
        RECT 1251.270 1414.780 1251.590 1414.840 ;
        RECT 1251.270 1387.100 1251.590 1387.160 ;
        RECT 1251.075 1386.960 1251.590 1387.100 ;
        RECT 1251.270 1386.900 1251.590 1386.960 ;
        RECT 1251.270 1345.280 1251.590 1345.340 ;
        RECT 1251.075 1345.140 1251.590 1345.280 ;
        RECT 1251.270 1345.080 1251.590 1345.140 ;
        RECT 1251.285 1297.340 1251.575 1297.385 ;
        RECT 1252.190 1297.340 1252.510 1297.400 ;
        RECT 1251.285 1297.200 1252.510 1297.340 ;
        RECT 1251.285 1297.155 1251.575 1297.200 ;
        RECT 1252.190 1297.140 1252.510 1297.200 ;
        RECT 1251.270 1249.060 1251.590 1249.120 ;
        RECT 1252.190 1249.060 1252.510 1249.120 ;
        RECT 1251.270 1248.920 1252.510 1249.060 ;
        RECT 1251.270 1248.860 1251.590 1248.920 ;
        RECT 1252.190 1248.860 1252.510 1248.920 ;
        RECT 1251.270 1207.380 1251.590 1207.640 ;
        RECT 1251.360 1207.240 1251.500 1207.380 ;
        RECT 1251.730 1207.240 1252.050 1207.300 ;
        RECT 1251.360 1207.100 1252.050 1207.240 ;
        RECT 1251.730 1207.040 1252.050 1207.100 ;
        RECT 1251.270 1152.500 1251.590 1152.560 ;
        RECT 1252.190 1152.500 1252.510 1152.560 ;
        RECT 1251.270 1152.360 1252.510 1152.500 ;
        RECT 1251.270 1152.300 1251.590 1152.360 ;
        RECT 1252.190 1152.300 1252.510 1152.360 ;
        RECT 1251.270 1140.940 1251.590 1141.000 ;
        RECT 1251.075 1140.800 1251.590 1140.940 ;
        RECT 1251.270 1140.740 1251.590 1140.800 ;
        RECT 1251.285 1104.220 1251.575 1104.265 ;
        RECT 1252.190 1104.220 1252.510 1104.280 ;
        RECT 1251.285 1104.080 1252.510 1104.220 ;
        RECT 1251.285 1104.035 1251.575 1104.080 ;
        RECT 1252.190 1104.020 1252.510 1104.080 ;
        RECT 1252.190 1097.080 1252.510 1097.140 ;
        RECT 1253.110 1097.080 1253.430 1097.140 ;
        RECT 1252.190 1096.940 1253.430 1097.080 ;
        RECT 1252.190 1096.880 1252.510 1096.940 ;
        RECT 1253.110 1096.880 1253.430 1096.940 ;
        RECT 1251.730 1014.800 1252.050 1014.860 ;
        RECT 1251.360 1014.660 1252.050 1014.800 ;
        RECT 1251.360 1014.520 1251.500 1014.660 ;
        RECT 1251.730 1014.600 1252.050 1014.660 ;
        RECT 1251.270 1014.260 1251.590 1014.520 ;
        RECT 1251.270 979.920 1251.590 980.180 ;
        RECT 1251.360 979.500 1251.500 979.920 ;
        RECT 1251.270 979.240 1251.590 979.500 ;
        RECT 1251.270 931.640 1251.590 931.900 ;
        RECT 1251.360 931.160 1251.500 931.640 ;
        RECT 1251.730 931.160 1252.050 931.220 ;
        RECT 1251.360 931.020 1252.050 931.160 ;
        RECT 1251.730 930.960 1252.050 931.020 ;
        RECT 1251.270 869.620 1251.590 869.680 ;
        RECT 1252.190 869.620 1252.510 869.680 ;
        RECT 1251.270 869.480 1252.510 869.620 ;
        RECT 1251.270 869.420 1251.590 869.480 ;
        RECT 1252.190 869.420 1252.510 869.480 ;
        RECT 1251.730 786.660 1252.050 786.720 ;
        RECT 1251.360 786.520 1252.050 786.660 ;
        RECT 1251.360 786.380 1251.500 786.520 ;
        RECT 1251.730 786.460 1252.050 786.520 ;
        RECT 1251.270 786.120 1251.590 786.380 ;
        RECT 1251.270 738.180 1251.590 738.440 ;
        RECT 1251.360 738.040 1251.500 738.180 ;
        RECT 1251.730 738.040 1252.050 738.100 ;
        RECT 1251.360 737.900 1252.050 738.040 ;
        RECT 1251.730 737.840 1252.050 737.900 ;
        RECT 1251.270 676.160 1251.590 676.220 ;
        RECT 1252.190 676.160 1252.510 676.220 ;
        RECT 1251.270 676.020 1252.510 676.160 ;
        RECT 1251.270 675.960 1251.590 676.020 ;
        RECT 1252.190 675.960 1252.510 676.020 ;
        RECT 1251.730 590.140 1252.050 590.200 ;
        RECT 1251.535 590.000 1252.050 590.140 ;
        RECT 1251.730 589.940 1252.050 590.000 ;
        RECT 1251.745 566.000 1252.035 566.045 ;
        RECT 1252.190 566.000 1252.510 566.060 ;
        RECT 1251.745 565.860 1252.510 566.000 ;
        RECT 1251.745 565.815 1252.035 565.860 ;
        RECT 1252.190 565.800 1252.510 565.860 ;
        RECT 1251.270 524.520 1251.590 524.580 ;
        RECT 1252.190 524.520 1252.510 524.580 ;
        RECT 1251.270 524.380 1252.510 524.520 ;
        RECT 1251.270 524.320 1251.590 524.380 ;
        RECT 1252.190 524.320 1252.510 524.380 ;
        RECT 1250.810 469.440 1251.130 469.500 ;
        RECT 1251.730 469.440 1252.050 469.500 ;
        RECT 1250.810 469.300 1252.050 469.440 ;
        RECT 1250.810 469.240 1251.130 469.300 ;
        RECT 1251.730 469.240 1252.050 469.300 ;
        RECT 1251.270 379.340 1251.590 379.400 ;
        RECT 1251.075 379.200 1251.590 379.340 ;
        RECT 1251.270 379.140 1251.590 379.200 ;
        RECT 1251.270 331.400 1251.590 331.460 ;
        RECT 1251.075 331.260 1251.590 331.400 ;
        RECT 1251.270 331.200 1251.590 331.260 ;
        RECT 1251.730 159.020 1252.050 159.080 ;
        RECT 1251.360 158.880 1252.050 159.020 ;
        RECT 1251.360 158.740 1251.500 158.880 ;
        RECT 1251.730 158.820 1252.050 158.880 ;
        RECT 1251.270 158.480 1251.590 158.740 ;
        RECT 1251.270 96.460 1251.590 96.520 ;
        RECT 1251.075 96.320 1251.590 96.460 ;
        RECT 1251.270 96.260 1251.590 96.320 ;
        RECT 392.910 59.740 393.230 59.800 ;
        RECT 1251.285 59.740 1251.575 59.785 ;
        RECT 392.910 59.600 1251.575 59.740 ;
        RECT 392.910 59.540 393.230 59.600 ;
        RECT 1251.285 59.555 1251.575 59.600 ;
        RECT 389.230 16.900 389.550 16.960 ;
        RECT 392.910 16.900 393.230 16.960 ;
        RECT 389.230 16.760 393.230 16.900 ;
        RECT 389.230 16.700 389.550 16.760 ;
        RECT 392.910 16.700 393.230 16.760 ;
      LAYER via ;
        RECT 1251.300 1586.820 1251.560 1587.080 ;
        RECT 1251.760 1538.880 1252.020 1539.140 ;
        RECT 1251.300 1414.780 1251.560 1415.040 ;
        RECT 1251.300 1386.900 1251.560 1387.160 ;
        RECT 1251.300 1345.080 1251.560 1345.340 ;
        RECT 1252.220 1297.140 1252.480 1297.400 ;
        RECT 1251.300 1248.860 1251.560 1249.120 ;
        RECT 1252.220 1248.860 1252.480 1249.120 ;
        RECT 1251.300 1207.380 1251.560 1207.640 ;
        RECT 1251.760 1207.040 1252.020 1207.300 ;
        RECT 1251.300 1152.300 1251.560 1152.560 ;
        RECT 1252.220 1152.300 1252.480 1152.560 ;
        RECT 1251.300 1140.740 1251.560 1141.000 ;
        RECT 1252.220 1104.020 1252.480 1104.280 ;
        RECT 1252.220 1096.880 1252.480 1097.140 ;
        RECT 1253.140 1096.880 1253.400 1097.140 ;
        RECT 1251.760 1014.600 1252.020 1014.860 ;
        RECT 1251.300 1014.260 1251.560 1014.520 ;
        RECT 1251.300 979.920 1251.560 980.180 ;
        RECT 1251.300 979.240 1251.560 979.500 ;
        RECT 1251.300 931.640 1251.560 931.900 ;
        RECT 1251.760 930.960 1252.020 931.220 ;
        RECT 1251.300 869.420 1251.560 869.680 ;
        RECT 1252.220 869.420 1252.480 869.680 ;
        RECT 1251.760 786.460 1252.020 786.720 ;
        RECT 1251.300 786.120 1251.560 786.380 ;
        RECT 1251.300 738.180 1251.560 738.440 ;
        RECT 1251.760 737.840 1252.020 738.100 ;
        RECT 1251.300 675.960 1251.560 676.220 ;
        RECT 1252.220 675.960 1252.480 676.220 ;
        RECT 1251.760 589.940 1252.020 590.200 ;
        RECT 1252.220 565.800 1252.480 566.060 ;
        RECT 1251.300 524.320 1251.560 524.580 ;
        RECT 1252.220 524.320 1252.480 524.580 ;
        RECT 1250.840 469.240 1251.100 469.500 ;
        RECT 1251.760 469.240 1252.020 469.500 ;
        RECT 1251.300 379.140 1251.560 379.400 ;
        RECT 1251.300 331.200 1251.560 331.460 ;
        RECT 1251.760 158.820 1252.020 159.080 ;
        RECT 1251.300 158.480 1251.560 158.740 ;
        RECT 1251.300 96.260 1251.560 96.520 ;
        RECT 392.940 59.540 393.200 59.800 ;
        RECT 389.260 16.700 389.520 16.960 ;
        RECT 392.940 16.700 393.200 16.960 ;
      LAYER met2 ;
        RECT 1254.510 1700.410 1254.790 1704.000 ;
        RECT 1254.120 1700.270 1254.790 1700.410 ;
        RECT 1254.120 1677.290 1254.260 1700.270 ;
        RECT 1254.510 1700.000 1254.790 1700.270 ;
        RECT 1251.360 1677.150 1254.260 1677.290 ;
        RECT 1251.360 1655.530 1251.500 1677.150 ;
        RECT 1251.360 1655.390 1251.960 1655.530 ;
        RECT 1251.820 1594.330 1251.960 1655.390 ;
        RECT 1251.360 1594.190 1251.960 1594.330 ;
        RECT 1251.360 1587.110 1251.500 1594.190 ;
        RECT 1251.300 1586.790 1251.560 1587.110 ;
        RECT 1251.760 1538.850 1252.020 1539.170 ;
        RECT 1251.820 1463.090 1251.960 1538.850 ;
        RECT 1251.360 1462.950 1251.960 1463.090 ;
        RECT 1251.360 1415.070 1251.500 1462.950 ;
        RECT 1251.300 1414.750 1251.560 1415.070 ;
        RECT 1251.300 1386.870 1251.560 1387.190 ;
        RECT 1251.360 1345.370 1251.500 1386.870 ;
        RECT 1251.300 1345.050 1251.560 1345.370 ;
        RECT 1252.220 1297.110 1252.480 1297.430 ;
        RECT 1252.280 1249.150 1252.420 1297.110 ;
        RECT 1251.300 1248.830 1251.560 1249.150 ;
        RECT 1252.220 1248.830 1252.480 1249.150 ;
        RECT 1251.360 1207.670 1251.500 1248.830 ;
        RECT 1251.300 1207.350 1251.560 1207.670 ;
        RECT 1251.760 1207.010 1252.020 1207.330 ;
        RECT 1251.820 1176.810 1251.960 1207.010 ;
        RECT 1251.820 1176.670 1252.420 1176.810 ;
        RECT 1252.280 1152.590 1252.420 1176.670 ;
        RECT 1251.300 1152.270 1251.560 1152.590 ;
        RECT 1252.220 1152.270 1252.480 1152.590 ;
        RECT 1251.360 1141.030 1251.500 1152.270 ;
        RECT 1251.300 1140.710 1251.560 1141.030 ;
        RECT 1252.220 1103.990 1252.480 1104.310 ;
        RECT 1252.280 1097.170 1252.420 1103.990 ;
        RECT 1252.220 1096.850 1252.480 1097.170 ;
        RECT 1253.140 1096.850 1253.400 1097.170 ;
        RECT 1253.200 1049.085 1253.340 1096.850 ;
        RECT 1251.750 1048.715 1252.030 1049.085 ;
        RECT 1253.130 1048.715 1253.410 1049.085 ;
        RECT 1251.820 1014.890 1251.960 1048.715 ;
        RECT 1251.760 1014.570 1252.020 1014.890 ;
        RECT 1251.300 1014.230 1251.560 1014.550 ;
        RECT 1251.360 980.210 1251.500 1014.230 ;
        RECT 1251.300 979.890 1251.560 980.210 ;
        RECT 1251.300 979.210 1251.560 979.530 ;
        RECT 1251.360 931.930 1251.500 979.210 ;
        RECT 1251.300 931.610 1251.560 931.930 ;
        RECT 1251.760 930.930 1252.020 931.250 ;
        RECT 1251.820 893.930 1251.960 930.930 ;
        RECT 1251.820 893.790 1252.420 893.930 ;
        RECT 1252.280 869.710 1252.420 893.790 ;
        RECT 1251.300 869.565 1251.560 869.710 ;
        RECT 1252.220 869.565 1252.480 869.710 ;
        RECT 1251.290 869.195 1251.570 869.565 ;
        RECT 1252.210 869.195 1252.490 869.565 ;
        RECT 1252.280 834.090 1252.420 869.195 ;
        RECT 1251.820 833.950 1252.420 834.090 ;
        RECT 1251.820 786.750 1251.960 833.950 ;
        RECT 1251.760 786.430 1252.020 786.750 ;
        RECT 1251.300 786.090 1251.560 786.410 ;
        RECT 1251.360 738.470 1251.500 786.090 ;
        RECT 1251.300 738.150 1251.560 738.470 ;
        RECT 1251.760 737.810 1252.020 738.130 ;
        RECT 1251.820 677.125 1251.960 737.810 ;
        RECT 1251.750 676.755 1252.030 677.125 ;
        RECT 1251.290 676.075 1251.570 676.445 ;
        RECT 1251.300 675.930 1251.560 676.075 ;
        RECT 1252.220 675.930 1252.480 676.250 ;
        RECT 1252.280 650.490 1252.420 675.930 ;
        RECT 1251.820 650.350 1252.420 650.490 ;
        RECT 1251.820 590.230 1251.960 650.350 ;
        RECT 1251.760 589.910 1252.020 590.230 ;
        RECT 1252.220 565.770 1252.480 566.090 ;
        RECT 1252.280 524.610 1252.420 565.770 ;
        RECT 1251.300 524.290 1251.560 524.610 ;
        RECT 1252.220 524.290 1252.480 524.610 ;
        RECT 1251.360 493.410 1251.500 524.290 ;
        RECT 1250.900 493.270 1251.500 493.410 ;
        RECT 1250.900 469.530 1251.040 493.270 ;
        RECT 1250.840 469.210 1251.100 469.530 ;
        RECT 1251.760 469.210 1252.020 469.530 ;
        RECT 1251.820 434.930 1251.960 469.210 ;
        RECT 1251.360 434.790 1251.960 434.930 ;
        RECT 1251.360 379.430 1251.500 434.790 ;
        RECT 1251.300 379.110 1251.560 379.430 ;
        RECT 1251.300 331.170 1251.560 331.490 ;
        RECT 1251.360 318.650 1251.500 331.170 ;
        RECT 1251.360 318.510 1251.960 318.650 ;
        RECT 1251.820 289.580 1251.960 318.510 ;
        RECT 1251.820 289.440 1252.420 289.580 ;
        RECT 1252.280 264.930 1252.420 289.440 ;
        RECT 1251.820 264.790 1252.420 264.930 ;
        RECT 1251.820 159.110 1251.960 264.790 ;
        RECT 1251.760 158.790 1252.020 159.110 ;
        RECT 1251.300 158.450 1251.560 158.770 ;
        RECT 1251.360 96.550 1251.500 158.450 ;
        RECT 1251.300 96.230 1251.560 96.550 ;
        RECT 392.940 59.510 393.200 59.830 ;
        RECT 393.000 16.990 393.140 59.510 ;
        RECT 389.260 16.670 389.520 16.990 ;
        RECT 392.940 16.670 393.200 16.990 ;
        RECT 389.320 2.400 389.460 16.670 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 1251.750 1048.760 1252.030 1049.040 ;
        RECT 1253.130 1048.760 1253.410 1049.040 ;
        RECT 1251.290 869.240 1251.570 869.520 ;
        RECT 1252.210 869.240 1252.490 869.520 ;
        RECT 1251.750 676.800 1252.030 677.080 ;
        RECT 1251.290 676.120 1251.570 676.400 ;
      LAYER met3 ;
        RECT 1251.725 1049.050 1252.055 1049.065 ;
        RECT 1253.105 1049.050 1253.435 1049.065 ;
        RECT 1251.725 1048.750 1253.435 1049.050 ;
        RECT 1251.725 1048.735 1252.055 1048.750 ;
        RECT 1253.105 1048.735 1253.435 1048.750 ;
        RECT 1251.265 869.530 1251.595 869.545 ;
        RECT 1252.185 869.530 1252.515 869.545 ;
        RECT 1251.265 869.230 1252.515 869.530 ;
        RECT 1251.265 869.215 1251.595 869.230 ;
        RECT 1252.185 869.215 1252.515 869.230 ;
        RECT 1251.725 677.090 1252.055 677.105 ;
        RECT 1251.510 676.775 1252.055 677.090 ;
        RECT 1251.510 676.425 1251.810 676.775 ;
        RECT 1251.265 676.110 1251.810 676.425 ;
        RECT 1251.265 676.095 1251.595 676.110 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1256.790 1679.500 1257.110 1679.560 ;
        RECT 1258.170 1679.500 1258.490 1679.560 ;
        RECT 1256.790 1679.360 1258.490 1679.500 ;
        RECT 1256.790 1679.300 1257.110 1679.360 ;
        RECT 1258.170 1679.300 1258.490 1679.360 ;
        RECT 413.610 60.080 413.930 60.140 ;
        RECT 1256.790 60.080 1257.110 60.140 ;
        RECT 413.610 59.940 1257.110 60.080 ;
        RECT 413.610 59.880 413.930 59.940 ;
        RECT 1256.790 59.880 1257.110 59.940 ;
        RECT 407.170 16.900 407.490 16.960 ;
        RECT 413.610 16.900 413.930 16.960 ;
        RECT 407.170 16.760 413.930 16.900 ;
        RECT 407.170 16.700 407.490 16.760 ;
        RECT 413.610 16.700 413.930 16.760 ;
      LAYER via ;
        RECT 1256.820 1679.300 1257.080 1679.560 ;
        RECT 1258.200 1679.300 1258.460 1679.560 ;
        RECT 413.640 59.880 413.900 60.140 ;
        RECT 1256.820 59.880 1257.080 60.140 ;
        RECT 407.200 16.700 407.460 16.960 ;
        RECT 413.640 16.700 413.900 16.960 ;
      LAYER met2 ;
        RECT 1259.570 1700.410 1259.850 1704.000 ;
        RECT 1258.260 1700.270 1259.850 1700.410 ;
        RECT 1258.260 1679.590 1258.400 1700.270 ;
        RECT 1259.570 1700.000 1259.850 1700.270 ;
        RECT 1256.820 1679.270 1257.080 1679.590 ;
        RECT 1258.200 1679.270 1258.460 1679.590 ;
        RECT 1256.880 60.170 1257.020 1679.270 ;
        RECT 413.640 59.850 413.900 60.170 ;
        RECT 1256.820 59.850 1257.080 60.170 ;
        RECT 413.700 16.990 413.840 59.850 ;
        RECT 407.200 16.670 407.460 16.990 ;
        RECT 413.640 16.670 413.900 16.990 ;
        RECT 407.260 2.400 407.400 16.670 ;
        RECT 407.050 -4.800 407.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 0.300 ;
=======
      LAYER met1 ;
        RECT 68.610 58.720 68.930 58.780 ;
        RECT 1167.550 58.720 1167.870 58.780 ;
        RECT 68.610 58.580 1167.870 58.720 ;
        RECT 68.610 58.520 68.930 58.580 ;
        RECT 1167.550 58.520 1167.870 58.580 ;
      LAYER via ;
        RECT 68.640 58.520 68.900 58.780 ;
        RECT 1167.580 58.520 1167.840 58.780 ;
      LAYER met2 ;
        RECT 1168.030 1700.410 1168.310 1704.000 ;
        RECT 1167.640 1700.270 1168.310 1700.410 ;
        RECT 1167.640 58.810 1167.780 1700.270 ;
        RECT 1168.030 1700.000 1168.310 1700.270 ;
        RECT 68.640 58.490 68.900 58.810 ;
        RECT 1167.580 58.490 1167.840 58.810 ;
        RECT 68.700 3.130 68.840 58.490 ;
        RECT 68.240 2.990 68.840 3.130 ;
        RECT 68.240 2.400 68.380 2.990 ;
        RECT 68.030 -4.800 68.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 0.300 ;
=======
      LAYER met1 ;
        RECT 427.410 60.420 427.730 60.480 ;
        RECT 1264.150 60.420 1264.470 60.480 ;
        RECT 427.410 60.280 1264.470 60.420 ;
        RECT 427.410 60.220 427.730 60.280 ;
        RECT 1264.150 60.220 1264.470 60.280 ;
        RECT 424.650 16.560 424.970 16.620 ;
        RECT 427.410 16.560 427.730 16.620 ;
        RECT 424.650 16.420 427.730 16.560 ;
        RECT 424.650 16.360 424.970 16.420 ;
        RECT 427.410 16.360 427.730 16.420 ;
      LAYER via ;
        RECT 427.440 60.220 427.700 60.480 ;
        RECT 1264.180 60.220 1264.440 60.480 ;
        RECT 424.680 16.360 424.940 16.620 ;
        RECT 427.440 16.360 427.700 16.620 ;
      LAYER met2 ;
        RECT 1264.170 1700.000 1264.450 1704.000 ;
        RECT 1264.240 60.510 1264.380 1700.000 ;
        RECT 427.440 60.190 427.700 60.510 ;
        RECT 1264.180 60.190 1264.440 60.510 ;
        RECT 427.500 16.650 427.640 60.190 ;
        RECT 424.680 16.330 424.940 16.650 ;
        RECT 427.440 16.330 427.700 16.650 ;
        RECT 424.740 2.400 424.880 16.330 ;
        RECT 424.530 -4.800 425.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1263.690 1678.140 1264.010 1678.200 ;
        RECT 1267.830 1678.140 1268.150 1678.200 ;
        RECT 1263.690 1678.000 1268.150 1678.140 ;
        RECT 1263.690 1677.940 1264.010 1678.000 ;
        RECT 1267.830 1677.940 1268.150 1678.000 ;
        RECT 448.110 60.760 448.430 60.820 ;
        RECT 1263.690 60.760 1264.010 60.820 ;
        RECT 448.110 60.620 1264.010 60.760 ;
        RECT 448.110 60.560 448.430 60.620 ;
        RECT 1263.690 60.560 1264.010 60.620 ;
        RECT 442.590 16.560 442.910 16.620 ;
        RECT 448.110 16.560 448.430 16.620 ;
        RECT 442.590 16.420 448.430 16.560 ;
        RECT 442.590 16.360 442.910 16.420 ;
        RECT 448.110 16.360 448.430 16.420 ;
      LAYER via ;
        RECT 1263.720 1677.940 1263.980 1678.200 ;
        RECT 1267.860 1677.940 1268.120 1678.200 ;
        RECT 448.140 60.560 448.400 60.820 ;
        RECT 1263.720 60.560 1263.980 60.820 ;
        RECT 442.620 16.360 442.880 16.620 ;
        RECT 448.140 16.360 448.400 16.620 ;
      LAYER met2 ;
        RECT 1269.230 1700.410 1269.510 1704.000 ;
        RECT 1267.920 1700.270 1269.510 1700.410 ;
        RECT 1267.920 1678.230 1268.060 1700.270 ;
        RECT 1269.230 1700.000 1269.510 1700.270 ;
        RECT 1263.720 1677.910 1263.980 1678.230 ;
        RECT 1267.860 1677.910 1268.120 1678.230 ;
        RECT 1263.780 60.850 1263.920 1677.910 ;
        RECT 448.140 60.530 448.400 60.850 ;
        RECT 1263.720 60.530 1263.980 60.850 ;
        RECT 448.200 16.650 448.340 60.530 ;
        RECT 442.620 16.330 442.880 16.650 ;
        RECT 448.140 16.330 448.400 16.650 ;
        RECT 442.680 2.400 442.820 16.330 ;
        RECT 442.470 -4.800 443.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 0.300 ;
=======
      LAYER li1 ;
        RECT 1272.045 1449.165 1272.215 1497.275 ;
        RECT 1271.585 710.685 1271.755 738.395 ;
        RECT 1271.585 469.285 1271.755 502.095 ;
        RECT 1271.585 179.605 1271.755 227.715 ;
        RECT 1272.045 60.945 1272.215 131.155 ;
      LAYER mcon ;
        RECT 1272.045 1497.105 1272.215 1497.275 ;
        RECT 1271.585 738.225 1271.755 738.395 ;
        RECT 1271.585 501.925 1271.755 502.095 ;
        RECT 1271.585 227.545 1271.755 227.715 ;
        RECT 1272.045 130.985 1272.215 131.155 ;
      LAYER met1 ;
        RECT 1271.510 1545.880 1271.830 1545.940 ;
        RECT 1271.970 1545.880 1272.290 1545.940 ;
        RECT 1271.510 1545.740 1272.290 1545.880 ;
        RECT 1271.510 1545.680 1271.830 1545.740 ;
        RECT 1271.970 1545.680 1272.290 1545.740 ;
        RECT 1271.510 1511.340 1271.830 1511.600 ;
        RECT 1271.600 1510.520 1271.740 1511.340 ;
        RECT 1271.970 1510.520 1272.290 1510.580 ;
        RECT 1271.600 1510.380 1272.290 1510.520 ;
        RECT 1271.970 1510.320 1272.290 1510.380 ;
        RECT 1271.970 1497.260 1272.290 1497.320 ;
        RECT 1271.775 1497.120 1272.290 1497.260 ;
        RECT 1271.970 1497.060 1272.290 1497.120 ;
        RECT 1271.970 1449.320 1272.290 1449.380 ;
        RECT 1271.775 1449.180 1272.290 1449.320 ;
        RECT 1271.970 1449.120 1272.290 1449.180 ;
        RECT 1271.510 1269.600 1271.830 1269.860 ;
        RECT 1271.600 1269.120 1271.740 1269.600 ;
        RECT 1271.970 1269.120 1272.290 1269.180 ;
        RECT 1271.600 1268.980 1272.290 1269.120 ;
        RECT 1271.970 1268.920 1272.290 1268.980 ;
        RECT 1271.970 1207.920 1272.290 1207.980 ;
        RECT 1271.600 1207.780 1272.290 1207.920 ;
        RECT 1271.600 1207.640 1271.740 1207.780 ;
        RECT 1271.970 1207.720 1272.290 1207.780 ;
        RECT 1271.510 1207.380 1271.830 1207.640 ;
        RECT 1271.510 1152.500 1271.830 1152.560 ;
        RECT 1271.970 1152.500 1272.290 1152.560 ;
        RECT 1271.510 1152.360 1272.290 1152.500 ;
        RECT 1271.510 1152.300 1271.830 1152.360 ;
        RECT 1271.970 1152.300 1272.290 1152.360 ;
        RECT 1271.510 966.180 1271.830 966.240 ;
        RECT 1271.970 966.180 1272.290 966.240 ;
        RECT 1271.510 966.040 1272.290 966.180 ;
        RECT 1271.510 965.980 1271.830 966.040 ;
        RECT 1271.970 965.980 1272.290 966.040 ;
        RECT 1270.590 959.040 1270.910 959.100 ;
        RECT 1271.970 959.040 1272.290 959.100 ;
        RECT 1270.590 958.900 1272.290 959.040 ;
        RECT 1270.590 958.840 1270.910 958.900 ;
        RECT 1271.970 958.840 1272.290 958.900 ;
        RECT 1271.510 910.760 1271.830 910.820 ;
        RECT 1272.430 910.760 1272.750 910.820 ;
        RECT 1271.510 910.620 1272.750 910.760 ;
        RECT 1271.510 910.560 1271.830 910.620 ;
        RECT 1272.430 910.560 1272.750 910.620 ;
        RECT 1271.510 759.260 1271.830 759.520 ;
        RECT 1271.600 758.840 1271.740 759.260 ;
        RECT 1271.510 758.580 1271.830 758.840 ;
        RECT 1271.510 738.380 1271.830 738.440 ;
        RECT 1271.315 738.240 1271.830 738.380 ;
        RECT 1271.510 738.180 1271.830 738.240 ;
        RECT 1271.525 710.840 1271.815 710.885 ;
        RECT 1272.430 710.840 1272.750 710.900 ;
        RECT 1271.525 710.700 1272.750 710.840 ;
        RECT 1271.525 710.655 1271.815 710.700 ;
        RECT 1272.430 710.640 1272.750 710.700 ;
        RECT 1271.510 572.940 1271.830 573.200 ;
        RECT 1271.600 572.800 1271.740 572.940 ;
        RECT 1271.970 572.800 1272.290 572.860 ;
        RECT 1271.600 572.660 1272.290 572.800 ;
        RECT 1271.970 572.600 1272.290 572.660 ;
        RECT 1271.510 502.080 1271.830 502.140 ;
        RECT 1271.315 501.940 1271.830 502.080 ;
        RECT 1271.510 501.880 1271.830 501.940 ;
        RECT 1271.525 469.440 1271.815 469.485 ;
        RECT 1271.970 469.440 1272.290 469.500 ;
        RECT 1271.525 469.300 1272.290 469.440 ;
        RECT 1271.525 469.255 1271.815 469.300 ;
        RECT 1271.970 469.240 1272.290 469.300 ;
        RECT 1271.510 283.120 1271.830 283.180 ;
        RECT 1272.430 283.120 1272.750 283.180 ;
        RECT 1271.510 282.980 1272.750 283.120 ;
        RECT 1271.510 282.920 1271.830 282.980 ;
        RECT 1272.430 282.920 1272.750 282.980 ;
        RECT 1271.510 227.700 1271.830 227.760 ;
        RECT 1271.315 227.560 1271.830 227.700 ;
        RECT 1271.510 227.500 1271.830 227.560 ;
        RECT 1271.525 179.760 1271.815 179.805 ;
        RECT 1272.430 179.760 1272.750 179.820 ;
        RECT 1271.525 179.620 1272.750 179.760 ;
        RECT 1271.525 179.575 1271.815 179.620 ;
        RECT 1272.430 179.560 1272.750 179.620 ;
        RECT 1271.970 131.140 1272.290 131.200 ;
        RECT 1271.775 131.000 1272.290 131.140 ;
        RECT 1271.970 130.940 1272.290 131.000 ;
        RECT 461.910 61.100 462.230 61.160 ;
        RECT 1271.985 61.100 1272.275 61.145 ;
        RECT 461.910 60.960 1272.275 61.100 ;
        RECT 461.910 60.900 462.230 60.960 ;
        RECT 1271.985 60.915 1272.275 60.960 ;
        RECT 460.530 2.960 460.850 3.020 ;
        RECT 461.910 2.960 462.230 3.020 ;
        RECT 460.530 2.820 462.230 2.960 ;
        RECT 460.530 2.760 460.850 2.820 ;
        RECT 461.910 2.760 462.230 2.820 ;
      LAYER via ;
        RECT 1271.540 1545.680 1271.800 1545.940 ;
        RECT 1272.000 1545.680 1272.260 1545.940 ;
        RECT 1271.540 1511.340 1271.800 1511.600 ;
        RECT 1272.000 1510.320 1272.260 1510.580 ;
        RECT 1272.000 1497.060 1272.260 1497.320 ;
        RECT 1272.000 1449.120 1272.260 1449.380 ;
        RECT 1271.540 1269.600 1271.800 1269.860 ;
        RECT 1272.000 1268.920 1272.260 1269.180 ;
        RECT 1272.000 1207.720 1272.260 1207.980 ;
        RECT 1271.540 1207.380 1271.800 1207.640 ;
        RECT 1271.540 1152.300 1271.800 1152.560 ;
        RECT 1272.000 1152.300 1272.260 1152.560 ;
        RECT 1271.540 965.980 1271.800 966.240 ;
        RECT 1272.000 965.980 1272.260 966.240 ;
        RECT 1270.620 958.840 1270.880 959.100 ;
        RECT 1272.000 958.840 1272.260 959.100 ;
        RECT 1271.540 910.560 1271.800 910.820 ;
        RECT 1272.460 910.560 1272.720 910.820 ;
        RECT 1271.540 759.260 1271.800 759.520 ;
        RECT 1271.540 758.580 1271.800 758.840 ;
        RECT 1271.540 738.180 1271.800 738.440 ;
        RECT 1272.460 710.640 1272.720 710.900 ;
        RECT 1271.540 572.940 1271.800 573.200 ;
        RECT 1272.000 572.600 1272.260 572.860 ;
        RECT 1271.540 501.880 1271.800 502.140 ;
        RECT 1272.000 469.240 1272.260 469.500 ;
        RECT 1271.540 282.920 1271.800 283.180 ;
        RECT 1272.460 282.920 1272.720 283.180 ;
        RECT 1271.540 227.500 1271.800 227.760 ;
        RECT 1272.460 179.560 1272.720 179.820 ;
        RECT 1272.000 130.940 1272.260 131.200 ;
        RECT 461.940 60.900 462.200 61.160 ;
        RECT 460.560 2.760 460.820 3.020 ;
        RECT 461.940 2.760 462.200 3.020 ;
      LAYER met2 ;
        RECT 1273.830 1700.000 1274.110 1704.000 ;
        RECT 1273.900 1678.140 1274.040 1700.000 ;
        RECT 1272.060 1678.000 1274.040 1678.140 ;
        RECT 1272.060 1605.210 1272.200 1678.000 ;
        RECT 1271.600 1605.070 1272.200 1605.210 ;
        RECT 1271.600 1603.850 1271.740 1605.070 ;
        RECT 1271.600 1603.710 1272.200 1603.850 ;
        RECT 1272.060 1545.970 1272.200 1603.710 ;
        RECT 1271.540 1545.650 1271.800 1545.970 ;
        RECT 1272.000 1545.650 1272.260 1545.970 ;
        RECT 1271.600 1511.630 1271.740 1545.650 ;
        RECT 1271.540 1511.310 1271.800 1511.630 ;
        RECT 1272.000 1510.290 1272.260 1510.610 ;
        RECT 1272.060 1497.350 1272.200 1510.290 ;
        RECT 1272.000 1497.030 1272.260 1497.350 ;
        RECT 1272.000 1449.090 1272.260 1449.410 ;
        RECT 1272.060 1402.005 1272.200 1449.090 ;
        RECT 1271.990 1401.635 1272.270 1402.005 ;
        RECT 1271.530 1400.955 1271.810 1401.325 ;
        RECT 1271.600 1269.890 1271.740 1400.955 ;
        RECT 1271.540 1269.570 1271.800 1269.890 ;
        RECT 1272.000 1268.890 1272.260 1269.210 ;
        RECT 1272.060 1208.010 1272.200 1268.890 ;
        RECT 1272.000 1207.690 1272.260 1208.010 ;
        RECT 1271.540 1207.350 1271.800 1207.670 ;
        RECT 1271.600 1152.590 1271.740 1207.350 ;
        RECT 1271.540 1152.270 1271.800 1152.590 ;
        RECT 1272.000 1152.270 1272.260 1152.590 ;
        RECT 1272.060 1112.210 1272.200 1152.270 ;
        RECT 1271.600 1112.070 1272.200 1112.210 ;
        RECT 1271.600 1110.850 1271.740 1112.070 ;
        RECT 1271.600 1110.710 1272.200 1110.850 ;
        RECT 1272.060 979.610 1272.200 1110.710 ;
        RECT 1271.600 979.470 1272.200 979.610 ;
        RECT 1271.600 966.270 1271.740 979.470 ;
        RECT 1271.540 965.950 1271.800 966.270 ;
        RECT 1272.000 965.950 1272.260 966.270 ;
        RECT 1272.060 959.130 1272.200 965.950 ;
        RECT 1270.620 958.810 1270.880 959.130 ;
        RECT 1272.000 958.810 1272.260 959.130 ;
        RECT 1270.680 911.045 1270.820 958.810 ;
        RECT 1270.610 910.675 1270.890 911.045 ;
        RECT 1271.530 910.675 1271.810 911.045 ;
        RECT 1271.540 910.530 1271.800 910.675 ;
        RECT 1272.460 910.530 1272.720 910.850 ;
        RECT 1272.520 821.285 1272.660 910.530 ;
        RECT 1271.530 820.915 1271.810 821.285 ;
        RECT 1272.450 820.915 1272.730 821.285 ;
        RECT 1271.600 759.550 1271.740 820.915 ;
        RECT 1271.540 759.230 1271.800 759.550 ;
        RECT 1271.540 758.550 1271.800 758.870 ;
        RECT 1271.600 738.470 1271.740 758.550 ;
        RECT 1271.540 738.150 1271.800 738.470 ;
        RECT 1272.460 710.610 1272.720 710.930 ;
        RECT 1272.520 689.250 1272.660 710.610 ;
        RECT 1272.060 689.110 1272.660 689.250 ;
        RECT 1272.060 628.845 1272.200 689.110 ;
        RECT 1271.990 628.475 1272.270 628.845 ;
        RECT 1271.530 627.795 1271.810 628.165 ;
        RECT 1271.600 573.230 1271.740 627.795 ;
        RECT 1271.540 572.910 1271.800 573.230 ;
        RECT 1272.000 572.570 1272.260 572.890 ;
        RECT 1272.060 548.490 1272.200 572.570 ;
        RECT 1271.600 548.350 1272.200 548.490 ;
        RECT 1271.600 502.170 1271.740 548.350 ;
        RECT 1271.540 501.850 1271.800 502.170 ;
        RECT 1272.000 469.210 1272.260 469.530 ;
        RECT 1272.060 414.530 1272.200 469.210 ;
        RECT 1272.060 414.390 1272.660 414.530 ;
        RECT 1272.520 283.210 1272.660 414.390 ;
        RECT 1271.540 282.890 1271.800 283.210 ;
        RECT 1272.460 282.890 1272.720 283.210 ;
        RECT 1271.600 227.790 1271.740 282.890 ;
        RECT 1271.540 227.470 1271.800 227.790 ;
        RECT 1272.460 179.530 1272.720 179.850 ;
        RECT 1272.520 131.650 1272.660 179.530 ;
        RECT 1272.060 131.510 1272.660 131.650 ;
        RECT 1272.060 131.230 1272.200 131.510 ;
        RECT 1272.000 130.910 1272.260 131.230 ;
        RECT 461.940 60.870 462.200 61.190 ;
        RECT 462.000 3.050 462.140 60.870 ;
        RECT 460.560 2.730 460.820 3.050 ;
        RECT 461.940 2.730 462.200 3.050 ;
        RECT 460.620 2.400 460.760 2.730 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 1271.990 1401.680 1272.270 1401.960 ;
        RECT 1271.530 1401.000 1271.810 1401.280 ;
        RECT 1270.610 910.720 1270.890 911.000 ;
        RECT 1271.530 910.720 1271.810 911.000 ;
        RECT 1271.530 820.960 1271.810 821.240 ;
        RECT 1272.450 820.960 1272.730 821.240 ;
        RECT 1271.990 628.520 1272.270 628.800 ;
        RECT 1271.530 627.840 1271.810 628.120 ;
      LAYER met3 ;
        RECT 1271.965 1401.970 1272.295 1401.985 ;
        RECT 1270.830 1401.670 1272.295 1401.970 ;
        RECT 1270.830 1401.290 1271.130 1401.670 ;
        RECT 1271.965 1401.655 1272.295 1401.670 ;
        RECT 1271.505 1401.290 1271.835 1401.305 ;
        RECT 1270.830 1400.990 1271.835 1401.290 ;
        RECT 1271.505 1400.975 1271.835 1400.990 ;
        RECT 1270.585 911.010 1270.915 911.025 ;
        RECT 1271.505 911.010 1271.835 911.025 ;
        RECT 1270.585 910.710 1271.835 911.010 ;
        RECT 1270.585 910.695 1270.915 910.710 ;
        RECT 1271.505 910.695 1271.835 910.710 ;
        RECT 1271.505 821.250 1271.835 821.265 ;
        RECT 1272.425 821.250 1272.755 821.265 ;
        RECT 1271.505 820.950 1272.755 821.250 ;
        RECT 1271.505 820.935 1271.835 820.950 ;
        RECT 1272.425 820.935 1272.755 820.950 ;
        RECT 1271.965 628.810 1272.295 628.825 ;
        RECT 1271.750 628.495 1272.295 628.810 ;
        RECT 1271.750 628.145 1272.050 628.495 ;
        RECT 1271.505 627.830 1272.050 628.145 ;
        RECT 1271.505 627.815 1271.835 627.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 0.300 ;
=======
      LAYER met1 ;
        RECT 482.610 61.440 482.930 61.500 ;
        RECT 1277.490 61.440 1277.810 61.500 ;
        RECT 482.610 61.300 1277.810 61.440 ;
        RECT 482.610 61.240 482.930 61.300 ;
        RECT 1277.490 61.240 1277.810 61.300 ;
        RECT 478.470 15.880 478.790 15.940 ;
        RECT 482.610 15.880 482.930 15.940 ;
        RECT 478.470 15.740 482.930 15.880 ;
        RECT 478.470 15.680 478.790 15.740 ;
        RECT 482.610 15.680 482.930 15.740 ;
      LAYER via ;
        RECT 482.640 61.240 482.900 61.500 ;
        RECT 1277.520 61.240 1277.780 61.500 ;
        RECT 478.500 15.680 478.760 15.940 ;
        RECT 482.640 15.680 482.900 15.940 ;
      LAYER met2 ;
        RECT 1278.890 1700.410 1279.170 1704.000 ;
        RECT 1277.580 1700.270 1279.170 1700.410 ;
        RECT 1277.580 61.530 1277.720 1700.270 ;
        RECT 1278.890 1700.000 1279.170 1700.270 ;
        RECT 482.640 61.210 482.900 61.530 ;
        RECT 1277.520 61.210 1277.780 61.530 ;
        RECT 482.700 15.970 482.840 61.210 ;
        RECT 478.500 15.650 478.760 15.970 ;
        RECT 482.640 15.650 482.900 15.970 ;
        RECT 478.560 2.400 478.700 15.650 ;
        RECT 478.350 -4.800 478.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 0.300 ;
=======
      LAYER met1 ;
        RECT 496.410 61.780 496.730 61.840 ;
        RECT 1284.850 61.780 1285.170 61.840 ;
        RECT 496.410 61.640 1285.170 61.780 ;
        RECT 496.410 61.580 496.730 61.640 ;
        RECT 1284.850 61.580 1285.170 61.640 ;
      LAYER via ;
        RECT 496.440 61.580 496.700 61.840 ;
        RECT 1284.880 61.580 1285.140 61.840 ;
      LAYER met2 ;
        RECT 1283.490 1700.410 1283.770 1704.000 ;
        RECT 1283.490 1700.270 1285.080 1700.410 ;
        RECT 1283.490 1700.000 1283.770 1700.270 ;
        RECT 1284.940 61.870 1285.080 1700.270 ;
        RECT 496.440 61.550 496.700 61.870 ;
        RECT 1284.880 61.550 1285.140 61.870 ;
        RECT 496.500 2.400 496.640 61.550 ;
        RECT 496.290 -4.800 496.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1284.390 1670.320 1284.710 1670.380 ;
        RECT 1287.150 1670.320 1287.470 1670.380 ;
        RECT 1284.390 1670.180 1287.470 1670.320 ;
        RECT 1284.390 1670.120 1284.710 1670.180 ;
        RECT 1287.150 1670.120 1287.470 1670.180 ;
        RECT 517.110 62.120 517.430 62.180 ;
        RECT 1284.390 62.120 1284.710 62.180 ;
        RECT 517.110 61.980 1284.710 62.120 ;
        RECT 517.110 61.920 517.430 61.980 ;
        RECT 1284.390 61.920 1284.710 61.980 ;
        RECT 513.890 15.880 514.210 15.940 ;
        RECT 517.110 15.880 517.430 15.940 ;
        RECT 513.890 15.740 517.430 15.880 ;
        RECT 513.890 15.680 514.210 15.740 ;
        RECT 517.110 15.680 517.430 15.740 ;
      LAYER via ;
        RECT 1284.420 1670.120 1284.680 1670.380 ;
        RECT 1287.180 1670.120 1287.440 1670.380 ;
        RECT 517.140 61.920 517.400 62.180 ;
        RECT 1284.420 61.920 1284.680 62.180 ;
        RECT 513.920 15.680 514.180 15.940 ;
        RECT 517.140 15.680 517.400 15.940 ;
      LAYER met2 ;
        RECT 1288.550 1700.410 1288.830 1704.000 ;
        RECT 1287.240 1700.270 1288.830 1700.410 ;
        RECT 1287.240 1670.410 1287.380 1700.270 ;
        RECT 1288.550 1700.000 1288.830 1700.270 ;
        RECT 1284.420 1670.090 1284.680 1670.410 ;
        RECT 1287.180 1670.090 1287.440 1670.410 ;
        RECT 1284.480 62.210 1284.620 1670.090 ;
        RECT 517.140 61.890 517.400 62.210 ;
        RECT 1284.420 61.890 1284.680 62.210 ;
        RECT 517.200 15.970 517.340 61.890 ;
        RECT 513.920 15.650 514.180 15.970 ;
        RECT 517.140 15.650 517.400 15.970 ;
        RECT 513.980 2.400 514.120 15.650 ;
        RECT 513.770 -4.800 514.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 0.300 ;
=======
      LAYER met1 ;
        RECT 537.810 58.380 538.130 58.440 ;
        RECT 1292.210 58.380 1292.530 58.440 ;
        RECT 537.810 58.240 1292.530 58.380 ;
        RECT 537.810 58.180 538.130 58.240 ;
        RECT 1292.210 58.180 1292.530 58.240 ;
        RECT 531.830 15.880 532.150 15.940 ;
        RECT 537.810 15.880 538.130 15.940 ;
        RECT 531.830 15.740 538.130 15.880 ;
        RECT 531.830 15.680 532.150 15.740 ;
        RECT 537.810 15.680 538.130 15.740 ;
      LAYER via ;
        RECT 537.840 58.180 538.100 58.440 ;
        RECT 1292.240 58.180 1292.500 58.440 ;
        RECT 531.860 15.680 532.120 15.940 ;
        RECT 537.840 15.680 538.100 15.940 ;
      LAYER met2 ;
        RECT 1293.150 1700.410 1293.430 1704.000 ;
        RECT 1292.300 1700.270 1293.430 1700.410 ;
        RECT 1292.300 58.470 1292.440 1700.270 ;
        RECT 1293.150 1700.000 1293.430 1700.270 ;
        RECT 537.840 58.150 538.100 58.470 ;
        RECT 1292.240 58.150 1292.500 58.470 ;
        RECT 537.900 15.970 538.040 58.150 ;
        RECT 531.860 15.650 532.120 15.970 ;
        RECT 537.840 15.650 538.100 15.970 ;
        RECT 531.920 2.400 532.060 15.650 ;
        RECT 531.710 -4.800 532.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 0.300 ;
=======
      LAYER met1 ;
        RECT 886.490 1684.940 886.810 1685.000 ;
        RECT 1298.190 1684.940 1298.510 1685.000 ;
        RECT 886.490 1684.800 1298.510 1684.940 ;
        RECT 886.490 1684.740 886.810 1684.800 ;
        RECT 1298.190 1684.740 1298.510 1684.800 ;
        RECT 549.770 26.420 550.090 26.480 ;
        RECT 886.490 26.420 886.810 26.480 ;
        RECT 549.770 26.280 886.810 26.420 ;
        RECT 549.770 26.220 550.090 26.280 ;
        RECT 886.490 26.220 886.810 26.280 ;
      LAYER via ;
        RECT 886.520 1684.740 886.780 1685.000 ;
        RECT 1298.220 1684.740 1298.480 1685.000 ;
        RECT 549.800 26.220 550.060 26.480 ;
        RECT 886.520 26.220 886.780 26.480 ;
      LAYER met2 ;
        RECT 1298.210 1700.000 1298.490 1704.000 ;
        RECT 1298.280 1685.030 1298.420 1700.000 ;
        RECT 886.520 1684.710 886.780 1685.030 ;
        RECT 1298.220 1684.710 1298.480 1685.030 ;
        RECT 886.580 26.510 886.720 1684.710 ;
        RECT 549.800 26.190 550.060 26.510 ;
        RECT 886.520 26.190 886.780 26.510 ;
        RECT 549.860 2.400 550.000 26.190 ;
        RECT 549.650 -4.800 550.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 0.300 ;
=======
      LAYER li1 ;
        RECT 1298.265 1338.665 1298.435 1345.975 ;
        RECT 1298.265 655.605 1298.435 703.375 ;
        RECT 1298.265 559.045 1298.435 607.155 ;
        RECT 1298.265 493.425 1298.435 517.395 ;
        RECT 1298.265 372.725 1298.435 380.035 ;
        RECT 1298.265 324.445 1298.435 331.415 ;
        RECT 600.905 15.045 601.075 17.935 ;
      LAYER mcon ;
        RECT 1298.265 1345.805 1298.435 1345.975 ;
        RECT 1298.265 703.205 1298.435 703.375 ;
        RECT 1298.265 606.985 1298.435 607.155 ;
        RECT 1298.265 517.225 1298.435 517.395 ;
        RECT 1298.265 379.865 1298.435 380.035 ;
        RECT 1298.265 331.245 1298.435 331.415 ;
        RECT 600.905 17.765 601.075 17.935 ;
      LAYER met1 ;
        RECT 1298.650 1387.100 1298.970 1387.160 ;
        RECT 1299.570 1387.100 1299.890 1387.160 ;
        RECT 1298.650 1386.960 1299.890 1387.100 ;
        RECT 1298.650 1386.900 1298.970 1386.960 ;
        RECT 1299.570 1386.900 1299.890 1386.960 ;
        RECT 1298.205 1345.960 1298.495 1346.005 ;
        RECT 1298.650 1345.960 1298.970 1346.020 ;
        RECT 1298.205 1345.820 1298.970 1345.960 ;
        RECT 1298.205 1345.775 1298.495 1345.820 ;
        RECT 1298.650 1345.760 1298.970 1345.820 ;
        RECT 1298.190 1338.820 1298.510 1338.880 ;
        RECT 1297.995 1338.680 1298.510 1338.820 ;
        RECT 1298.190 1338.620 1298.510 1338.680 ;
        RECT 1298.190 1152.500 1298.510 1152.560 ;
        RECT 1298.650 1152.500 1298.970 1152.560 ;
        RECT 1298.190 1152.360 1298.970 1152.500 ;
        RECT 1298.190 1152.300 1298.510 1152.360 ;
        RECT 1298.650 1152.300 1298.970 1152.360 ;
        RECT 1298.650 1125.300 1298.970 1125.360 ;
        RECT 1298.280 1125.160 1298.970 1125.300 ;
        RECT 1298.280 1124.680 1298.420 1125.160 ;
        RECT 1298.650 1125.100 1298.970 1125.160 ;
        RECT 1298.190 1124.420 1298.510 1124.680 ;
        RECT 1298.190 959.380 1298.510 959.440 ;
        RECT 1298.650 959.380 1298.970 959.440 ;
        RECT 1298.190 959.240 1298.970 959.380 ;
        RECT 1298.190 959.180 1298.510 959.240 ;
        RECT 1298.650 959.180 1298.970 959.240 ;
        RECT 1297.270 958.700 1297.590 958.760 ;
        RECT 1298.190 958.700 1298.510 958.760 ;
        RECT 1297.270 958.560 1298.510 958.700 ;
        RECT 1297.270 958.500 1297.590 958.560 ;
        RECT 1298.190 958.500 1298.510 958.560 ;
        RECT 1298.650 710.500 1298.970 710.560 ;
        RECT 1299.110 710.500 1299.430 710.560 ;
        RECT 1298.650 710.360 1299.430 710.500 ;
        RECT 1298.650 710.300 1298.970 710.360 ;
        RECT 1299.110 710.300 1299.430 710.360 ;
        RECT 1298.650 703.500 1298.970 703.760 ;
        RECT 1298.205 703.360 1298.495 703.405 ;
        RECT 1298.740 703.360 1298.880 703.500 ;
        RECT 1298.205 703.220 1298.880 703.360 ;
        RECT 1298.205 703.175 1298.495 703.220 ;
        RECT 1298.190 655.760 1298.510 655.820 ;
        RECT 1297.995 655.620 1298.510 655.760 ;
        RECT 1298.190 655.560 1298.510 655.620 ;
        RECT 1297.270 638.420 1297.590 638.480 ;
        RECT 1298.190 638.420 1298.510 638.480 ;
        RECT 1297.270 638.280 1298.510 638.420 ;
        RECT 1297.270 638.220 1297.590 638.280 ;
        RECT 1298.190 638.220 1298.510 638.280 ;
        RECT 1298.190 607.140 1298.510 607.200 ;
        RECT 1297.995 607.000 1298.510 607.140 ;
        RECT 1298.190 606.940 1298.510 607.000 ;
        RECT 1298.205 559.200 1298.495 559.245 ;
        RECT 1299.110 559.200 1299.430 559.260 ;
        RECT 1298.205 559.060 1299.430 559.200 ;
        RECT 1298.205 559.015 1298.495 559.060 ;
        RECT 1299.110 559.000 1299.430 559.060 ;
        RECT 1298.190 542.540 1298.510 542.600 ;
        RECT 1299.110 542.540 1299.430 542.600 ;
        RECT 1298.190 542.400 1299.430 542.540 ;
        RECT 1298.190 542.340 1298.510 542.400 ;
        RECT 1299.110 542.340 1299.430 542.400 ;
        RECT 1298.190 517.380 1298.510 517.440 ;
        RECT 1297.995 517.240 1298.510 517.380 ;
        RECT 1298.190 517.180 1298.510 517.240 ;
        RECT 1298.190 493.580 1298.510 493.640 ;
        RECT 1297.995 493.440 1298.510 493.580 ;
        RECT 1298.190 493.380 1298.510 493.440 ;
        RECT 1298.190 434.760 1298.510 434.820 ;
        RECT 1298.650 434.760 1298.970 434.820 ;
        RECT 1298.190 434.620 1298.970 434.760 ;
        RECT 1298.190 434.560 1298.510 434.620 ;
        RECT 1298.650 434.560 1298.970 434.620 ;
        RECT 1298.205 380.020 1298.495 380.065 ;
        RECT 1298.650 380.020 1298.970 380.080 ;
        RECT 1298.205 379.880 1298.970 380.020 ;
        RECT 1298.205 379.835 1298.495 379.880 ;
        RECT 1298.650 379.820 1298.970 379.880 ;
        RECT 1298.190 372.880 1298.510 372.940 ;
        RECT 1297.995 372.740 1298.510 372.880 ;
        RECT 1298.190 372.680 1298.510 372.740 ;
        RECT 1298.190 331.400 1298.510 331.460 ;
        RECT 1297.995 331.260 1298.510 331.400 ;
        RECT 1298.190 331.200 1298.510 331.260 ;
        RECT 1298.190 324.600 1298.510 324.660 ;
        RECT 1297.995 324.460 1298.510 324.600 ;
        RECT 1298.190 324.400 1298.510 324.460 ;
        RECT 1298.650 145.080 1298.970 145.140 ;
        RECT 1299.110 145.080 1299.430 145.140 ;
        RECT 1298.650 144.940 1299.430 145.080 ;
        RECT 1298.650 144.880 1298.970 144.940 ;
        RECT 1299.110 144.880 1299.430 144.940 ;
        RECT 567.710 17.920 568.030 17.980 ;
        RECT 600.845 17.920 601.135 17.965 ;
        RECT 567.710 17.780 601.135 17.920 ;
        RECT 567.710 17.720 568.030 17.780 ;
        RECT 600.845 17.735 601.135 17.780 ;
        RECT 600.845 15.200 601.135 15.245 ;
        RECT 1298.190 15.200 1298.510 15.260 ;
        RECT 600.845 15.060 1298.510 15.200 ;
        RECT 600.845 15.015 601.135 15.060 ;
        RECT 1298.190 15.000 1298.510 15.060 ;
      LAYER via ;
        RECT 1298.680 1386.900 1298.940 1387.160 ;
        RECT 1299.600 1386.900 1299.860 1387.160 ;
        RECT 1298.680 1345.760 1298.940 1346.020 ;
        RECT 1298.220 1338.620 1298.480 1338.880 ;
        RECT 1298.220 1152.300 1298.480 1152.560 ;
        RECT 1298.680 1152.300 1298.940 1152.560 ;
        RECT 1298.680 1125.100 1298.940 1125.360 ;
        RECT 1298.220 1124.420 1298.480 1124.680 ;
        RECT 1298.220 959.180 1298.480 959.440 ;
        RECT 1298.680 959.180 1298.940 959.440 ;
        RECT 1297.300 958.500 1297.560 958.760 ;
        RECT 1298.220 958.500 1298.480 958.760 ;
        RECT 1298.680 710.300 1298.940 710.560 ;
        RECT 1299.140 710.300 1299.400 710.560 ;
        RECT 1298.680 703.500 1298.940 703.760 ;
        RECT 1298.220 655.560 1298.480 655.820 ;
        RECT 1297.300 638.220 1297.560 638.480 ;
        RECT 1298.220 638.220 1298.480 638.480 ;
        RECT 1298.220 606.940 1298.480 607.200 ;
        RECT 1299.140 559.000 1299.400 559.260 ;
        RECT 1298.220 542.340 1298.480 542.600 ;
        RECT 1299.140 542.340 1299.400 542.600 ;
        RECT 1298.220 517.180 1298.480 517.440 ;
        RECT 1298.220 493.380 1298.480 493.640 ;
        RECT 1298.220 434.560 1298.480 434.820 ;
        RECT 1298.680 434.560 1298.940 434.820 ;
        RECT 1298.680 379.820 1298.940 380.080 ;
        RECT 1298.220 372.680 1298.480 372.940 ;
        RECT 1298.220 331.200 1298.480 331.460 ;
        RECT 1298.220 324.400 1298.480 324.660 ;
        RECT 1298.680 144.880 1298.940 145.140 ;
        RECT 1299.140 144.880 1299.400 145.140 ;
        RECT 567.740 17.720 568.000 17.980 ;
        RECT 1298.220 15.000 1298.480 15.260 ;
      LAYER met2 ;
        RECT 1302.810 1700.410 1303.090 1704.000 ;
        RECT 1302.420 1700.270 1303.090 1700.410 ;
        RECT 1302.420 1656.210 1302.560 1700.270 ;
        RECT 1302.810 1700.000 1303.090 1700.270 ;
        RECT 1298.740 1656.070 1302.560 1656.210 ;
        RECT 1298.740 1435.325 1298.880 1656.070 ;
        RECT 1298.670 1434.955 1298.950 1435.325 ;
        RECT 1299.590 1434.955 1299.870 1435.325 ;
        RECT 1299.660 1387.190 1299.800 1434.955 ;
        RECT 1298.680 1386.870 1298.940 1387.190 ;
        RECT 1299.600 1386.870 1299.860 1387.190 ;
        RECT 1298.740 1346.050 1298.880 1386.870 ;
        RECT 1298.680 1345.730 1298.940 1346.050 ;
        RECT 1298.220 1338.590 1298.480 1338.910 ;
        RECT 1298.280 1152.590 1298.420 1338.590 ;
        RECT 1298.220 1152.270 1298.480 1152.590 ;
        RECT 1298.680 1152.270 1298.940 1152.590 ;
        RECT 1298.740 1125.390 1298.880 1152.270 ;
        RECT 1298.680 1125.070 1298.940 1125.390 ;
        RECT 1298.220 1124.390 1298.480 1124.710 ;
        RECT 1298.280 1007.490 1298.420 1124.390 ;
        RECT 1298.280 1007.350 1298.880 1007.490 ;
        RECT 1298.740 959.470 1298.880 1007.350 ;
        RECT 1298.220 959.150 1298.480 959.470 ;
        RECT 1298.680 959.150 1298.940 959.470 ;
        RECT 1298.280 958.790 1298.420 959.150 ;
        RECT 1297.300 958.470 1297.560 958.790 ;
        RECT 1298.220 958.470 1298.480 958.790 ;
        RECT 1297.360 911.045 1297.500 958.470 ;
        RECT 1297.290 910.675 1297.570 911.045 ;
        RECT 1298.670 910.675 1298.950 911.045 ;
        RECT 1298.740 886.450 1298.880 910.675 ;
        RECT 1298.740 886.310 1299.340 886.450 ;
        RECT 1299.200 821.285 1299.340 886.310 ;
        RECT 1298.210 820.915 1298.490 821.285 ;
        RECT 1299.130 820.915 1299.410 821.285 ;
        RECT 1298.280 766.090 1298.420 820.915 ;
        RECT 1298.280 765.950 1298.880 766.090 ;
        RECT 1298.740 741.610 1298.880 765.950 ;
        RECT 1298.740 741.470 1299.340 741.610 ;
        RECT 1299.200 710.590 1299.340 741.470 ;
        RECT 1298.680 710.270 1298.940 710.590 ;
        RECT 1299.140 710.270 1299.400 710.590 ;
        RECT 1298.740 703.790 1298.880 710.270 ;
        RECT 1298.680 703.470 1298.940 703.790 ;
        RECT 1298.220 655.530 1298.480 655.850 ;
        RECT 1298.280 638.510 1298.420 655.530 ;
        RECT 1297.300 638.190 1297.560 638.510 ;
        RECT 1298.220 638.190 1298.480 638.510 ;
        RECT 1297.360 614.565 1297.500 638.190 ;
        RECT 1297.290 614.195 1297.570 614.565 ;
        RECT 1298.210 614.195 1298.490 614.565 ;
        RECT 1298.280 607.230 1298.420 614.195 ;
        RECT 1298.220 606.910 1298.480 607.230 ;
        RECT 1299.140 558.970 1299.400 559.290 ;
        RECT 1299.200 542.630 1299.340 558.970 ;
        RECT 1298.220 542.310 1298.480 542.630 ;
        RECT 1299.140 542.310 1299.400 542.630 ;
        RECT 1298.280 517.470 1298.420 542.310 ;
        RECT 1298.220 517.150 1298.480 517.470 ;
        RECT 1298.220 493.350 1298.480 493.670 ;
        RECT 1298.280 434.850 1298.420 493.350 ;
        RECT 1298.220 434.530 1298.480 434.850 ;
        RECT 1298.680 434.530 1298.940 434.850 ;
        RECT 1298.740 380.110 1298.880 434.530 ;
        RECT 1298.680 379.790 1298.940 380.110 ;
        RECT 1298.220 372.650 1298.480 372.970 ;
        RECT 1298.280 331.490 1298.420 372.650 ;
        RECT 1298.220 331.170 1298.480 331.490 ;
        RECT 1298.220 324.370 1298.480 324.690 ;
        RECT 1298.280 269.010 1298.420 324.370 ;
        RECT 1298.280 268.870 1298.880 269.010 ;
        RECT 1298.740 210.530 1298.880 268.870 ;
        RECT 1298.740 210.390 1299.800 210.530 ;
        RECT 1299.660 192.850 1299.800 210.390 ;
        RECT 1299.200 192.710 1299.800 192.850 ;
        RECT 1299.200 145.170 1299.340 192.710 ;
        RECT 1298.680 144.850 1298.940 145.170 ;
        RECT 1299.140 144.850 1299.400 145.170 ;
        RECT 1298.740 62.290 1298.880 144.850 ;
        RECT 1298.280 62.150 1298.880 62.290 ;
        RECT 567.740 17.690 568.000 18.010 ;
        RECT 567.800 2.400 567.940 17.690 ;
        RECT 1298.280 15.290 1298.420 62.150 ;
        RECT 1298.220 14.970 1298.480 15.290 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 1298.670 1435.000 1298.950 1435.280 ;
        RECT 1299.590 1435.000 1299.870 1435.280 ;
        RECT 1297.290 910.720 1297.570 911.000 ;
        RECT 1298.670 910.720 1298.950 911.000 ;
        RECT 1298.210 820.960 1298.490 821.240 ;
        RECT 1299.130 820.960 1299.410 821.240 ;
        RECT 1297.290 614.240 1297.570 614.520 ;
        RECT 1298.210 614.240 1298.490 614.520 ;
      LAYER met3 ;
        RECT 1298.645 1435.290 1298.975 1435.305 ;
        RECT 1299.565 1435.290 1299.895 1435.305 ;
        RECT 1298.645 1434.990 1299.895 1435.290 ;
        RECT 1298.645 1434.975 1298.975 1434.990 ;
        RECT 1299.565 1434.975 1299.895 1434.990 ;
        RECT 1297.265 911.010 1297.595 911.025 ;
        RECT 1298.645 911.010 1298.975 911.025 ;
        RECT 1297.265 910.710 1298.975 911.010 ;
        RECT 1297.265 910.695 1297.595 910.710 ;
        RECT 1298.645 910.695 1298.975 910.710 ;
        RECT 1298.185 821.250 1298.515 821.265 ;
        RECT 1299.105 821.250 1299.435 821.265 ;
        RECT 1298.185 820.950 1299.435 821.250 ;
        RECT 1298.185 820.935 1298.515 820.950 ;
        RECT 1299.105 820.935 1299.435 820.950 ;
        RECT 1297.265 614.530 1297.595 614.545 ;
        RECT 1298.185 614.530 1298.515 614.545 ;
        RECT 1297.265 614.230 1298.515 614.530 ;
        RECT 1297.265 614.215 1297.595 614.230 ;
        RECT 1298.185 614.215 1298.515 614.230 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 0.300 ;
=======
      LAYER met1 ;
        RECT 927.890 1684.600 928.210 1684.660 ;
        RECT 1307.850 1684.600 1308.170 1684.660 ;
        RECT 927.890 1684.460 1308.170 1684.600 ;
        RECT 927.890 1684.400 928.210 1684.460 ;
        RECT 1307.850 1684.400 1308.170 1684.460 ;
        RECT 586.110 27.100 586.430 27.160 ;
        RECT 927.890 27.100 928.210 27.160 ;
        RECT 586.110 26.960 928.210 27.100 ;
        RECT 586.110 26.900 586.430 26.960 ;
        RECT 927.890 26.900 928.210 26.960 ;
      LAYER via ;
        RECT 927.920 1684.400 928.180 1684.660 ;
        RECT 1307.880 1684.400 1308.140 1684.660 ;
        RECT 586.140 26.900 586.400 27.160 ;
        RECT 927.920 26.900 928.180 27.160 ;
      LAYER met2 ;
        RECT 1307.870 1700.000 1308.150 1704.000 ;
        RECT 1307.940 1684.690 1308.080 1700.000 ;
        RECT 927.920 1684.370 928.180 1684.690 ;
        RECT 1307.880 1684.370 1308.140 1684.690 ;
        RECT 927.980 27.190 928.120 1684.370 ;
        RECT 586.140 26.870 586.400 27.190 ;
        RECT 927.920 26.870 928.180 27.190 ;
        RECT 586.200 14.010 586.340 26.870 ;
        RECT 585.740 13.870 586.340 14.010 ;
        RECT 585.740 2.400 585.880 13.870 ;
        RECT 585.530 -4.800 586.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 91.490 -4.800 92.050 0.300 ;
=======
        RECT 1174.470 1700.410 1174.750 1704.000 ;
        RECT 1173.160 1700.270 1174.750 1700.410 ;
        RECT 1173.160 19.565 1173.300 1700.270 ;
        RECT 1174.470 1700.000 1174.750 1700.270 ;
        RECT 91.630 19.195 91.910 19.565 ;
        RECT 1173.090 19.195 1173.370 19.565 ;
        RECT 91.700 2.400 91.840 19.195 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 91.630 19.240 91.910 19.520 ;
        RECT 1173.090 19.240 1173.370 19.520 ;
      LAYER met3 ;
        RECT 91.605 19.530 91.935 19.545 ;
        RECT 1173.065 19.530 1173.395 19.545 ;
        RECT 91.605 19.230 1173.395 19.530 ;
        RECT 91.605 19.215 91.935 19.230 ;
        RECT 1173.065 19.215 1173.395 19.230 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 0.300 ;
=======
      LAYER met1 ;
        RECT 941.690 1684.260 942.010 1684.320 ;
        RECT 1312.450 1684.260 1312.770 1684.320 ;
        RECT 941.690 1684.120 1312.770 1684.260 ;
        RECT 941.690 1684.060 942.010 1684.120 ;
        RECT 1312.450 1684.060 1312.770 1684.120 ;
        RECT 603.130 23.700 603.450 23.760 ;
        RECT 941.690 23.700 942.010 23.760 ;
        RECT 603.130 23.560 942.010 23.700 ;
        RECT 603.130 23.500 603.450 23.560 ;
        RECT 941.690 23.500 942.010 23.560 ;
      LAYER via ;
        RECT 941.720 1684.060 941.980 1684.320 ;
        RECT 1312.480 1684.060 1312.740 1684.320 ;
        RECT 603.160 23.500 603.420 23.760 ;
        RECT 941.720 23.500 941.980 23.760 ;
      LAYER met2 ;
        RECT 1312.470 1700.000 1312.750 1704.000 ;
        RECT 1312.540 1684.350 1312.680 1700.000 ;
        RECT 941.720 1684.030 941.980 1684.350 ;
        RECT 1312.480 1684.030 1312.740 1684.350 ;
        RECT 941.780 23.790 941.920 1684.030 ;
        RECT 603.160 23.470 603.420 23.790 ;
        RECT 941.720 23.470 941.980 23.790 ;
        RECT 603.220 2.400 603.360 23.470 ;
        RECT 603.010 -4.800 603.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 0.300 ;
=======
      LAYER met1 ;
        RECT 1312.910 1700.580 1313.230 1700.640 ;
        RECT 1316.130 1700.580 1316.450 1700.640 ;
        RECT 1312.910 1700.440 1316.450 1700.580 ;
        RECT 1312.910 1700.380 1313.230 1700.440 ;
        RECT 1316.130 1700.380 1316.450 1700.440 ;
        RECT 621.070 14.180 621.390 14.240 ;
        RECT 1312.910 14.180 1313.230 14.240 ;
        RECT 621.070 14.040 626.820 14.180 ;
        RECT 621.070 13.980 621.390 14.040 ;
        RECT 626.680 13.840 626.820 14.040 ;
        RECT 632.660 14.040 1313.230 14.180 ;
        RECT 632.660 13.840 632.800 14.040 ;
        RECT 1312.910 13.980 1313.230 14.040 ;
        RECT 626.680 13.700 632.800 13.840 ;
      LAYER via ;
        RECT 1312.940 1700.380 1313.200 1700.640 ;
        RECT 1316.160 1700.380 1316.420 1700.640 ;
        RECT 621.100 13.980 621.360 14.240 ;
        RECT 1312.940 13.980 1313.200 14.240 ;
      LAYER met2 ;
        RECT 1317.530 1701.090 1317.810 1704.000 ;
        RECT 1316.220 1700.950 1317.810 1701.090 ;
        RECT 1316.220 1700.670 1316.360 1700.950 ;
        RECT 1312.940 1700.350 1313.200 1700.670 ;
        RECT 1316.160 1700.350 1316.420 1700.670 ;
        RECT 1313.000 14.270 1313.140 1700.350 ;
        RECT 1317.530 1700.000 1317.810 1700.950 ;
        RECT 621.100 13.950 621.360 14.270 ;
        RECT 1312.940 13.950 1313.200 14.270 ;
        RECT 621.160 2.400 621.300 13.950 ;
        RECT 620.950 -4.800 621.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 0.300 ;
=======
      LAYER met1 ;
        RECT 115.530 17.580 115.850 17.640 ;
        RECT 115.530 17.440 1148.920 17.580 ;
        RECT 115.530 17.380 115.850 17.440 ;
        RECT 1148.780 17.240 1148.920 17.440 ;
        RECT 1179.510 17.240 1179.830 17.300 ;
        RECT 1148.780 17.100 1179.830 17.240 ;
        RECT 1179.510 17.040 1179.830 17.100 ;
      LAYER via ;
        RECT 115.560 17.380 115.820 17.640 ;
        RECT 1179.540 17.040 1179.800 17.300 ;
      LAYER met2 ;
        RECT 1180.910 1700.410 1181.190 1704.000 ;
        RECT 1180.060 1700.270 1181.190 1700.410 ;
        RECT 1180.060 17.920 1180.200 1700.270 ;
        RECT 1180.910 1700.000 1181.190 1700.270 ;
        RECT 1179.600 17.780 1180.200 17.920 ;
        RECT 115.560 17.350 115.820 17.670 ;
        RECT 115.620 2.400 115.760 17.350 ;
        RECT 1179.600 17.330 1179.740 17.780 ;
        RECT 1179.540 17.010 1179.800 17.330 ;
        RECT 115.410 -4.800 115.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 0.300 ;
=======
      LAYER li1 ;
        RECT 276.145 16.405 276.315 18.275 ;
        RECT 323.985 16.405 324.155 18.275 ;
        RECT 372.745 15.385 372.915 18.275 ;
        RECT 420.585 15.385 420.755 18.275 ;
        RECT 469.345 15.045 469.515 18.275 ;
        RECT 517.185 15.045 517.355 18.275 ;
        RECT 565.945 15.045 566.115 18.275 ;
        RECT 599.525 14.875 599.695 15.215 ;
        RECT 599.525 14.705 601.535 14.875 ;
        RECT 613.785 14.705 613.955 18.275 ;
        RECT 662.545 18.105 662.715 21.335 ;
        RECT 709.925 20.995 710.095 21.335 ;
        RECT 709.925 20.825 710.555 20.995 ;
        RECT 710.385 18.105 710.555 20.825 ;
        RECT 759.145 18.105 759.315 21.335 ;
        RECT 806.985 18.105 807.155 21.335 ;
        RECT 855.745 18.105 855.915 20.995 ;
        RECT 903.585 18.105 903.755 20.995 ;
        RECT 952.345 18.105 952.515 20.995 ;
        RECT 1000.185 18.105 1000.355 20.995 ;
        RECT 1048.945 18.105 1049.115 20.995 ;
        RECT 1096.785 18.105 1096.955 20.995 ;
      LAYER mcon ;
        RECT 662.545 21.165 662.715 21.335 ;
        RECT 709.925 21.165 710.095 21.335 ;
        RECT 759.145 21.165 759.315 21.335 ;
        RECT 276.145 18.105 276.315 18.275 ;
        RECT 323.985 18.105 324.155 18.275 ;
        RECT 372.745 18.105 372.915 18.275 ;
        RECT 420.585 18.105 420.755 18.275 ;
        RECT 469.345 18.105 469.515 18.275 ;
        RECT 517.185 18.105 517.355 18.275 ;
        RECT 565.945 18.105 566.115 18.275 ;
        RECT 613.785 18.105 613.955 18.275 ;
        RECT 806.985 21.165 807.155 21.335 ;
        RECT 855.745 20.825 855.915 20.995 ;
        RECT 903.585 20.825 903.755 20.995 ;
        RECT 952.345 20.825 952.515 20.995 ;
        RECT 1000.185 20.825 1000.355 20.995 ;
        RECT 1048.945 20.825 1049.115 20.995 ;
        RECT 1096.785 20.825 1096.955 20.995 ;
        RECT 599.525 15.045 599.695 15.215 ;
        RECT 601.365 14.705 601.535 14.875 ;
      LAYER met1 ;
        RECT 662.485 21.320 662.775 21.365 ;
        RECT 709.865 21.320 710.155 21.365 ;
        RECT 662.485 21.180 710.155 21.320 ;
        RECT 662.485 21.135 662.775 21.180 ;
        RECT 709.865 21.135 710.155 21.180 ;
        RECT 759.085 21.320 759.375 21.365 ;
        RECT 806.925 21.320 807.215 21.365 ;
        RECT 759.085 21.180 807.215 21.320 ;
        RECT 759.085 21.135 759.375 21.180 ;
        RECT 806.925 21.135 807.215 21.180 ;
        RECT 855.685 20.980 855.975 21.025 ;
        RECT 903.525 20.980 903.815 21.025 ;
        RECT 855.685 20.840 903.815 20.980 ;
        RECT 855.685 20.795 855.975 20.840 ;
        RECT 903.525 20.795 903.815 20.840 ;
        RECT 952.285 20.980 952.575 21.025 ;
        RECT 1000.125 20.980 1000.415 21.025 ;
        RECT 952.285 20.840 1000.415 20.980 ;
        RECT 952.285 20.795 952.575 20.840 ;
        RECT 1000.125 20.795 1000.415 20.840 ;
        RECT 1048.885 20.980 1049.175 21.025 ;
        RECT 1096.725 20.980 1097.015 21.025 ;
        RECT 1048.885 20.840 1097.015 20.980 ;
        RECT 1048.885 20.795 1049.175 20.840 ;
        RECT 1096.725 20.795 1097.015 20.840 ;
        RECT 139.450 18.260 139.770 18.320 ;
        RECT 276.085 18.260 276.375 18.305 ;
        RECT 139.450 18.120 276.375 18.260 ;
        RECT 139.450 18.060 139.770 18.120 ;
        RECT 276.085 18.075 276.375 18.120 ;
        RECT 323.925 18.260 324.215 18.305 ;
        RECT 372.685 18.260 372.975 18.305 ;
        RECT 323.925 18.120 372.975 18.260 ;
        RECT 323.925 18.075 324.215 18.120 ;
        RECT 372.685 18.075 372.975 18.120 ;
        RECT 420.525 18.260 420.815 18.305 ;
        RECT 469.285 18.260 469.575 18.305 ;
        RECT 420.525 18.120 469.575 18.260 ;
        RECT 420.525 18.075 420.815 18.120 ;
        RECT 469.285 18.075 469.575 18.120 ;
        RECT 517.125 18.260 517.415 18.305 ;
        RECT 565.885 18.260 566.175 18.305 ;
        RECT 517.125 18.120 566.175 18.260 ;
        RECT 517.125 18.075 517.415 18.120 ;
        RECT 565.885 18.075 566.175 18.120 ;
        RECT 613.725 18.260 614.015 18.305 ;
        RECT 662.485 18.260 662.775 18.305 ;
        RECT 613.725 18.120 662.775 18.260 ;
        RECT 613.725 18.075 614.015 18.120 ;
        RECT 662.485 18.075 662.775 18.120 ;
        RECT 710.325 18.260 710.615 18.305 ;
        RECT 759.085 18.260 759.375 18.305 ;
        RECT 710.325 18.120 759.375 18.260 ;
        RECT 710.325 18.075 710.615 18.120 ;
        RECT 759.085 18.075 759.375 18.120 ;
        RECT 806.925 18.260 807.215 18.305 ;
        RECT 855.685 18.260 855.975 18.305 ;
        RECT 806.925 18.120 855.975 18.260 ;
        RECT 806.925 18.075 807.215 18.120 ;
        RECT 855.685 18.075 855.975 18.120 ;
        RECT 903.525 18.260 903.815 18.305 ;
        RECT 952.285 18.260 952.575 18.305 ;
        RECT 903.525 18.120 952.575 18.260 ;
        RECT 903.525 18.075 903.815 18.120 ;
        RECT 952.285 18.075 952.575 18.120 ;
        RECT 1000.125 18.260 1000.415 18.305 ;
        RECT 1048.885 18.260 1049.175 18.305 ;
        RECT 1000.125 18.120 1049.175 18.260 ;
        RECT 1000.125 18.075 1000.415 18.120 ;
        RECT 1048.885 18.075 1049.175 18.120 ;
        RECT 1096.725 18.260 1097.015 18.305 ;
        RECT 1186.870 18.260 1187.190 18.320 ;
        RECT 1096.725 18.120 1187.190 18.260 ;
        RECT 1096.725 18.075 1097.015 18.120 ;
        RECT 1186.870 18.060 1187.190 18.120 ;
        RECT 276.085 16.560 276.375 16.605 ;
        RECT 323.925 16.560 324.215 16.605 ;
        RECT 276.085 16.420 324.215 16.560 ;
        RECT 276.085 16.375 276.375 16.420 ;
        RECT 323.925 16.375 324.215 16.420 ;
        RECT 372.685 15.540 372.975 15.585 ;
        RECT 420.525 15.540 420.815 15.585 ;
        RECT 372.685 15.400 420.815 15.540 ;
        RECT 372.685 15.355 372.975 15.400 ;
        RECT 420.525 15.355 420.815 15.400 ;
        RECT 469.285 15.200 469.575 15.245 ;
        RECT 517.125 15.200 517.415 15.245 ;
        RECT 469.285 15.060 517.415 15.200 ;
        RECT 469.285 15.015 469.575 15.060 ;
        RECT 517.125 15.015 517.415 15.060 ;
        RECT 565.885 15.200 566.175 15.245 ;
        RECT 599.465 15.200 599.755 15.245 ;
        RECT 565.885 15.060 599.755 15.200 ;
        RECT 565.885 15.015 566.175 15.060 ;
        RECT 599.465 15.015 599.755 15.060 ;
        RECT 601.305 14.860 601.595 14.905 ;
        RECT 613.725 14.860 614.015 14.905 ;
        RECT 601.305 14.720 614.015 14.860 ;
        RECT 601.305 14.675 601.595 14.720 ;
        RECT 613.725 14.675 614.015 14.720 ;
      LAYER via ;
        RECT 139.480 18.060 139.740 18.320 ;
        RECT 1186.900 18.060 1187.160 18.320 ;
      LAYER met2 ;
        RECT 1187.350 1700.410 1187.630 1704.000 ;
        RECT 1186.960 1700.270 1187.630 1700.410 ;
        RECT 1186.960 18.350 1187.100 1700.270 ;
        RECT 1187.350 1700.000 1187.630 1700.270 ;
        RECT 139.480 18.030 139.740 18.350 ;
        RECT 1186.900 18.030 1187.160 18.350 ;
        RECT 139.540 2.400 139.680 18.030 ;
        RECT 139.330 -4.800 139.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 157.270 -4.800 157.830 0.300 ;
=======
        RECT 1191.950 1700.000 1192.230 1704.000 ;
        RECT 1192.020 1688.965 1192.160 1700.000 ;
        RECT 158.330 1688.595 158.610 1688.965 ;
        RECT 1191.950 1688.595 1192.230 1688.965 ;
        RECT 158.400 17.410 158.540 1688.595 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 158.330 1688.640 158.610 1688.920 ;
        RECT 1191.950 1688.640 1192.230 1688.920 ;
      LAYER met3 ;
        RECT 158.305 1688.930 158.635 1688.945 ;
        RECT 1191.925 1688.930 1192.255 1688.945 ;
        RECT 158.305 1688.630 1192.255 1688.930 ;
        RECT 158.305 1688.615 158.635 1688.630 ;
        RECT 1191.925 1688.615 1192.255 1688.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1194.230 1693.440 1194.550 1693.500 ;
        RECT 1196.990 1693.440 1197.310 1693.500 ;
        RECT 1194.230 1693.300 1197.310 1693.440 ;
        RECT 1194.230 1693.240 1194.550 1693.300 ;
        RECT 1196.990 1693.240 1197.310 1693.300 ;
        RECT 174.870 18.940 175.190 19.000 ;
        RECT 1194.230 18.940 1194.550 19.000 ;
        RECT 174.870 18.800 1194.550 18.940 ;
        RECT 174.870 18.740 175.190 18.800 ;
        RECT 1194.230 18.740 1194.550 18.800 ;
      LAYER via ;
        RECT 1194.260 1693.240 1194.520 1693.500 ;
        RECT 1197.020 1693.240 1197.280 1693.500 ;
        RECT 174.900 18.740 175.160 19.000 ;
        RECT 1194.260 18.740 1194.520 19.000 ;
      LAYER met2 ;
        RECT 1197.010 1700.000 1197.290 1704.000 ;
        RECT 1197.080 1693.530 1197.220 1700.000 ;
        RECT 1194.260 1693.210 1194.520 1693.530 ;
        RECT 1197.020 1693.210 1197.280 1693.530 ;
        RECT 1194.320 19.030 1194.460 1693.210 ;
        RECT 174.900 18.710 175.160 19.030 ;
        RECT 1194.260 18.710 1194.520 19.030 ;
        RECT 174.960 2.400 175.100 18.710 ;
        RECT 174.750 -4.800 175.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1201.590 1687.320 1201.910 1687.380 ;
        RECT 1187.420 1687.180 1201.910 1687.320 ;
        RECT 192.810 1686.980 193.130 1687.040 ;
        RECT 1187.420 1686.980 1187.560 1687.180 ;
        RECT 1201.590 1687.120 1201.910 1687.180 ;
        RECT 192.810 1686.840 1187.560 1686.980 ;
        RECT 192.810 1686.780 193.130 1686.840 ;
      LAYER via ;
        RECT 192.840 1686.780 193.100 1687.040 ;
        RECT 1201.620 1687.120 1201.880 1687.380 ;
      LAYER met2 ;
        RECT 1201.610 1700.000 1201.890 1704.000 ;
        RECT 1201.680 1687.410 1201.820 1700.000 ;
        RECT 1201.620 1687.090 1201.880 1687.410 ;
        RECT 192.840 1686.750 193.100 1687.070 ;
        RECT 192.900 2.400 193.040 1686.750 ;
        RECT 192.690 -4.800 193.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 0.300 ;
=======
      LAYER li1 ;
        RECT 1201.665 786.505 1201.835 814.215 ;
        RECT 1201.665 524.365 1201.835 572.475 ;
        RECT 1202.125 276.165 1202.295 324.275 ;
        RECT 1202.125 179.605 1202.295 227.715 ;
        RECT 1202.125 65.365 1202.295 131.155 ;
      LAYER mcon ;
        RECT 1201.665 814.045 1201.835 814.215 ;
        RECT 1201.665 572.305 1201.835 572.475 ;
        RECT 1202.125 324.105 1202.295 324.275 ;
        RECT 1202.125 227.545 1202.295 227.715 ;
        RECT 1202.125 130.985 1202.295 131.155 ;
      LAYER met1 ;
        RECT 1202.050 1028.200 1202.370 1028.460 ;
        RECT 1202.140 1027.780 1202.280 1028.200 ;
        RECT 1202.050 1027.520 1202.370 1027.780 ;
        RECT 1202.510 1006.980 1202.830 1007.040 ;
        RECT 1204.350 1006.980 1204.670 1007.040 ;
        RECT 1202.510 1006.840 1204.670 1006.980 ;
        RECT 1202.510 1006.780 1202.830 1006.840 ;
        RECT 1204.350 1006.780 1204.670 1006.840 ;
        RECT 1202.050 869.420 1202.370 869.680 ;
        RECT 1202.140 868.940 1202.280 869.420 ;
        RECT 1202.510 868.940 1202.830 869.000 ;
        RECT 1202.140 868.800 1202.830 868.940 ;
        RECT 1202.510 868.740 1202.830 868.800 ;
        RECT 1201.590 845.480 1201.910 845.540 ;
        RECT 1202.510 845.480 1202.830 845.540 ;
        RECT 1201.590 845.340 1202.830 845.480 ;
        RECT 1201.590 845.280 1201.910 845.340 ;
        RECT 1202.510 845.280 1202.830 845.340 ;
        RECT 1201.590 814.200 1201.910 814.260 ;
        RECT 1201.395 814.060 1201.910 814.200 ;
        RECT 1201.590 814.000 1201.910 814.060 ;
        RECT 1201.590 786.660 1201.910 786.720 ;
        RECT 1201.395 786.520 1201.910 786.660 ;
        RECT 1201.590 786.460 1201.910 786.520 ;
        RECT 1201.605 572.460 1201.895 572.505 ;
        RECT 1202.050 572.460 1202.370 572.520 ;
        RECT 1201.605 572.320 1202.370 572.460 ;
        RECT 1201.605 572.275 1201.895 572.320 ;
        RECT 1202.050 572.260 1202.370 572.320 ;
        RECT 1201.590 524.520 1201.910 524.580 ;
        RECT 1201.395 524.380 1201.910 524.520 ;
        RECT 1201.590 524.320 1201.910 524.380 ;
        RECT 1201.590 427.620 1201.910 427.680 ;
        RECT 1202.050 427.620 1202.370 427.680 ;
        RECT 1201.590 427.480 1202.370 427.620 ;
        RECT 1201.590 427.420 1201.910 427.480 ;
        RECT 1202.050 427.420 1202.370 427.480 ;
        RECT 1201.590 331.060 1201.910 331.120 ;
        RECT 1202.050 331.060 1202.370 331.120 ;
        RECT 1201.590 330.920 1202.370 331.060 ;
        RECT 1201.590 330.860 1201.910 330.920 ;
        RECT 1202.050 330.860 1202.370 330.920 ;
        RECT 1202.050 324.260 1202.370 324.320 ;
        RECT 1201.855 324.120 1202.370 324.260 ;
        RECT 1202.050 324.060 1202.370 324.120 ;
        RECT 1202.050 276.320 1202.370 276.380 ;
        RECT 1201.855 276.180 1202.370 276.320 ;
        RECT 1202.050 276.120 1202.370 276.180 ;
        RECT 1201.590 234.300 1201.910 234.560 ;
        RECT 1201.680 234.160 1201.820 234.300 ;
        RECT 1202.050 234.160 1202.370 234.220 ;
        RECT 1201.680 234.020 1202.370 234.160 ;
        RECT 1202.050 233.960 1202.370 234.020 ;
        RECT 1202.050 227.700 1202.370 227.760 ;
        RECT 1201.855 227.560 1202.370 227.700 ;
        RECT 1202.050 227.500 1202.370 227.560 ;
        RECT 1202.050 179.760 1202.370 179.820 ;
        RECT 1201.855 179.620 1202.370 179.760 ;
        RECT 1202.050 179.560 1202.370 179.620 ;
        RECT 1201.590 131.140 1201.910 131.200 ;
        RECT 1202.065 131.140 1202.355 131.185 ;
        RECT 1201.590 131.000 1202.355 131.140 ;
        RECT 1201.590 130.940 1201.910 131.000 ;
        RECT 1202.065 130.955 1202.355 131.000 ;
        RECT 1202.065 65.520 1202.355 65.565 ;
        RECT 1202.970 65.520 1203.290 65.580 ;
        RECT 1202.065 65.380 1203.290 65.520 ;
        RECT 1202.065 65.335 1202.355 65.380 ;
        RECT 1202.970 65.320 1203.290 65.380 ;
        RECT 210.750 19.620 211.070 19.680 ;
        RECT 1201.590 19.620 1201.910 19.680 ;
        RECT 210.750 19.480 1201.910 19.620 ;
        RECT 210.750 19.420 211.070 19.480 ;
        RECT 1201.590 19.420 1201.910 19.480 ;
      LAYER via ;
        RECT 1202.080 1028.200 1202.340 1028.460 ;
        RECT 1202.080 1027.520 1202.340 1027.780 ;
        RECT 1202.540 1006.780 1202.800 1007.040 ;
        RECT 1204.380 1006.780 1204.640 1007.040 ;
        RECT 1202.080 869.420 1202.340 869.680 ;
        RECT 1202.540 868.740 1202.800 869.000 ;
        RECT 1201.620 845.280 1201.880 845.540 ;
        RECT 1202.540 845.280 1202.800 845.540 ;
        RECT 1201.620 814.000 1201.880 814.260 ;
        RECT 1201.620 786.460 1201.880 786.720 ;
        RECT 1202.080 572.260 1202.340 572.520 ;
        RECT 1201.620 524.320 1201.880 524.580 ;
        RECT 1201.620 427.420 1201.880 427.680 ;
        RECT 1202.080 427.420 1202.340 427.680 ;
        RECT 1201.620 330.860 1201.880 331.120 ;
        RECT 1202.080 330.860 1202.340 331.120 ;
        RECT 1202.080 324.060 1202.340 324.320 ;
        RECT 1202.080 276.120 1202.340 276.380 ;
        RECT 1201.620 234.300 1201.880 234.560 ;
        RECT 1202.080 233.960 1202.340 234.220 ;
        RECT 1202.080 227.500 1202.340 227.760 ;
        RECT 1202.080 179.560 1202.340 179.820 ;
        RECT 1201.620 130.940 1201.880 131.200 ;
        RECT 1203.000 65.320 1203.260 65.580 ;
        RECT 210.780 19.420 211.040 19.680 ;
        RECT 1201.620 19.420 1201.880 19.680 ;
      LAYER met2 ;
        RECT 1206.670 1700.410 1206.950 1704.000 ;
        RECT 1205.360 1700.270 1206.950 1700.410 ;
        RECT 1205.360 1677.290 1205.500 1700.270 ;
        RECT 1206.670 1700.000 1206.950 1700.270 ;
        RECT 1201.680 1677.150 1205.500 1677.290 ;
        RECT 1201.680 1655.530 1201.820 1677.150 ;
        RECT 1201.680 1655.390 1202.280 1655.530 ;
        RECT 1202.140 1511.370 1202.280 1655.390 ;
        RECT 1201.680 1511.230 1202.280 1511.370 ;
        RECT 1201.680 1510.690 1201.820 1511.230 ;
        RECT 1201.680 1510.550 1202.280 1510.690 ;
        RECT 1202.140 1414.810 1202.280 1510.550 ;
        RECT 1201.680 1414.670 1202.280 1414.810 ;
        RECT 1201.680 1414.130 1201.820 1414.670 ;
        RECT 1201.680 1413.990 1202.280 1414.130 ;
        RECT 1202.140 1318.250 1202.280 1413.990 ;
        RECT 1201.680 1318.110 1202.280 1318.250 ;
        RECT 1201.680 1317.570 1201.820 1318.110 ;
        RECT 1201.680 1317.430 1202.280 1317.570 ;
        RECT 1202.140 1221.690 1202.280 1317.430 ;
        RECT 1201.680 1221.550 1202.280 1221.690 ;
        RECT 1201.680 1221.010 1201.820 1221.550 ;
        RECT 1201.680 1220.870 1202.280 1221.010 ;
        RECT 1202.140 1125.130 1202.280 1220.870 ;
        RECT 1201.680 1124.990 1202.280 1125.130 ;
        RECT 1201.680 1124.450 1201.820 1124.990 ;
        RECT 1201.680 1124.310 1202.280 1124.450 ;
        RECT 1202.140 1028.490 1202.280 1124.310 ;
        RECT 1202.080 1028.170 1202.340 1028.490 ;
        RECT 1202.080 1027.490 1202.340 1027.810 ;
        RECT 1202.140 1014.290 1202.280 1027.490 ;
        RECT 1202.140 1014.150 1202.740 1014.290 ;
        RECT 1202.600 1007.070 1202.740 1014.150 ;
        RECT 1202.540 1006.750 1202.800 1007.070 ;
        RECT 1204.380 1006.750 1204.640 1007.070 ;
        RECT 1204.440 959.325 1204.580 1006.750 ;
        RECT 1203.450 958.955 1203.730 959.325 ;
        RECT 1204.370 958.955 1204.650 959.325 ;
        RECT 1203.520 911.045 1203.660 958.955 ;
        RECT 1202.070 910.675 1202.350 911.045 ;
        RECT 1203.450 910.675 1203.730 911.045 ;
        RECT 1202.140 869.710 1202.280 910.675 ;
        RECT 1202.080 869.390 1202.340 869.710 ;
        RECT 1202.540 868.710 1202.800 869.030 ;
        RECT 1202.600 845.570 1202.740 868.710 ;
        RECT 1201.620 845.250 1201.880 845.570 ;
        RECT 1202.540 845.250 1202.800 845.570 ;
        RECT 1201.680 814.290 1201.820 845.250 ;
        RECT 1201.620 813.970 1201.880 814.290 ;
        RECT 1201.620 786.430 1201.880 786.750 ;
        RECT 1201.680 700.810 1201.820 786.430 ;
        RECT 1201.680 700.670 1202.280 700.810 ;
        RECT 1202.140 628.845 1202.280 700.670 ;
        RECT 1202.070 628.475 1202.350 628.845 ;
        RECT 1201.610 627.795 1201.890 628.165 ;
        RECT 1201.680 596.770 1201.820 627.795 ;
        RECT 1201.680 596.630 1202.280 596.770 ;
        RECT 1202.140 572.550 1202.280 596.630 ;
        RECT 1202.080 572.230 1202.340 572.550 ;
        RECT 1201.620 524.290 1201.880 524.610 ;
        RECT 1201.680 476.240 1201.820 524.290 ;
        RECT 1201.680 476.100 1202.280 476.240 ;
        RECT 1202.140 435.725 1202.280 476.100 ;
        RECT 1202.070 435.355 1202.350 435.725 ;
        RECT 1201.610 434.675 1201.890 435.045 ;
        RECT 1201.680 427.710 1201.820 434.675 ;
        RECT 1201.620 427.390 1201.880 427.710 ;
        RECT 1202.080 427.390 1202.340 427.710 ;
        RECT 1202.140 379.680 1202.280 427.390 ;
        RECT 1202.140 379.540 1202.740 379.680 ;
        RECT 1202.600 331.570 1202.740 379.540 ;
        RECT 1201.680 331.430 1202.740 331.570 ;
        RECT 1201.680 331.150 1201.820 331.430 ;
        RECT 1201.620 330.830 1201.880 331.150 ;
        RECT 1202.080 330.830 1202.340 331.150 ;
        RECT 1202.140 324.350 1202.280 330.830 ;
        RECT 1202.080 324.030 1202.340 324.350 ;
        RECT 1202.080 276.090 1202.340 276.410 ;
        RECT 1202.140 258.810 1202.280 276.090 ;
        RECT 1201.680 258.670 1202.280 258.810 ;
        RECT 1201.680 234.590 1201.820 258.670 ;
        RECT 1201.620 234.270 1201.880 234.590 ;
        RECT 1202.080 233.930 1202.340 234.250 ;
        RECT 1202.140 227.790 1202.280 233.930 ;
        RECT 1202.080 227.470 1202.340 227.790 ;
        RECT 1202.080 179.530 1202.340 179.850 ;
        RECT 1202.140 138.450 1202.280 179.530 ;
        RECT 1201.680 138.310 1202.280 138.450 ;
        RECT 1201.680 131.230 1201.820 138.310 ;
        RECT 1201.620 130.910 1201.880 131.230 ;
        RECT 1203.000 65.290 1203.260 65.610 ;
        RECT 1203.060 42.005 1203.200 65.290 ;
        RECT 1202.070 41.635 1202.350 42.005 ;
        RECT 1202.990 41.635 1203.270 42.005 ;
        RECT 1202.140 41.210 1202.280 41.635 ;
        RECT 1201.680 41.070 1202.280 41.210 ;
        RECT 1201.680 19.710 1201.820 41.070 ;
        RECT 210.780 19.390 211.040 19.710 ;
        RECT 1201.620 19.390 1201.880 19.710 ;
        RECT 210.840 2.400 210.980 19.390 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 1203.450 959.000 1203.730 959.280 ;
        RECT 1204.370 959.000 1204.650 959.280 ;
        RECT 1202.070 910.720 1202.350 911.000 ;
        RECT 1203.450 910.720 1203.730 911.000 ;
        RECT 1202.070 628.520 1202.350 628.800 ;
        RECT 1201.610 627.840 1201.890 628.120 ;
        RECT 1202.070 435.400 1202.350 435.680 ;
        RECT 1201.610 434.720 1201.890 435.000 ;
        RECT 1202.070 41.680 1202.350 41.960 ;
        RECT 1202.990 41.680 1203.270 41.960 ;
      LAYER met3 ;
        RECT 1203.425 959.290 1203.755 959.305 ;
        RECT 1204.345 959.290 1204.675 959.305 ;
        RECT 1203.425 958.990 1204.675 959.290 ;
        RECT 1203.425 958.975 1203.755 958.990 ;
        RECT 1204.345 958.975 1204.675 958.990 ;
        RECT 1202.045 911.010 1202.375 911.025 ;
        RECT 1203.425 911.010 1203.755 911.025 ;
        RECT 1202.045 910.710 1203.755 911.010 ;
        RECT 1202.045 910.695 1202.375 910.710 ;
        RECT 1203.425 910.695 1203.755 910.710 ;
        RECT 1202.045 628.810 1202.375 628.825 ;
        RECT 1201.830 628.495 1202.375 628.810 ;
        RECT 1201.830 628.145 1202.130 628.495 ;
        RECT 1201.585 627.830 1202.130 628.145 ;
        RECT 1201.585 627.815 1201.915 627.830 ;
        RECT 1202.045 435.690 1202.375 435.705 ;
        RECT 1201.830 435.375 1202.375 435.690 ;
        RECT 1201.830 435.025 1202.130 435.375 ;
        RECT 1201.585 434.710 1202.130 435.025 ;
        RECT 1201.585 434.695 1201.915 434.710 ;
        RECT 1202.045 41.970 1202.375 41.985 ;
        RECT 1202.965 41.970 1203.295 41.985 ;
        RECT 1202.045 41.670 1203.295 41.970 ;
        RECT 1202.045 41.655 1202.375 41.670 ;
        RECT 1202.965 41.655 1203.295 41.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 0.300 ;
=======
      LAYER li1 ;
        RECT 1186.945 1687.165 1187.115 1689.035 ;
      LAYER mcon ;
        RECT 1186.945 1688.865 1187.115 1689.035 ;
      LAYER met1 ;
        RECT 1186.885 1689.020 1187.175 1689.065 ;
        RECT 1211.250 1689.020 1211.570 1689.080 ;
        RECT 1186.885 1688.880 1211.570 1689.020 ;
        RECT 1186.885 1688.835 1187.175 1688.880 ;
        RECT 1211.250 1688.820 1211.570 1688.880 ;
        RECT 234.210 1687.320 234.530 1687.380 ;
        RECT 1186.885 1687.320 1187.175 1687.365 ;
        RECT 234.210 1687.180 1187.175 1687.320 ;
        RECT 234.210 1687.120 234.530 1687.180 ;
        RECT 1186.885 1687.135 1187.175 1687.180 ;
        RECT 228.690 16.900 229.010 16.960 ;
        RECT 234.210 16.900 234.530 16.960 ;
        RECT 228.690 16.760 234.530 16.900 ;
        RECT 228.690 16.700 229.010 16.760 ;
        RECT 234.210 16.700 234.530 16.760 ;
      LAYER via ;
        RECT 1211.280 1688.820 1211.540 1689.080 ;
        RECT 234.240 1687.120 234.500 1687.380 ;
        RECT 228.720 16.700 228.980 16.960 ;
        RECT 234.240 16.700 234.500 16.960 ;
      LAYER met2 ;
        RECT 1211.270 1700.000 1211.550 1704.000 ;
        RECT 1211.340 1689.110 1211.480 1700.000 ;
        RECT 1211.280 1688.790 1211.540 1689.110 ;
        RECT 234.240 1687.090 234.500 1687.410 ;
        RECT 234.300 16.990 234.440 1687.090 ;
        RECT 228.720 16.670 228.980 16.990 ;
        RECT 234.240 16.670 234.500 16.990 ;
        RECT 228.780 2.400 228.920 16.670 ;
        RECT 228.570 -4.800 229.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 0.300 ;
=======
      LAYER li1 ;
        RECT 1162.105 1538.925 1162.275 1587.035 ;
        RECT 1161.185 1497.445 1161.355 1511.555 ;
        RECT 1161.185 1442.025 1161.355 1490.475 ;
        RECT 1161.645 966.365 1161.815 980.135 ;
        RECT 1161.645 303.365 1161.815 337.875 ;
      LAYER mcon ;
        RECT 1162.105 1586.865 1162.275 1587.035 ;
        RECT 1161.185 1511.385 1161.355 1511.555 ;
        RECT 1161.185 1490.305 1161.355 1490.475 ;
        RECT 1161.645 979.965 1161.815 980.135 ;
        RECT 1161.645 337.705 1161.815 337.875 ;
      LAYER met1 ;
        RECT 1161.570 1607.900 1161.890 1608.160 ;
        RECT 1161.660 1607.420 1161.800 1607.900 ;
        RECT 1162.030 1607.420 1162.350 1607.480 ;
        RECT 1161.660 1607.280 1162.350 1607.420 ;
        RECT 1162.030 1607.220 1162.350 1607.280 ;
        RECT 1162.045 1587.020 1162.335 1587.065 ;
        RECT 1162.490 1587.020 1162.810 1587.080 ;
        RECT 1162.045 1586.880 1162.810 1587.020 ;
        RECT 1162.045 1586.835 1162.335 1586.880 ;
        RECT 1162.490 1586.820 1162.810 1586.880 ;
        RECT 1162.030 1539.080 1162.350 1539.140 ;
        RECT 1161.835 1538.940 1162.350 1539.080 ;
        RECT 1162.030 1538.880 1162.350 1538.940 ;
        RECT 1161.125 1511.540 1161.415 1511.585 ;
        RECT 1162.030 1511.540 1162.350 1511.600 ;
        RECT 1161.125 1511.400 1162.350 1511.540 ;
        RECT 1161.125 1511.355 1161.415 1511.400 ;
        RECT 1162.030 1511.340 1162.350 1511.400 ;
        RECT 1161.110 1497.600 1161.430 1497.660 ;
        RECT 1160.915 1497.460 1161.430 1497.600 ;
        RECT 1161.110 1497.400 1161.430 1497.460 ;
        RECT 1161.110 1490.460 1161.430 1490.520 ;
        RECT 1160.915 1490.320 1161.430 1490.460 ;
        RECT 1161.110 1490.260 1161.430 1490.320 ;
        RECT 1161.125 1442.180 1161.415 1442.225 ;
        RECT 1162.490 1442.180 1162.810 1442.240 ;
        RECT 1161.125 1442.040 1162.810 1442.180 ;
        RECT 1161.125 1441.995 1161.415 1442.040 ;
        RECT 1162.490 1441.980 1162.810 1442.040 ;
        RECT 1162.030 1345.620 1162.350 1345.680 ;
        RECT 1162.490 1345.620 1162.810 1345.680 ;
        RECT 1162.030 1345.480 1162.810 1345.620 ;
        RECT 1162.030 1345.420 1162.350 1345.480 ;
        RECT 1162.490 1345.420 1162.810 1345.480 ;
        RECT 1161.570 1304.820 1161.890 1304.880 ;
        RECT 1162.030 1304.820 1162.350 1304.880 ;
        RECT 1161.570 1304.680 1162.350 1304.820 ;
        RECT 1161.570 1304.620 1161.890 1304.680 ;
        RECT 1162.030 1304.620 1162.350 1304.680 ;
        RECT 1161.570 1304.140 1161.890 1304.200 ;
        RECT 1162.030 1304.140 1162.350 1304.200 ;
        RECT 1161.570 1304.000 1162.350 1304.140 ;
        RECT 1161.570 1303.940 1161.890 1304.000 ;
        RECT 1162.030 1303.940 1162.350 1304.000 ;
        RECT 1161.570 1159.300 1161.890 1159.360 ;
        RECT 1162.030 1159.300 1162.350 1159.360 ;
        RECT 1161.570 1159.160 1162.350 1159.300 ;
        RECT 1161.570 1159.100 1161.890 1159.160 ;
        RECT 1162.030 1159.100 1162.350 1159.160 ;
        RECT 1161.570 1062.740 1161.890 1062.800 ;
        RECT 1162.030 1062.740 1162.350 1062.800 ;
        RECT 1161.570 1062.600 1162.350 1062.740 ;
        RECT 1161.570 1062.540 1161.890 1062.600 ;
        RECT 1162.030 1062.540 1162.350 1062.600 ;
        RECT 1161.570 980.120 1161.890 980.180 ;
        RECT 1161.375 979.980 1161.890 980.120 ;
        RECT 1161.570 979.920 1161.890 979.980 ;
        RECT 1161.570 966.520 1161.890 966.580 ;
        RECT 1161.375 966.380 1161.890 966.520 ;
        RECT 1161.570 966.320 1161.890 966.380 ;
        RECT 1161.570 931.980 1161.890 932.240 ;
        RECT 1161.660 931.560 1161.800 931.980 ;
        RECT 1161.570 931.300 1161.890 931.560 ;
        RECT 1161.570 869.620 1161.890 869.680 ;
        RECT 1162.030 869.620 1162.350 869.680 ;
        RECT 1161.570 869.480 1162.350 869.620 ;
        RECT 1161.570 869.420 1161.890 869.480 ;
        RECT 1162.030 869.420 1162.350 869.480 ;
        RECT 1161.110 786.660 1161.430 786.720 ;
        RECT 1162.030 786.660 1162.350 786.720 ;
        RECT 1161.110 786.520 1162.350 786.660 ;
        RECT 1161.110 786.460 1161.430 786.520 ;
        RECT 1162.030 786.460 1162.350 786.520 ;
        RECT 1161.570 689.900 1161.890 690.160 ;
        RECT 1161.660 689.760 1161.800 689.900 ;
        RECT 1162.030 689.760 1162.350 689.820 ;
        RECT 1161.660 689.620 1162.350 689.760 ;
        RECT 1162.030 689.560 1162.350 689.620 ;
        RECT 1161.570 593.340 1161.890 593.600 ;
        RECT 1161.660 593.200 1161.800 593.340 ;
        RECT 1162.030 593.200 1162.350 593.260 ;
        RECT 1161.660 593.060 1162.350 593.200 ;
        RECT 1162.030 593.000 1162.350 593.060 ;
        RECT 1161.570 517.380 1161.890 517.440 ;
        RECT 1162.030 517.380 1162.350 517.440 ;
        RECT 1161.570 517.240 1162.350 517.380 ;
        RECT 1161.570 517.180 1161.890 517.240 ;
        RECT 1162.030 517.180 1162.350 517.240 ;
        RECT 1161.570 337.860 1161.890 337.920 ;
        RECT 1161.375 337.720 1161.890 337.860 ;
        RECT 1161.570 337.660 1161.890 337.720 ;
        RECT 1161.570 303.520 1161.890 303.580 ;
        RECT 1161.375 303.380 1161.890 303.520 ;
        RECT 1161.570 303.320 1161.890 303.380 ;
      LAYER via ;
        RECT 1161.600 1607.900 1161.860 1608.160 ;
        RECT 1162.060 1607.220 1162.320 1607.480 ;
        RECT 1162.520 1586.820 1162.780 1587.080 ;
        RECT 1162.060 1538.880 1162.320 1539.140 ;
        RECT 1162.060 1511.340 1162.320 1511.600 ;
        RECT 1161.140 1497.400 1161.400 1497.660 ;
        RECT 1161.140 1490.260 1161.400 1490.520 ;
        RECT 1162.520 1441.980 1162.780 1442.240 ;
        RECT 1162.060 1345.420 1162.320 1345.680 ;
        RECT 1162.520 1345.420 1162.780 1345.680 ;
        RECT 1161.600 1304.620 1161.860 1304.880 ;
        RECT 1162.060 1304.620 1162.320 1304.880 ;
        RECT 1161.600 1303.940 1161.860 1304.200 ;
        RECT 1162.060 1303.940 1162.320 1304.200 ;
        RECT 1161.600 1159.100 1161.860 1159.360 ;
        RECT 1162.060 1159.100 1162.320 1159.360 ;
        RECT 1161.600 1062.540 1161.860 1062.800 ;
        RECT 1162.060 1062.540 1162.320 1062.800 ;
        RECT 1161.600 979.920 1161.860 980.180 ;
        RECT 1161.600 966.320 1161.860 966.580 ;
        RECT 1161.600 931.980 1161.860 932.240 ;
        RECT 1161.600 931.300 1161.860 931.560 ;
        RECT 1161.600 869.420 1161.860 869.680 ;
        RECT 1162.060 869.420 1162.320 869.680 ;
        RECT 1161.140 786.460 1161.400 786.720 ;
        RECT 1162.060 786.460 1162.320 786.720 ;
        RECT 1161.600 689.900 1161.860 690.160 ;
        RECT 1162.060 689.560 1162.320 689.820 ;
        RECT 1161.600 593.340 1161.860 593.600 ;
        RECT 1162.060 593.000 1162.320 593.260 ;
        RECT 1161.600 517.180 1161.860 517.440 ;
        RECT 1162.060 517.180 1162.320 517.440 ;
        RECT 1161.600 337.660 1161.860 337.920 ;
        RECT 1161.600 303.320 1161.860 303.580 ;
      LAYER met2 ;
        RECT 1162.970 1700.410 1163.250 1704.000 ;
        RECT 1162.580 1700.270 1163.250 1700.410 ;
        RECT 1162.580 1688.850 1162.720 1700.270 ;
        RECT 1162.970 1700.000 1163.250 1700.270 ;
        RECT 1161.660 1688.710 1162.720 1688.850 ;
        RECT 1161.660 1608.190 1161.800 1688.710 ;
        RECT 1161.600 1607.870 1161.860 1608.190 ;
        RECT 1162.060 1607.190 1162.320 1607.510 ;
        RECT 1162.120 1594.330 1162.260 1607.190 ;
        RECT 1162.120 1594.190 1162.720 1594.330 ;
        RECT 1162.580 1587.110 1162.720 1594.190 ;
        RECT 1162.520 1586.790 1162.780 1587.110 ;
        RECT 1162.060 1538.850 1162.320 1539.170 ;
        RECT 1162.120 1511.630 1162.260 1538.850 ;
        RECT 1162.060 1511.310 1162.320 1511.630 ;
        RECT 1161.140 1497.370 1161.400 1497.690 ;
        RECT 1161.200 1490.550 1161.340 1497.370 ;
        RECT 1161.140 1490.230 1161.400 1490.550 ;
        RECT 1162.520 1441.950 1162.780 1442.270 ;
        RECT 1162.580 1345.710 1162.720 1441.950 ;
        RECT 1162.060 1345.390 1162.320 1345.710 ;
        RECT 1162.520 1345.390 1162.780 1345.710 ;
        RECT 1162.120 1304.910 1162.260 1345.390 ;
        RECT 1161.600 1304.590 1161.860 1304.910 ;
        RECT 1162.060 1304.590 1162.320 1304.910 ;
        RECT 1161.660 1304.230 1161.800 1304.590 ;
        RECT 1161.600 1303.910 1161.860 1304.230 ;
        RECT 1162.060 1303.910 1162.320 1304.230 ;
        RECT 1162.120 1221.010 1162.260 1303.910 ;
        RECT 1161.660 1220.870 1162.260 1221.010 ;
        RECT 1161.660 1159.390 1161.800 1220.870 ;
        RECT 1161.600 1159.070 1161.860 1159.390 ;
        RECT 1162.060 1159.070 1162.320 1159.390 ;
        RECT 1162.120 1124.450 1162.260 1159.070 ;
        RECT 1161.660 1124.310 1162.260 1124.450 ;
        RECT 1161.660 1062.830 1161.800 1124.310 ;
        RECT 1161.600 1062.510 1161.860 1062.830 ;
        RECT 1162.060 1062.510 1162.320 1062.830 ;
        RECT 1162.120 1027.890 1162.260 1062.510 ;
        RECT 1161.660 1027.750 1162.260 1027.890 ;
        RECT 1161.660 980.210 1161.800 1027.750 ;
        RECT 1161.600 979.890 1161.860 980.210 ;
        RECT 1161.600 966.290 1161.860 966.610 ;
        RECT 1161.660 932.270 1161.800 966.290 ;
        RECT 1161.600 931.950 1161.860 932.270 ;
        RECT 1161.600 931.270 1161.860 931.590 ;
        RECT 1161.660 869.710 1161.800 931.270 ;
        RECT 1161.600 869.390 1161.860 869.710 ;
        RECT 1162.060 869.390 1162.320 869.710 ;
        RECT 1162.120 845.650 1162.260 869.390 ;
        RECT 1161.660 845.510 1162.260 845.650 ;
        RECT 1161.660 787.170 1161.800 845.510 ;
        RECT 1161.200 787.030 1161.800 787.170 ;
        RECT 1161.200 786.750 1161.340 787.030 ;
        RECT 1161.140 786.430 1161.400 786.750 ;
        RECT 1162.060 786.430 1162.320 786.750 ;
        RECT 1162.120 725.405 1162.260 786.430 ;
        RECT 1162.050 725.035 1162.330 725.405 ;
        RECT 1161.590 724.355 1161.870 724.725 ;
        RECT 1161.660 690.190 1161.800 724.355 ;
        RECT 1161.600 689.870 1161.860 690.190 ;
        RECT 1162.060 689.530 1162.320 689.850 ;
        RECT 1162.120 641.650 1162.260 689.530 ;
        RECT 1161.660 641.510 1162.260 641.650 ;
        RECT 1161.660 593.630 1161.800 641.510 ;
        RECT 1161.600 593.310 1161.860 593.630 ;
        RECT 1162.060 592.970 1162.320 593.290 ;
        RECT 1162.120 545.090 1162.260 592.970 ;
        RECT 1161.660 544.950 1162.260 545.090 ;
        RECT 1161.660 517.470 1161.800 544.950 ;
        RECT 1161.600 517.150 1161.860 517.470 ;
        RECT 1162.060 517.150 1162.320 517.470 ;
        RECT 1162.120 362.170 1162.260 517.150 ;
        RECT 1161.660 362.030 1162.260 362.170 ;
        RECT 1161.660 337.950 1161.800 362.030 ;
        RECT 1161.600 337.630 1161.860 337.950 ;
        RECT 1161.600 303.290 1161.860 303.610 ;
        RECT 1161.660 265.610 1161.800 303.290 ;
        RECT 1161.200 265.470 1161.800 265.610 ;
        RECT 1161.200 254.730 1161.340 265.470 ;
        RECT 1161.200 254.590 1162.260 254.730 ;
        RECT 1162.120 207.130 1162.260 254.590 ;
        RECT 1161.200 206.990 1162.260 207.130 ;
        RECT 1161.200 206.450 1161.340 206.990 ;
        RECT 1161.200 206.310 1161.800 206.450 ;
        RECT 1161.660 72.490 1161.800 206.310 ;
        RECT 1161.660 72.350 1162.260 72.490 ;
        RECT 1162.120 17.525 1162.260 72.350 ;
        RECT 50.230 17.155 50.510 17.525 ;
        RECT 1162.050 17.155 1162.330 17.525 ;
        RECT 50.300 2.400 50.440 17.155 ;
        RECT 50.090 -4.800 50.650 2.400 ;
      LAYER via2 ;
        RECT 1162.050 725.080 1162.330 725.360 ;
        RECT 1161.590 724.400 1161.870 724.680 ;
        RECT 50.230 17.200 50.510 17.480 ;
        RECT 1162.050 17.200 1162.330 17.480 ;
      LAYER met3 ;
        RECT 1162.025 725.370 1162.355 725.385 ;
        RECT 1161.350 725.070 1162.355 725.370 ;
        RECT 1161.350 724.705 1161.650 725.070 ;
        RECT 1162.025 725.055 1162.355 725.070 ;
        RECT 1161.350 724.390 1161.895 724.705 ;
        RECT 1161.565 724.375 1161.895 724.390 ;
        RECT 50.205 17.490 50.535 17.505 ;
        RECT 1162.025 17.490 1162.355 17.505 ;
        RECT 50.205 17.190 1162.355 17.490 ;
        RECT 50.205 17.175 50.535 17.190 ;
        RECT 1162.025 17.175 1162.355 17.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 0.300 ;
=======
      LAYER li1 ;
        RECT 1177.285 1688.185 1177.455 1690.735 ;
        RECT 1197.525 1689.205 1197.695 1690.735 ;
      LAYER mcon ;
        RECT 1177.285 1690.565 1177.455 1690.735 ;
        RECT 1197.525 1690.565 1197.695 1690.735 ;
      LAYER met1 ;
        RECT 1177.225 1690.720 1177.515 1690.765 ;
        RECT 1197.465 1690.720 1197.755 1690.765 ;
        RECT 1177.225 1690.580 1197.755 1690.720 ;
        RECT 1177.225 1690.535 1177.515 1690.580 ;
        RECT 1197.465 1690.535 1197.755 1690.580 ;
        RECT 1197.465 1689.360 1197.755 1689.405 ;
        RECT 1217.690 1689.360 1218.010 1689.420 ;
        RECT 1197.465 1689.220 1218.010 1689.360 ;
        RECT 1197.465 1689.175 1197.755 1689.220 ;
        RECT 1217.690 1689.160 1218.010 1689.220 ;
        RECT 254.910 1688.340 255.230 1688.400 ;
        RECT 1177.225 1688.340 1177.515 1688.385 ;
        RECT 254.910 1688.200 1177.515 1688.340 ;
        RECT 254.910 1688.140 255.230 1688.200 ;
        RECT 1177.225 1688.155 1177.515 1688.200 ;
        RECT 252.610 16.900 252.930 16.960 ;
        RECT 254.910 16.900 255.230 16.960 ;
        RECT 252.610 16.760 255.230 16.900 ;
        RECT 252.610 16.700 252.930 16.760 ;
        RECT 254.910 16.700 255.230 16.760 ;
      LAYER via ;
        RECT 1217.720 1689.160 1217.980 1689.420 ;
        RECT 254.940 1688.140 255.200 1688.400 ;
        RECT 252.640 16.700 252.900 16.960 ;
        RECT 254.940 16.700 255.200 16.960 ;
      LAYER met2 ;
        RECT 1217.710 1700.000 1217.990 1704.000 ;
        RECT 1217.780 1689.450 1217.920 1700.000 ;
        RECT 1217.720 1689.130 1217.980 1689.450 ;
        RECT 254.940 1688.110 255.200 1688.430 ;
        RECT 255.000 16.990 255.140 1688.110 ;
        RECT 252.640 16.670 252.900 16.990 ;
        RECT 254.940 16.670 255.200 16.990 ;
        RECT 252.700 2.400 252.840 16.670 ;
        RECT 252.490 -4.800 253.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 0.300 ;
=======
      LAYER li1 ;
        RECT 1222.825 1573.265 1222.995 1683.595 ;
        RECT 1222.825 1490.645 1222.995 1538.755 ;
        RECT 1222.825 1255.365 1222.995 1283.415 ;
        RECT 1222.825 966.025 1222.995 1025.015 ;
        RECT 1223.285 821.185 1223.455 845.495 ;
        RECT 1222.825 331.245 1222.995 379.355 ;
      LAYER mcon ;
        RECT 1222.825 1683.425 1222.995 1683.595 ;
        RECT 1222.825 1538.585 1222.995 1538.755 ;
        RECT 1222.825 1283.245 1222.995 1283.415 ;
        RECT 1222.825 1024.845 1222.995 1025.015 ;
        RECT 1223.285 845.325 1223.455 845.495 ;
        RECT 1222.825 379.185 1222.995 379.355 ;
      LAYER met1 ;
        RECT 1222.750 1683.580 1223.070 1683.640 ;
        RECT 1222.555 1683.440 1223.070 1683.580 ;
        RECT 1222.750 1683.380 1223.070 1683.440 ;
        RECT 1222.765 1573.420 1223.055 1573.465 ;
        RECT 1223.210 1573.420 1223.530 1573.480 ;
        RECT 1222.765 1573.280 1223.530 1573.420 ;
        RECT 1222.765 1573.235 1223.055 1573.280 ;
        RECT 1223.210 1573.220 1223.530 1573.280 ;
        RECT 1222.765 1538.740 1223.055 1538.785 ;
        RECT 1223.210 1538.740 1223.530 1538.800 ;
        RECT 1222.765 1538.600 1223.530 1538.740 ;
        RECT 1222.765 1538.555 1223.055 1538.600 ;
        RECT 1223.210 1538.540 1223.530 1538.600 ;
        RECT 1222.750 1490.800 1223.070 1490.860 ;
        RECT 1222.555 1490.660 1223.070 1490.800 ;
        RECT 1222.750 1490.600 1223.070 1490.660 ;
        RECT 1222.750 1462.720 1223.070 1462.980 ;
        RECT 1222.840 1462.240 1222.980 1462.720 ;
        RECT 1223.210 1462.240 1223.530 1462.300 ;
        RECT 1222.840 1462.100 1223.530 1462.240 ;
        RECT 1223.210 1462.040 1223.530 1462.100 ;
        RECT 1223.210 1404.100 1223.530 1404.160 ;
        RECT 1224.130 1404.100 1224.450 1404.160 ;
        RECT 1223.210 1403.960 1224.450 1404.100 ;
        RECT 1223.210 1403.900 1223.530 1403.960 ;
        RECT 1224.130 1403.900 1224.450 1403.960 ;
        RECT 1223.210 1338.820 1223.530 1338.880 ;
        RECT 1222.840 1338.680 1223.530 1338.820 ;
        RECT 1222.840 1338.540 1222.980 1338.680 ;
        RECT 1223.210 1338.620 1223.530 1338.680 ;
        RECT 1222.750 1338.280 1223.070 1338.540 ;
        RECT 1222.750 1331.680 1223.070 1331.740 ;
        RECT 1223.670 1331.680 1223.990 1331.740 ;
        RECT 1222.750 1331.540 1223.990 1331.680 ;
        RECT 1222.750 1331.480 1223.070 1331.540 ;
        RECT 1223.670 1331.480 1223.990 1331.540 ;
        RECT 1222.750 1283.400 1223.070 1283.460 ;
        RECT 1222.555 1283.260 1223.070 1283.400 ;
        RECT 1222.750 1283.200 1223.070 1283.260 ;
        RECT 1222.765 1255.520 1223.055 1255.565 ;
        RECT 1223.670 1255.520 1223.990 1255.580 ;
        RECT 1222.765 1255.380 1223.990 1255.520 ;
        RECT 1222.765 1255.335 1223.055 1255.380 ;
        RECT 1223.670 1255.320 1223.990 1255.380 ;
        RECT 1223.210 1159.300 1223.530 1159.360 ;
        RECT 1223.670 1159.300 1223.990 1159.360 ;
        RECT 1223.210 1159.160 1223.990 1159.300 ;
        RECT 1223.210 1159.100 1223.530 1159.160 ;
        RECT 1223.670 1159.100 1223.990 1159.160 ;
        RECT 1222.750 1104.220 1223.070 1104.280 ;
        RECT 1224.130 1104.220 1224.450 1104.280 ;
        RECT 1222.750 1104.080 1224.450 1104.220 ;
        RECT 1222.750 1104.020 1223.070 1104.080 ;
        RECT 1224.130 1104.020 1224.450 1104.080 ;
        RECT 1222.750 1103.540 1223.070 1103.600 ;
        RECT 1224.130 1103.540 1224.450 1103.600 ;
        RECT 1222.750 1103.400 1224.450 1103.540 ;
        RECT 1222.750 1103.340 1223.070 1103.400 ;
        RECT 1224.130 1103.340 1224.450 1103.400 ;
        RECT 1222.765 1025.000 1223.055 1025.045 ;
        RECT 1223.670 1025.000 1223.990 1025.060 ;
        RECT 1222.765 1024.860 1223.990 1025.000 ;
        RECT 1222.765 1024.815 1223.055 1024.860 ;
        RECT 1223.670 1024.800 1223.990 1024.860 ;
        RECT 1222.765 966.180 1223.055 966.225 ;
        RECT 1223.210 966.180 1223.530 966.240 ;
        RECT 1222.765 966.040 1223.530 966.180 ;
        RECT 1222.765 965.995 1223.055 966.040 ;
        RECT 1223.210 965.980 1223.530 966.040 ;
        RECT 1222.750 917.900 1223.070 917.960 ;
        RECT 1224.130 917.900 1224.450 917.960 ;
        RECT 1222.750 917.760 1224.450 917.900 ;
        RECT 1222.750 917.700 1223.070 917.760 ;
        RECT 1224.130 917.700 1224.450 917.760 ;
        RECT 1222.750 869.620 1223.070 869.680 ;
        RECT 1223.210 869.620 1223.530 869.680 ;
        RECT 1222.750 869.480 1223.530 869.620 ;
        RECT 1222.750 869.420 1223.070 869.480 ;
        RECT 1223.210 869.420 1223.530 869.480 ;
        RECT 1223.210 845.480 1223.530 845.540 ;
        RECT 1223.015 845.340 1223.530 845.480 ;
        RECT 1223.210 845.280 1223.530 845.340 ;
        RECT 1223.225 821.340 1223.515 821.385 ;
        RECT 1223.670 821.340 1223.990 821.400 ;
        RECT 1223.225 821.200 1223.990 821.340 ;
        RECT 1223.225 821.155 1223.515 821.200 ;
        RECT 1223.670 821.140 1223.990 821.200 ;
        RECT 1222.750 724.440 1223.070 724.500 ;
        RECT 1223.670 724.440 1223.990 724.500 ;
        RECT 1222.750 724.300 1223.990 724.440 ;
        RECT 1222.750 724.240 1223.070 724.300 ;
        RECT 1223.670 724.240 1223.990 724.300 ;
        RECT 1222.750 531.320 1223.070 531.380 ;
        RECT 1223.670 531.320 1223.990 531.380 ;
        RECT 1222.750 531.180 1223.990 531.320 ;
        RECT 1222.750 531.120 1223.070 531.180 ;
        RECT 1223.670 531.120 1223.990 531.180 ;
        RECT 1222.750 434.560 1223.070 434.820 ;
        RECT 1222.840 434.420 1222.980 434.560 ;
        RECT 1223.210 434.420 1223.530 434.480 ;
        RECT 1222.840 434.280 1223.530 434.420 ;
        RECT 1223.210 434.220 1223.530 434.280 ;
        RECT 1222.765 379.340 1223.055 379.385 ;
        RECT 1223.210 379.340 1223.530 379.400 ;
        RECT 1222.765 379.200 1223.530 379.340 ;
        RECT 1222.765 379.155 1223.055 379.200 ;
        RECT 1223.210 379.140 1223.530 379.200 ;
        RECT 1222.750 331.400 1223.070 331.460 ;
        RECT 1222.555 331.260 1223.070 331.400 ;
        RECT 1222.750 331.200 1223.070 331.260 ;
        RECT 1223.210 241.980 1223.530 242.040 ;
        RECT 1222.840 241.840 1223.530 241.980 ;
        RECT 1222.840 241.700 1222.980 241.840 ;
        RECT 1223.210 241.780 1223.530 241.840 ;
        RECT 1222.750 241.440 1223.070 241.700 ;
        RECT 1222.750 186.560 1223.070 186.620 ;
        RECT 1223.210 186.560 1223.530 186.620 ;
        RECT 1222.750 186.420 1223.530 186.560 ;
        RECT 1222.750 186.360 1223.070 186.420 ;
        RECT 1223.210 186.360 1223.530 186.420 ;
        RECT 1223.210 158.820 1223.530 159.080 ;
        RECT 1223.300 158.400 1223.440 158.820 ;
        RECT 1223.210 158.140 1223.530 158.400 ;
        RECT 270.090 20.300 270.410 20.360 ;
        RECT 1223.210 20.300 1223.530 20.360 ;
        RECT 270.090 20.160 1223.530 20.300 ;
        RECT 270.090 20.100 270.410 20.160 ;
        RECT 1223.210 20.100 1223.530 20.160 ;
      LAYER via ;
        RECT 1222.780 1683.380 1223.040 1683.640 ;
        RECT 1223.240 1573.220 1223.500 1573.480 ;
        RECT 1223.240 1538.540 1223.500 1538.800 ;
        RECT 1222.780 1490.600 1223.040 1490.860 ;
        RECT 1222.780 1462.720 1223.040 1462.980 ;
        RECT 1223.240 1462.040 1223.500 1462.300 ;
        RECT 1223.240 1403.900 1223.500 1404.160 ;
        RECT 1224.160 1403.900 1224.420 1404.160 ;
        RECT 1223.240 1338.620 1223.500 1338.880 ;
        RECT 1222.780 1338.280 1223.040 1338.540 ;
        RECT 1222.780 1331.480 1223.040 1331.740 ;
        RECT 1223.700 1331.480 1223.960 1331.740 ;
        RECT 1222.780 1283.200 1223.040 1283.460 ;
        RECT 1223.700 1255.320 1223.960 1255.580 ;
        RECT 1223.240 1159.100 1223.500 1159.360 ;
        RECT 1223.700 1159.100 1223.960 1159.360 ;
        RECT 1222.780 1104.020 1223.040 1104.280 ;
        RECT 1224.160 1104.020 1224.420 1104.280 ;
        RECT 1222.780 1103.340 1223.040 1103.600 ;
        RECT 1224.160 1103.340 1224.420 1103.600 ;
        RECT 1223.700 1024.800 1223.960 1025.060 ;
        RECT 1223.240 965.980 1223.500 966.240 ;
        RECT 1222.780 917.700 1223.040 917.960 ;
        RECT 1224.160 917.700 1224.420 917.960 ;
        RECT 1222.780 869.420 1223.040 869.680 ;
        RECT 1223.240 869.420 1223.500 869.680 ;
        RECT 1223.240 845.280 1223.500 845.540 ;
        RECT 1223.700 821.140 1223.960 821.400 ;
        RECT 1222.780 724.240 1223.040 724.500 ;
        RECT 1223.700 724.240 1223.960 724.500 ;
        RECT 1222.780 531.120 1223.040 531.380 ;
        RECT 1223.700 531.120 1223.960 531.380 ;
        RECT 1222.780 434.560 1223.040 434.820 ;
        RECT 1223.240 434.220 1223.500 434.480 ;
        RECT 1223.240 379.140 1223.500 379.400 ;
        RECT 1222.780 331.200 1223.040 331.460 ;
        RECT 1223.240 241.780 1223.500 242.040 ;
        RECT 1222.780 241.440 1223.040 241.700 ;
        RECT 1222.780 186.360 1223.040 186.620 ;
        RECT 1223.240 186.360 1223.500 186.620 ;
        RECT 1223.240 158.820 1223.500 159.080 ;
        RECT 1223.240 158.140 1223.500 158.400 ;
        RECT 270.120 20.100 270.380 20.360 ;
        RECT 1223.240 20.100 1223.500 20.360 ;
      LAYER met2 ;
        RECT 1222.770 1700.000 1223.050 1704.000 ;
        RECT 1222.840 1683.670 1222.980 1700.000 ;
        RECT 1222.780 1683.350 1223.040 1683.670 ;
        RECT 1223.240 1573.190 1223.500 1573.510 ;
        RECT 1223.300 1538.830 1223.440 1573.190 ;
        RECT 1223.240 1538.510 1223.500 1538.830 ;
        RECT 1222.780 1490.570 1223.040 1490.890 ;
        RECT 1222.840 1463.010 1222.980 1490.570 ;
        RECT 1222.780 1462.690 1223.040 1463.010 ;
        RECT 1223.240 1462.010 1223.500 1462.330 ;
        RECT 1223.300 1404.190 1223.440 1462.010 ;
        RECT 1223.240 1403.870 1223.500 1404.190 ;
        RECT 1224.160 1403.870 1224.420 1404.190 ;
        RECT 1224.220 1380.245 1224.360 1403.870 ;
        RECT 1223.230 1379.875 1223.510 1380.245 ;
        RECT 1224.150 1379.875 1224.430 1380.245 ;
        RECT 1223.300 1338.910 1223.440 1379.875 ;
        RECT 1223.240 1338.590 1223.500 1338.910 ;
        RECT 1222.780 1338.250 1223.040 1338.570 ;
        RECT 1222.840 1331.770 1222.980 1338.250 ;
        RECT 1222.780 1331.450 1223.040 1331.770 ;
        RECT 1223.700 1331.450 1223.960 1331.770 ;
        RECT 1223.760 1283.685 1223.900 1331.450 ;
        RECT 1222.770 1283.315 1223.050 1283.685 ;
        RECT 1223.690 1283.315 1223.970 1283.685 ;
        RECT 1222.780 1283.170 1223.040 1283.315 ;
        RECT 1223.700 1255.290 1223.960 1255.610 ;
        RECT 1223.760 1159.390 1223.900 1255.290 ;
        RECT 1223.240 1159.070 1223.500 1159.390 ;
        RECT 1223.700 1159.070 1223.960 1159.390 ;
        RECT 1223.300 1152.445 1223.440 1159.070 ;
        RECT 1223.230 1152.075 1223.510 1152.445 ;
        RECT 1224.150 1152.075 1224.430 1152.445 ;
        RECT 1224.220 1104.310 1224.360 1152.075 ;
        RECT 1222.780 1103.990 1223.040 1104.310 ;
        RECT 1224.160 1103.990 1224.420 1104.310 ;
        RECT 1222.840 1103.630 1222.980 1103.990 ;
        RECT 1222.780 1103.310 1223.040 1103.630 ;
        RECT 1224.160 1103.310 1224.420 1103.630 ;
        RECT 1224.220 1062.570 1224.360 1103.310 ;
        RECT 1223.760 1062.430 1224.360 1062.570 ;
        RECT 1223.760 1025.090 1223.900 1062.430 ;
        RECT 1223.700 1024.770 1223.960 1025.090 ;
        RECT 1223.240 966.125 1223.500 966.270 ;
        RECT 1223.230 965.755 1223.510 966.125 ;
        RECT 1224.150 965.755 1224.430 966.125 ;
        RECT 1224.220 917.990 1224.360 965.755 ;
        RECT 1222.780 917.670 1223.040 917.990 ;
        RECT 1224.160 917.670 1224.420 917.990 ;
        RECT 1222.840 869.710 1222.980 917.670 ;
        RECT 1222.780 869.390 1223.040 869.710 ;
        RECT 1223.240 869.390 1223.500 869.710 ;
        RECT 1223.300 845.570 1223.440 869.390 ;
        RECT 1223.240 845.250 1223.500 845.570 ;
        RECT 1223.700 821.110 1223.960 821.430 ;
        RECT 1223.760 766.090 1223.900 821.110 ;
        RECT 1223.300 765.950 1223.900 766.090 ;
        RECT 1223.300 724.610 1223.440 765.950 ;
        RECT 1222.840 724.530 1223.440 724.610 ;
        RECT 1222.780 724.470 1223.440 724.530 ;
        RECT 1222.780 724.210 1223.040 724.470 ;
        RECT 1223.700 724.210 1223.960 724.530 ;
        RECT 1223.760 688.570 1223.900 724.210 ;
        RECT 1223.300 688.430 1223.900 688.570 ;
        RECT 1223.300 651.850 1223.440 688.430 ;
        RECT 1222.840 651.710 1223.440 651.850 ;
        RECT 1222.840 531.410 1222.980 651.710 ;
        RECT 1222.780 531.090 1223.040 531.410 ;
        RECT 1223.700 531.090 1223.960 531.410 ;
        RECT 1223.760 495.450 1223.900 531.090 ;
        RECT 1223.300 495.310 1223.900 495.450 ;
        RECT 1223.300 458.730 1223.440 495.310 ;
        RECT 1222.840 458.590 1223.440 458.730 ;
        RECT 1222.840 434.850 1222.980 458.590 ;
        RECT 1222.780 434.530 1223.040 434.850 ;
        RECT 1223.240 434.190 1223.500 434.510 ;
        RECT 1223.300 379.430 1223.440 434.190 ;
        RECT 1223.240 379.110 1223.500 379.430 ;
        RECT 1222.780 331.170 1223.040 331.490 ;
        RECT 1222.840 331.005 1222.980 331.170 ;
        RECT 1222.770 330.635 1223.050 331.005 ;
        RECT 1223.230 329.955 1223.510 330.325 ;
        RECT 1223.300 242.070 1223.440 329.955 ;
        RECT 1223.240 241.750 1223.500 242.070 ;
        RECT 1222.780 241.410 1223.040 241.730 ;
        RECT 1222.840 186.650 1222.980 241.410 ;
        RECT 1222.780 186.330 1223.040 186.650 ;
        RECT 1223.240 186.330 1223.500 186.650 ;
        RECT 1223.300 159.110 1223.440 186.330 ;
        RECT 1223.240 158.790 1223.500 159.110 ;
        RECT 1223.240 158.110 1223.500 158.430 ;
        RECT 1223.300 20.390 1223.440 158.110 ;
        RECT 270.120 20.070 270.380 20.390 ;
        RECT 1223.240 20.070 1223.500 20.390 ;
        RECT 270.180 2.400 270.320 20.070 ;
        RECT 269.970 -4.800 270.530 2.400 ;
      LAYER via2 ;
        RECT 1223.230 1379.920 1223.510 1380.200 ;
        RECT 1224.150 1379.920 1224.430 1380.200 ;
        RECT 1222.770 1283.360 1223.050 1283.640 ;
        RECT 1223.690 1283.360 1223.970 1283.640 ;
        RECT 1223.230 1152.120 1223.510 1152.400 ;
        RECT 1224.150 1152.120 1224.430 1152.400 ;
        RECT 1223.230 965.800 1223.510 966.080 ;
        RECT 1224.150 965.800 1224.430 966.080 ;
        RECT 1222.770 330.680 1223.050 330.960 ;
        RECT 1223.230 330.000 1223.510 330.280 ;
      LAYER met3 ;
        RECT 1223.205 1380.210 1223.535 1380.225 ;
        RECT 1224.125 1380.210 1224.455 1380.225 ;
        RECT 1223.205 1379.910 1224.455 1380.210 ;
        RECT 1223.205 1379.895 1223.535 1379.910 ;
        RECT 1224.125 1379.895 1224.455 1379.910 ;
        RECT 1222.745 1283.650 1223.075 1283.665 ;
        RECT 1223.665 1283.650 1223.995 1283.665 ;
        RECT 1222.745 1283.350 1223.995 1283.650 ;
        RECT 1222.745 1283.335 1223.075 1283.350 ;
        RECT 1223.665 1283.335 1223.995 1283.350 ;
        RECT 1223.205 1152.410 1223.535 1152.425 ;
        RECT 1224.125 1152.410 1224.455 1152.425 ;
        RECT 1223.205 1152.110 1224.455 1152.410 ;
        RECT 1223.205 1152.095 1223.535 1152.110 ;
        RECT 1224.125 1152.095 1224.455 1152.110 ;
        RECT 1223.205 966.090 1223.535 966.105 ;
        RECT 1224.125 966.090 1224.455 966.105 ;
        RECT 1223.205 965.790 1224.455 966.090 ;
        RECT 1223.205 965.775 1223.535 965.790 ;
        RECT 1224.125 965.775 1224.455 965.790 ;
        RECT 1222.745 330.970 1223.075 330.985 ;
        RECT 1222.070 330.670 1223.075 330.970 ;
        RECT 1222.070 330.290 1222.370 330.670 ;
        RECT 1222.745 330.655 1223.075 330.670 ;
        RECT 1223.205 330.290 1223.535 330.305 ;
        RECT 1222.070 329.990 1223.535 330.290 ;
        RECT 1223.205 329.975 1223.535 329.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 0.300 ;
=======
      LAYER met1 ;
        RECT 1227.350 1689.360 1227.670 1689.420 ;
        RECT 1218.240 1689.220 1227.670 1689.360 ;
        RECT 289.410 1688.680 289.730 1688.740 ;
        RECT 1218.240 1688.680 1218.380 1689.220 ;
        RECT 1227.350 1689.160 1227.670 1689.220 ;
        RECT 289.410 1688.540 1218.380 1688.680 ;
        RECT 289.410 1688.480 289.730 1688.540 ;
      LAYER via ;
        RECT 289.440 1688.480 289.700 1688.740 ;
        RECT 1227.380 1689.160 1227.640 1689.420 ;
      LAYER met2 ;
        RECT 1227.370 1700.000 1227.650 1704.000 ;
        RECT 1227.440 1689.450 1227.580 1700.000 ;
        RECT 1227.380 1689.130 1227.640 1689.450 ;
        RECT 289.440 1688.450 289.700 1688.770 ;
        RECT 289.500 17.410 289.640 1688.450 ;
        RECT 288.120 17.270 289.640 17.410 ;
        RECT 288.120 2.400 288.260 17.270 ;
        RECT 287.910 -4.800 288.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 0.300 ;
=======
      LAYER li1 ;
        RECT 1178.665 1687.505 1178.835 1689.035 ;
      LAYER mcon ;
        RECT 1178.665 1688.865 1178.835 1689.035 ;
      LAYER met1 ;
        RECT 310.110 1689.020 310.430 1689.080 ;
        RECT 1178.605 1689.020 1178.895 1689.065 ;
        RECT 310.110 1688.880 1178.895 1689.020 ;
        RECT 310.110 1688.820 310.430 1688.880 ;
        RECT 1178.605 1688.835 1178.895 1688.880 ;
        RECT 1178.605 1687.660 1178.895 1687.705 ;
        RECT 1232.410 1687.660 1232.730 1687.720 ;
        RECT 1178.605 1687.520 1232.730 1687.660 ;
        RECT 1178.605 1687.475 1178.895 1687.520 ;
        RECT 1232.410 1687.460 1232.730 1687.520 ;
        RECT 305.970 16.900 306.290 16.960 ;
        RECT 310.110 16.900 310.430 16.960 ;
        RECT 305.970 16.760 310.430 16.900 ;
        RECT 305.970 16.700 306.290 16.760 ;
        RECT 310.110 16.700 310.430 16.760 ;
      LAYER via ;
        RECT 310.140 1688.820 310.400 1689.080 ;
        RECT 1232.440 1687.460 1232.700 1687.720 ;
        RECT 306.000 16.700 306.260 16.960 ;
        RECT 310.140 16.700 310.400 16.960 ;
      LAYER met2 ;
        RECT 1232.430 1700.000 1232.710 1704.000 ;
        RECT 310.140 1688.790 310.400 1689.110 ;
        RECT 310.200 16.990 310.340 1688.790 ;
        RECT 1232.500 1687.750 1232.640 1700.000 ;
        RECT 1232.440 1687.430 1232.700 1687.750 ;
        RECT 306.000 16.670 306.260 16.990 ;
        RECT 310.140 16.670 310.400 16.990 ;
        RECT 306.060 2.400 306.200 16.670 ;
        RECT 305.850 -4.800 306.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 0.300 ;
=======
      LAYER li1 ;
        RECT 1197.065 1686.825 1197.235 1689.375 ;
      LAYER mcon ;
        RECT 1197.065 1689.205 1197.235 1689.375 ;
      LAYER met1 ;
        RECT 323.910 1689.360 324.230 1689.420 ;
        RECT 1197.005 1689.360 1197.295 1689.405 ;
        RECT 323.910 1689.220 1197.295 1689.360 ;
        RECT 323.910 1689.160 324.230 1689.220 ;
        RECT 1197.005 1689.175 1197.295 1689.220 ;
        RECT 1197.005 1686.980 1197.295 1687.025 ;
        RECT 1237.010 1686.980 1237.330 1687.040 ;
        RECT 1197.005 1686.840 1237.330 1686.980 ;
        RECT 1197.005 1686.795 1197.295 1686.840 ;
        RECT 1237.010 1686.780 1237.330 1686.840 ;
      LAYER via ;
        RECT 323.940 1689.160 324.200 1689.420 ;
        RECT 1237.040 1686.780 1237.300 1687.040 ;
      LAYER met2 ;
        RECT 1237.030 1700.000 1237.310 1704.000 ;
        RECT 323.940 1689.130 324.200 1689.450 ;
        RECT 324.000 2.400 324.140 1689.130 ;
        RECT 1237.100 1687.070 1237.240 1700.000 ;
        RECT 1237.040 1686.750 1237.300 1687.070 ;
        RECT 323.790 -4.800 324.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 0.300 ;
=======
      LAYER met1 ;
        RECT 341.390 20.640 341.710 20.700 ;
        RECT 1242.070 20.640 1242.390 20.700 ;
        RECT 341.390 20.500 1242.390 20.640 ;
        RECT 341.390 20.440 341.710 20.500 ;
        RECT 1242.070 20.440 1242.390 20.500 ;
      LAYER via ;
        RECT 341.420 20.440 341.680 20.700 ;
        RECT 1242.100 20.440 1242.360 20.700 ;
      LAYER met2 ;
        RECT 1242.090 1700.000 1242.370 1704.000 ;
        RECT 1242.160 20.730 1242.300 1700.000 ;
        RECT 341.420 20.410 341.680 20.730 ;
        RECT 1242.100 20.410 1242.360 20.730 ;
        RECT 341.480 2.400 341.620 20.410 ;
        RECT 341.270 -4.800 341.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 0.300 ;
=======
      LAYER met1 ;
        RECT 365.310 1689.700 365.630 1689.760 ;
        RECT 1246.670 1689.700 1246.990 1689.760 ;
        RECT 365.310 1689.560 1246.990 1689.700 ;
        RECT 365.310 1689.500 365.630 1689.560 ;
        RECT 1246.670 1689.500 1246.990 1689.560 ;
        RECT 359.330 16.900 359.650 16.960 ;
        RECT 365.310 16.900 365.630 16.960 ;
        RECT 359.330 16.760 365.630 16.900 ;
        RECT 359.330 16.700 359.650 16.760 ;
        RECT 365.310 16.700 365.630 16.760 ;
      LAYER via ;
        RECT 365.340 1689.500 365.600 1689.760 ;
        RECT 1246.700 1689.500 1246.960 1689.760 ;
        RECT 359.360 16.700 359.620 16.960 ;
        RECT 365.340 16.700 365.600 16.960 ;
      LAYER met2 ;
        RECT 1246.690 1700.000 1246.970 1704.000 ;
        RECT 1246.760 1689.790 1246.900 1700.000 ;
        RECT 365.340 1689.470 365.600 1689.790 ;
        RECT 1246.700 1689.470 1246.960 1689.790 ;
        RECT 365.400 16.990 365.540 1689.470 ;
        RECT 359.360 16.670 359.620 16.990 ;
        RECT 365.340 16.670 365.600 16.990 ;
        RECT 359.420 2.400 359.560 16.670 ;
        RECT 359.210 -4.800 359.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 0.300 ;
=======
      LAYER li1 ;
        RECT 414.145 15.725 414.315 16.915 ;
      LAYER mcon ;
        RECT 414.145 16.745 414.315 16.915 ;
      LAYER met1 ;
        RECT 1248.970 1700.920 1249.290 1700.980 ;
        RECT 1250.350 1700.920 1250.670 1700.980 ;
        RECT 1248.970 1700.780 1250.670 1700.920 ;
        RECT 1248.970 1700.720 1249.290 1700.780 ;
        RECT 1250.350 1700.720 1250.670 1700.780 ;
        RECT 1248.970 1435.520 1249.290 1435.780 ;
        RECT 1249.060 1435.100 1249.200 1435.520 ;
        RECT 1248.970 1434.840 1249.290 1435.100 ;
        RECT 414.085 16.900 414.375 16.945 ;
        RECT 1248.970 16.900 1249.290 16.960 ;
        RECT 414.085 16.760 1249.290 16.900 ;
        RECT 414.085 16.715 414.375 16.760 ;
        RECT 1248.970 16.700 1249.290 16.760 ;
        RECT 377.270 15.880 377.590 15.940 ;
        RECT 414.085 15.880 414.375 15.925 ;
        RECT 377.270 15.740 414.375 15.880 ;
        RECT 377.270 15.680 377.590 15.740 ;
        RECT 414.085 15.695 414.375 15.740 ;
      LAYER via ;
        RECT 1249.000 1700.720 1249.260 1700.980 ;
        RECT 1250.380 1700.720 1250.640 1700.980 ;
        RECT 1249.000 1435.520 1249.260 1435.780 ;
        RECT 1249.000 1434.840 1249.260 1435.100 ;
        RECT 1249.000 16.700 1249.260 16.960 ;
        RECT 377.300 15.680 377.560 15.940 ;
      LAYER met2 ;
        RECT 1251.290 1701.090 1251.570 1704.000 ;
        RECT 1250.440 1701.010 1251.570 1701.090 ;
        RECT 1249.000 1700.690 1249.260 1701.010 ;
        RECT 1250.380 1700.950 1251.570 1701.010 ;
        RECT 1250.380 1700.690 1250.640 1700.950 ;
        RECT 1249.060 1435.810 1249.200 1700.690 ;
        RECT 1251.290 1700.000 1251.570 1700.950 ;
        RECT 1249.000 1435.490 1249.260 1435.810 ;
        RECT 1249.000 1434.810 1249.260 1435.130 ;
        RECT 1249.060 16.990 1249.200 1434.810 ;
        RECT 1249.000 16.670 1249.260 16.990 ;
        RECT 377.300 15.650 377.560 15.970 ;
        RECT 377.360 2.400 377.500 15.650 ;
        RECT 377.150 -4.800 377.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 0.300 ;
=======
      LAYER met1 ;
        RECT 399.810 1690.040 400.130 1690.100 ;
        RECT 1256.330 1690.040 1256.650 1690.100 ;
        RECT 399.810 1689.900 1256.650 1690.040 ;
        RECT 399.810 1689.840 400.130 1689.900 ;
        RECT 1256.330 1689.840 1256.650 1689.900 ;
        RECT 395.210 16.900 395.530 16.960 ;
        RECT 399.810 16.900 400.130 16.960 ;
        RECT 395.210 16.760 400.130 16.900 ;
        RECT 395.210 16.700 395.530 16.760 ;
        RECT 399.810 16.700 400.130 16.760 ;
      LAYER via ;
        RECT 399.840 1689.840 400.100 1690.100 ;
        RECT 1256.360 1689.840 1256.620 1690.100 ;
        RECT 395.240 16.700 395.500 16.960 ;
        RECT 399.840 16.700 400.100 16.960 ;
      LAYER met2 ;
        RECT 1256.350 1700.000 1256.630 1704.000 ;
        RECT 1256.420 1690.130 1256.560 1700.000 ;
        RECT 399.840 1689.810 400.100 1690.130 ;
        RECT 1256.360 1689.810 1256.620 1690.130 ;
        RECT 399.900 16.990 400.040 1689.810 ;
        RECT 395.240 16.670 395.500 16.990 ;
        RECT 399.840 16.670 400.100 16.990 ;
        RECT 395.300 2.400 395.440 16.670 ;
        RECT 395.090 -4.800 395.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1257.250 1678.140 1257.570 1678.200 ;
        RECT 1260.010 1678.140 1260.330 1678.200 ;
        RECT 1257.250 1678.000 1260.330 1678.140 ;
        RECT 1257.250 1677.940 1257.570 1678.000 ;
        RECT 1260.010 1677.940 1260.330 1678.000 ;
        RECT 1256.790 16.560 1257.110 16.620 ;
        RECT 448.660 16.420 1257.110 16.560 ;
        RECT 413.150 16.220 413.470 16.280 ;
        RECT 448.660 16.220 448.800 16.420 ;
        RECT 1256.790 16.360 1257.110 16.420 ;
        RECT 413.150 16.080 448.800 16.220 ;
        RECT 413.150 16.020 413.470 16.080 ;
      LAYER via ;
        RECT 1257.280 1677.940 1257.540 1678.200 ;
        RECT 1260.040 1677.940 1260.300 1678.200 ;
        RECT 413.180 16.020 413.440 16.280 ;
        RECT 1256.820 16.360 1257.080 16.620 ;
      LAYER met2 ;
        RECT 1260.950 1700.410 1261.230 1704.000 ;
        RECT 1260.100 1700.270 1261.230 1700.410 ;
        RECT 1260.100 1678.230 1260.240 1700.270 ;
        RECT 1260.950 1700.000 1261.230 1700.270 ;
        RECT 1257.280 1677.910 1257.540 1678.230 ;
        RECT 1260.040 1677.910 1260.300 1678.230 ;
        RECT 1257.340 26.250 1257.480 1677.910 ;
        RECT 1256.880 26.110 1257.480 26.250 ;
        RECT 1256.880 16.650 1257.020 26.110 ;
        RECT 1256.820 16.330 1257.080 16.650 ;
        RECT 413.180 15.990 413.440 16.310 ;
        RECT 413.240 2.400 413.380 15.990 ;
        RECT 413.030 -4.800 413.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 74.010 -4.800 74.570 0.300 ;
=======
        RECT 1169.410 1700.410 1169.690 1704.000 ;
        RECT 1169.020 1700.270 1169.690 1700.410 ;
        RECT 1169.020 18.885 1169.160 1700.270 ;
        RECT 1169.410 1700.000 1169.690 1700.270 ;
        RECT 74.150 18.515 74.430 18.885 ;
        RECT 1168.950 18.515 1169.230 18.885 ;
        RECT 74.220 2.400 74.360 18.515 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 74.150 18.560 74.430 18.840 ;
        RECT 1168.950 18.560 1169.230 18.840 ;
      LAYER met3 ;
        RECT 74.125 18.850 74.455 18.865 ;
        RECT 1168.925 18.850 1169.255 18.865 ;
        RECT 74.125 18.550 1169.255 18.850 ;
        RECT 74.125 18.535 74.455 18.550 ;
        RECT 1168.925 18.535 1169.255 18.550 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 0.300 ;
=======
      LAYER met1 ;
        RECT 434.310 1690.380 434.630 1690.440 ;
        RECT 1265.990 1690.380 1266.310 1690.440 ;
        RECT 434.310 1690.240 1266.310 1690.380 ;
        RECT 434.310 1690.180 434.630 1690.240 ;
        RECT 1265.990 1690.180 1266.310 1690.240 ;
        RECT 430.630 16.560 430.950 16.620 ;
        RECT 434.310 16.560 434.630 16.620 ;
        RECT 430.630 16.420 434.630 16.560 ;
        RECT 430.630 16.360 430.950 16.420 ;
        RECT 434.310 16.360 434.630 16.420 ;
      LAYER via ;
        RECT 434.340 1690.180 434.600 1690.440 ;
        RECT 1266.020 1690.180 1266.280 1690.440 ;
        RECT 430.660 16.360 430.920 16.620 ;
        RECT 434.340 16.360 434.600 16.620 ;
      LAYER met2 ;
        RECT 1266.010 1700.000 1266.290 1704.000 ;
        RECT 1266.080 1690.470 1266.220 1700.000 ;
        RECT 434.340 1690.150 434.600 1690.470 ;
        RECT 1266.020 1690.150 1266.280 1690.470 ;
        RECT 434.400 16.650 434.540 1690.150 ;
        RECT 430.660 16.330 430.920 16.650 ;
        RECT 434.340 16.330 434.600 16.650 ;
        RECT 430.720 2.400 430.860 16.330 ;
        RECT 430.510 -4.800 431.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 0.300 ;
=======
      LAYER met1 ;
        RECT 455.010 1686.640 455.330 1686.700 ;
        RECT 1270.590 1686.640 1270.910 1686.700 ;
        RECT 455.010 1686.500 1270.910 1686.640 ;
        RECT 455.010 1686.440 455.330 1686.500 ;
        RECT 1270.590 1686.440 1270.910 1686.500 ;
        RECT 448.570 15.880 448.890 15.940 ;
        RECT 455.010 15.880 455.330 15.940 ;
        RECT 448.570 15.740 455.330 15.880 ;
        RECT 448.570 15.680 448.890 15.740 ;
        RECT 455.010 15.680 455.330 15.740 ;
      LAYER via ;
        RECT 455.040 1686.440 455.300 1686.700 ;
        RECT 1270.620 1686.440 1270.880 1686.700 ;
        RECT 448.600 15.680 448.860 15.940 ;
        RECT 455.040 15.680 455.300 15.940 ;
      LAYER met2 ;
        RECT 1270.610 1700.000 1270.890 1704.000 ;
        RECT 1270.680 1686.730 1270.820 1700.000 ;
        RECT 455.040 1686.410 455.300 1686.730 ;
        RECT 1270.620 1686.410 1270.880 1686.730 ;
        RECT 455.100 15.970 455.240 1686.410 ;
        RECT 448.600 15.650 448.860 15.970 ;
        RECT 455.040 15.650 455.300 15.970 ;
        RECT 448.660 2.400 448.800 15.650 ;
        RECT 448.450 -4.800 449.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 0.300 ;
=======
      LAYER met1 ;
        RECT 1271.050 1673.040 1271.370 1673.100 ;
        RECT 1274.270 1673.040 1274.590 1673.100 ;
        RECT 1271.050 1672.900 1274.590 1673.040 ;
        RECT 1271.050 1672.840 1271.370 1672.900 ;
        RECT 1274.270 1672.840 1274.590 1672.900 ;
        RECT 466.510 16.220 466.830 16.280 ;
        RECT 1271.050 16.220 1271.370 16.280 ;
        RECT 466.510 16.080 1271.370 16.220 ;
        RECT 466.510 16.020 466.830 16.080 ;
        RECT 1271.050 16.020 1271.370 16.080 ;
      LAYER via ;
        RECT 1271.080 1672.840 1271.340 1673.100 ;
        RECT 1274.300 1672.840 1274.560 1673.100 ;
        RECT 466.540 16.020 466.800 16.280 ;
        RECT 1271.080 16.020 1271.340 16.280 ;
      LAYER met2 ;
        RECT 1275.670 1700.410 1275.950 1704.000 ;
        RECT 1274.360 1700.270 1275.950 1700.410 ;
        RECT 1274.360 1673.130 1274.500 1700.270 ;
        RECT 1275.670 1700.000 1275.950 1700.270 ;
        RECT 1271.080 1672.810 1271.340 1673.130 ;
        RECT 1274.300 1672.810 1274.560 1673.130 ;
        RECT 1271.140 16.310 1271.280 1672.810 ;
        RECT 466.540 15.990 466.800 16.310 ;
        RECT 1271.080 15.990 1271.340 16.310 ;
        RECT 466.600 2.400 466.740 15.990 ;
        RECT 466.390 -4.800 466.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 0.300 ;
=======
      LAYER met1 ;
        RECT 489.510 1686.300 489.830 1686.360 ;
        RECT 1280.250 1686.300 1280.570 1686.360 ;
        RECT 489.510 1686.160 1280.570 1686.300 ;
        RECT 489.510 1686.100 489.830 1686.160 ;
        RECT 1280.250 1686.100 1280.570 1686.160 ;
        RECT 484.450 15.880 484.770 15.940 ;
        RECT 489.510 15.880 489.830 15.940 ;
        RECT 484.450 15.740 489.830 15.880 ;
        RECT 484.450 15.680 484.770 15.740 ;
        RECT 489.510 15.680 489.830 15.740 ;
      LAYER via ;
        RECT 489.540 1686.100 489.800 1686.360 ;
        RECT 1280.280 1686.100 1280.540 1686.360 ;
        RECT 484.480 15.680 484.740 15.940 ;
        RECT 489.540 15.680 489.800 15.940 ;
      LAYER met2 ;
        RECT 1280.270 1700.000 1280.550 1704.000 ;
        RECT 1280.340 1686.390 1280.480 1700.000 ;
        RECT 489.540 1686.070 489.800 1686.390 ;
        RECT 1280.280 1686.070 1280.540 1686.390 ;
        RECT 489.600 15.970 489.740 1686.070 ;
        RECT 484.480 15.650 484.740 15.970 ;
        RECT 489.540 15.650 489.800 15.970 ;
        RECT 484.540 2.400 484.680 15.650 ;
        RECT 484.330 -4.800 484.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 0.300 ;
=======
      LAYER met1 ;
        RECT 1285.310 15.880 1285.630 15.940 ;
        RECT 559.060 15.740 1285.630 15.880 ;
        RECT 502.390 15.540 502.710 15.600 ;
        RECT 559.060 15.540 559.200 15.740 ;
        RECT 1285.310 15.680 1285.630 15.740 ;
        RECT 502.390 15.400 559.200 15.540 ;
        RECT 502.390 15.340 502.710 15.400 ;
      LAYER via ;
        RECT 502.420 15.340 502.680 15.600 ;
        RECT 1285.340 15.680 1285.600 15.940 ;
      LAYER met2 ;
        RECT 1285.330 1700.000 1285.610 1704.000 ;
        RECT 1285.400 15.970 1285.540 1700.000 ;
        RECT 1285.340 15.650 1285.600 15.970 ;
        RECT 502.420 15.310 502.680 15.630 ;
        RECT 502.480 2.400 502.620 15.310 ;
        RECT 502.270 -4.800 502.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 0.300 ;
=======
      LAYER met1 ;
        RECT 524.010 1685.960 524.330 1686.020 ;
        RECT 1289.910 1685.960 1290.230 1686.020 ;
        RECT 524.010 1685.820 1290.230 1685.960 ;
        RECT 524.010 1685.760 524.330 1685.820 ;
        RECT 1289.910 1685.760 1290.230 1685.820 ;
        RECT 519.870 15.880 520.190 15.940 ;
        RECT 524.010 15.880 524.330 15.940 ;
        RECT 519.870 15.740 524.330 15.880 ;
        RECT 519.870 15.680 520.190 15.740 ;
        RECT 524.010 15.680 524.330 15.740 ;
      LAYER via ;
        RECT 524.040 1685.760 524.300 1686.020 ;
        RECT 1289.940 1685.760 1290.200 1686.020 ;
        RECT 519.900 15.680 520.160 15.940 ;
        RECT 524.040 15.680 524.300 15.940 ;
      LAYER met2 ;
        RECT 1289.930 1700.000 1290.210 1704.000 ;
        RECT 1290.000 1686.050 1290.140 1700.000 ;
        RECT 524.040 1685.730 524.300 1686.050 ;
        RECT 1289.940 1685.730 1290.200 1686.050 ;
        RECT 524.100 15.970 524.240 1685.730 ;
        RECT 519.900 15.650 520.160 15.970 ;
        RECT 524.040 15.650 524.300 15.970 ;
        RECT 519.960 2.400 520.100 15.650 ;
        RECT 519.750 -4.800 520.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1290.370 1678.480 1290.690 1678.540 ;
        RECT 1293.590 1678.480 1293.910 1678.540 ;
        RECT 1290.370 1678.340 1293.910 1678.480 ;
        RECT 1290.370 1678.280 1290.690 1678.340 ;
        RECT 1293.590 1678.280 1293.910 1678.340 ;
        RECT 1290.370 15.540 1290.690 15.600 ;
        RECT 600.460 15.400 1290.690 15.540 ;
        RECT 537.810 14.860 538.130 14.920 ;
        RECT 600.460 14.860 600.600 15.400 ;
        RECT 1290.370 15.340 1290.690 15.400 ;
        RECT 537.810 14.720 600.600 14.860 ;
        RECT 537.810 14.660 538.130 14.720 ;
      LAYER via ;
        RECT 1290.400 1678.280 1290.660 1678.540 ;
        RECT 1293.620 1678.280 1293.880 1678.540 ;
        RECT 537.840 14.660 538.100 14.920 ;
        RECT 1290.400 15.340 1290.660 15.600 ;
      LAYER met2 ;
        RECT 1294.990 1700.410 1295.270 1704.000 ;
        RECT 1293.680 1700.270 1295.270 1700.410 ;
        RECT 1293.680 1678.570 1293.820 1700.270 ;
        RECT 1294.990 1700.000 1295.270 1700.270 ;
        RECT 1290.400 1678.250 1290.660 1678.570 ;
        RECT 1293.620 1678.250 1293.880 1678.570 ;
        RECT 1290.460 15.630 1290.600 1678.250 ;
        RECT 1290.400 15.310 1290.660 15.630 ;
        RECT 537.840 14.630 538.100 14.950 ;
        RECT 537.900 2.400 538.040 14.630 ;
        RECT 537.690 -4.800 538.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 0.300 ;
=======
      LAYER met1 ;
        RECT 558.510 1685.620 558.830 1685.680 ;
        RECT 1299.570 1685.620 1299.890 1685.680 ;
        RECT 558.510 1685.480 1299.890 1685.620 ;
        RECT 558.510 1685.420 558.830 1685.480 ;
        RECT 1299.570 1685.420 1299.890 1685.480 ;
        RECT 555.750 15.880 556.070 15.940 ;
        RECT 558.510 15.880 558.830 15.940 ;
        RECT 555.750 15.740 558.830 15.880 ;
        RECT 555.750 15.680 556.070 15.740 ;
        RECT 558.510 15.680 558.830 15.740 ;
      LAYER via ;
        RECT 558.540 1685.420 558.800 1685.680 ;
        RECT 1299.600 1685.420 1299.860 1685.680 ;
        RECT 555.780 15.680 556.040 15.940 ;
        RECT 558.540 15.680 558.800 15.940 ;
      LAYER met2 ;
        RECT 1299.590 1700.000 1299.870 1704.000 ;
        RECT 1299.660 1685.710 1299.800 1700.000 ;
        RECT 558.540 1685.390 558.800 1685.710 ;
        RECT 1299.600 1685.390 1299.860 1685.710 ;
        RECT 558.600 15.970 558.740 1685.390 ;
        RECT 555.780 15.650 556.040 15.970 ;
        RECT 558.540 15.650 558.800 15.970 ;
        RECT 555.840 2.400 555.980 15.650 ;
        RECT 555.630 -4.800 556.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 0.300 ;
=======
      LAYER met1 ;
        RECT 579.210 1685.280 579.530 1685.340 ;
        RECT 1304.630 1685.280 1304.950 1685.340 ;
        RECT 579.210 1685.140 1304.950 1685.280 ;
        RECT 579.210 1685.080 579.530 1685.140 ;
        RECT 1304.630 1685.080 1304.950 1685.140 ;
        RECT 573.690 15.540 574.010 15.600 ;
        RECT 579.210 15.540 579.530 15.600 ;
        RECT 573.690 15.400 579.530 15.540 ;
        RECT 573.690 15.340 574.010 15.400 ;
        RECT 579.210 15.340 579.530 15.400 ;
      LAYER via ;
        RECT 579.240 1685.080 579.500 1685.340 ;
        RECT 1304.660 1685.080 1304.920 1685.340 ;
        RECT 573.720 15.340 573.980 15.600 ;
        RECT 579.240 15.340 579.500 15.600 ;
      LAYER met2 ;
        RECT 1304.650 1700.000 1304.930 1704.000 ;
        RECT 1304.720 1685.370 1304.860 1700.000 ;
        RECT 579.240 1685.050 579.500 1685.370 ;
        RECT 1304.660 1685.050 1304.920 1685.370 ;
        RECT 579.300 15.630 579.440 1685.050 ;
        RECT 573.720 15.310 573.980 15.630 ;
        RECT 579.240 15.310 579.500 15.630 ;
        RECT 573.780 2.400 573.920 15.310 ;
        RECT 573.570 -4.800 574.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1305.090 1675.760 1305.410 1675.820 ;
        RECT 1308.310 1675.760 1308.630 1675.820 ;
        RECT 1305.090 1675.620 1308.630 1675.760 ;
        RECT 1305.090 1675.560 1305.410 1675.620 ;
        RECT 1308.310 1675.560 1308.630 1675.620 ;
        RECT 1304.630 14.860 1304.950 14.920 ;
        RECT 631.740 14.720 1304.950 14.860 ;
        RECT 591.170 14.520 591.490 14.580 ;
        RECT 631.740 14.520 631.880 14.720 ;
        RECT 1304.630 14.660 1304.950 14.720 ;
        RECT 591.170 14.380 631.880 14.520 ;
        RECT 591.170 14.320 591.490 14.380 ;
      LAYER via ;
        RECT 1305.120 1675.560 1305.380 1675.820 ;
        RECT 1308.340 1675.560 1308.600 1675.820 ;
        RECT 591.200 14.320 591.460 14.580 ;
        RECT 1304.660 14.660 1304.920 14.920 ;
      LAYER met2 ;
        RECT 1309.250 1700.410 1309.530 1704.000 ;
        RECT 1308.400 1700.270 1309.530 1700.410 ;
        RECT 1308.400 1675.850 1308.540 1700.270 ;
        RECT 1309.250 1700.000 1309.530 1700.270 ;
        RECT 1305.120 1675.530 1305.380 1675.850 ;
        RECT 1308.340 1675.530 1308.600 1675.850 ;
        RECT 1305.180 20.810 1305.320 1675.530 ;
        RECT 1304.720 20.670 1305.320 20.810 ;
        RECT 1304.720 14.950 1304.860 20.670 ;
        RECT 1304.660 14.630 1304.920 14.950 ;
        RECT 591.200 14.290 591.460 14.610 ;
        RECT 591.260 2.400 591.400 14.290 ;
        RECT 591.050 -4.800 591.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 97.470 -4.800 98.030 0.300 ;
=======
        RECT 1175.850 1700.410 1176.130 1704.000 ;
        RECT 1175.000 1700.270 1176.130 1700.410 ;
        RECT 1175.000 1678.140 1175.140 1700.270 ;
        RECT 1175.850 1700.000 1176.130 1700.270 ;
        RECT 1173.620 1678.000 1175.140 1678.140 ;
        RECT 1173.620 20.245 1173.760 1678.000 ;
        RECT 97.610 19.875 97.890 20.245 ;
        RECT 1173.550 19.875 1173.830 20.245 ;
        RECT 97.680 2.400 97.820 19.875 ;
        RECT 97.470 -4.800 98.030 2.400 ;
      LAYER via2 ;
        RECT 97.610 19.920 97.890 20.200 ;
        RECT 1173.550 19.920 1173.830 20.200 ;
      LAYER met3 ;
        RECT 97.585 20.210 97.915 20.225 ;
        RECT 1173.525 20.210 1173.855 20.225 ;
        RECT 97.585 19.910 1173.855 20.210 ;
        RECT 97.585 19.895 97.915 19.910 ;
        RECT 1173.525 19.895 1173.855 19.910 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 0.300 ;
=======
      LAYER met1 ;
        RECT 955.490 1683.920 955.810 1683.980 ;
        RECT 1314.290 1683.920 1314.610 1683.980 ;
        RECT 955.490 1683.780 1314.610 1683.920 ;
        RECT 955.490 1683.720 955.810 1683.780 ;
        RECT 1314.290 1683.720 1314.610 1683.780 ;
        RECT 609.110 27.440 609.430 27.500 ;
        RECT 955.490 27.440 955.810 27.500 ;
        RECT 609.110 27.300 955.810 27.440 ;
        RECT 609.110 27.240 609.430 27.300 ;
        RECT 955.490 27.240 955.810 27.300 ;
      LAYER via ;
        RECT 955.520 1683.720 955.780 1683.980 ;
        RECT 1314.320 1683.720 1314.580 1683.980 ;
        RECT 609.140 27.240 609.400 27.500 ;
        RECT 955.520 27.240 955.780 27.500 ;
      LAYER met2 ;
        RECT 1314.310 1700.000 1314.590 1704.000 ;
        RECT 1314.380 1684.010 1314.520 1700.000 ;
        RECT 955.520 1683.690 955.780 1684.010 ;
        RECT 1314.320 1683.690 1314.580 1684.010 ;
        RECT 955.580 27.530 955.720 1683.690 ;
        RECT 609.140 27.210 609.400 27.530 ;
        RECT 955.520 27.210 955.780 27.530 ;
        RECT 609.200 2.400 609.340 27.210 ;
        RECT 608.990 -4.800 609.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1317.970 14.520 1318.290 14.580 ;
        RECT 632.200 14.380 1318.290 14.520 ;
        RECT 627.050 14.180 627.370 14.240 ;
        RECT 632.200 14.180 632.340 14.380 ;
        RECT 1317.970 14.320 1318.290 14.380 ;
        RECT 627.050 14.040 632.340 14.180 ;
        RECT 627.050 13.980 627.370 14.040 ;
      LAYER via ;
        RECT 627.080 13.980 627.340 14.240 ;
        RECT 1318.000 14.320 1318.260 14.580 ;
      LAYER met2 ;
        RECT 1318.910 1700.410 1319.190 1704.000 ;
        RECT 1318.060 1700.270 1319.190 1700.410 ;
        RECT 1318.060 14.610 1318.200 1700.270 ;
        RECT 1318.910 1700.000 1319.190 1700.270 ;
        RECT 1318.000 14.290 1318.260 14.610 ;
        RECT 627.080 13.950 627.340 14.270 ;
        RECT 627.140 2.400 627.280 13.950 ;
        RECT 626.930 -4.800 627.490 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 0.300 ;
=======
      LAYER li1 ;
        RECT 227.845 16.405 228.015 17.935 ;
        RECT 275.685 16.405 275.855 17.935 ;
        RECT 276.605 16.065 276.775 17.935 ;
        RECT 323.525 16.065 323.695 17.935 ;
        RECT 373.205 15.045 373.375 17.935 ;
        RECT 420.125 15.045 420.295 17.935 ;
        RECT 469.805 14.705 469.975 17.935 ;
        RECT 516.725 14.705 516.895 17.935 ;
        RECT 566.405 14.365 566.575 17.935 ;
        RECT 613.325 14.025 613.495 17.935 ;
        RECT 663.005 17.765 663.175 21.675 ;
        RECT 709.465 17.935 709.635 21.675 ;
        RECT 709.465 17.765 710.095 17.935 ;
        RECT 856.205 17.765 856.375 21.335 ;
        RECT 903.125 17.765 903.295 21.335 ;
        RECT 952.805 17.765 952.975 21.335 ;
        RECT 999.725 17.765 999.895 21.335 ;
        RECT 1049.405 17.765 1049.575 21.335 ;
        RECT 1096.325 17.765 1096.495 21.335 ;
      LAYER mcon ;
        RECT 663.005 21.505 663.175 21.675 ;
        RECT 227.845 17.765 228.015 17.935 ;
        RECT 275.685 17.765 275.855 17.935 ;
        RECT 276.605 17.765 276.775 17.935 ;
        RECT 323.525 17.765 323.695 17.935 ;
        RECT 373.205 17.765 373.375 17.935 ;
        RECT 420.125 17.765 420.295 17.935 ;
        RECT 469.805 17.765 469.975 17.935 ;
        RECT 516.725 17.765 516.895 17.935 ;
        RECT 566.405 17.765 566.575 17.935 ;
        RECT 613.325 17.765 613.495 17.935 ;
        RECT 709.465 21.505 709.635 21.675 ;
        RECT 856.205 21.165 856.375 21.335 ;
        RECT 709.925 17.765 710.095 17.935 ;
        RECT 903.125 21.165 903.295 21.335 ;
        RECT 952.805 21.165 952.975 21.335 ;
        RECT 999.725 21.165 999.895 21.335 ;
        RECT 1049.405 21.165 1049.575 21.335 ;
        RECT 1096.325 21.165 1096.495 21.335 ;
      LAYER met1 ;
        RECT 662.945 21.660 663.235 21.705 ;
        RECT 709.405 21.660 709.695 21.705 ;
        RECT 662.945 21.520 709.695 21.660 ;
        RECT 662.945 21.475 663.235 21.520 ;
        RECT 709.405 21.475 709.695 21.520 ;
        RECT 856.145 21.320 856.435 21.365 ;
        RECT 903.065 21.320 903.355 21.365 ;
        RECT 856.145 21.180 903.355 21.320 ;
        RECT 856.145 21.135 856.435 21.180 ;
        RECT 903.065 21.135 903.355 21.180 ;
        RECT 952.745 21.320 953.035 21.365 ;
        RECT 999.665 21.320 999.955 21.365 ;
        RECT 952.745 21.180 999.955 21.320 ;
        RECT 952.745 21.135 953.035 21.180 ;
        RECT 999.665 21.135 999.955 21.180 ;
        RECT 1049.345 21.320 1049.635 21.365 ;
        RECT 1096.265 21.320 1096.555 21.365 ;
        RECT 1049.345 21.180 1096.555 21.320 ;
        RECT 1049.345 21.135 1049.635 21.180 ;
        RECT 1096.265 21.135 1096.555 21.180 ;
        RECT 121.510 18.600 121.830 18.660 ;
        RECT 121.510 18.460 139.220 18.600 ;
        RECT 121.510 18.400 121.830 18.460 ;
        RECT 139.080 17.920 139.220 18.460 ;
        RECT 227.785 17.920 228.075 17.965 ;
        RECT 139.080 17.780 228.075 17.920 ;
        RECT 227.785 17.735 228.075 17.780 ;
        RECT 275.625 17.920 275.915 17.965 ;
        RECT 276.545 17.920 276.835 17.965 ;
        RECT 275.625 17.780 276.835 17.920 ;
        RECT 275.625 17.735 275.915 17.780 ;
        RECT 276.545 17.735 276.835 17.780 ;
        RECT 323.465 17.920 323.755 17.965 ;
        RECT 373.145 17.920 373.435 17.965 ;
        RECT 323.465 17.780 373.435 17.920 ;
        RECT 323.465 17.735 323.755 17.780 ;
        RECT 373.145 17.735 373.435 17.780 ;
        RECT 420.065 17.920 420.355 17.965 ;
        RECT 469.745 17.920 470.035 17.965 ;
        RECT 420.065 17.780 470.035 17.920 ;
        RECT 420.065 17.735 420.355 17.780 ;
        RECT 469.745 17.735 470.035 17.780 ;
        RECT 516.665 17.920 516.955 17.965 ;
        RECT 566.345 17.920 566.635 17.965 ;
        RECT 516.665 17.780 566.635 17.920 ;
        RECT 516.665 17.735 516.955 17.780 ;
        RECT 566.345 17.735 566.635 17.780 ;
        RECT 613.265 17.920 613.555 17.965 ;
        RECT 662.945 17.920 663.235 17.965 ;
        RECT 613.265 17.780 663.235 17.920 ;
        RECT 613.265 17.735 613.555 17.780 ;
        RECT 662.945 17.735 663.235 17.780 ;
        RECT 709.865 17.920 710.155 17.965 ;
        RECT 759.530 17.920 759.850 17.980 ;
        RECT 709.865 17.780 759.850 17.920 ;
        RECT 709.865 17.735 710.155 17.780 ;
        RECT 759.530 17.720 759.850 17.780 ;
        RECT 806.450 17.920 806.770 17.980 ;
        RECT 856.145 17.920 856.435 17.965 ;
        RECT 806.450 17.780 856.435 17.920 ;
        RECT 806.450 17.720 806.770 17.780 ;
        RECT 856.145 17.735 856.435 17.780 ;
        RECT 903.065 17.920 903.355 17.965 ;
        RECT 952.745 17.920 953.035 17.965 ;
        RECT 903.065 17.780 953.035 17.920 ;
        RECT 903.065 17.735 903.355 17.780 ;
        RECT 952.745 17.735 953.035 17.780 ;
        RECT 999.665 17.920 999.955 17.965 ;
        RECT 1049.345 17.920 1049.635 17.965 ;
        RECT 999.665 17.780 1049.635 17.920 ;
        RECT 999.665 17.735 999.955 17.780 ;
        RECT 1049.345 17.735 1049.635 17.780 ;
        RECT 1096.265 17.920 1096.555 17.965 ;
        RECT 1180.430 17.920 1180.750 17.980 ;
        RECT 1096.265 17.780 1180.750 17.920 ;
        RECT 1096.265 17.735 1096.555 17.780 ;
        RECT 1180.430 17.720 1180.750 17.780 ;
        RECT 227.785 16.560 228.075 16.605 ;
        RECT 275.625 16.560 275.915 16.605 ;
        RECT 227.785 16.420 275.915 16.560 ;
        RECT 227.785 16.375 228.075 16.420 ;
        RECT 275.625 16.375 275.915 16.420 ;
        RECT 276.545 16.220 276.835 16.265 ;
        RECT 323.465 16.220 323.755 16.265 ;
        RECT 276.545 16.080 323.755 16.220 ;
        RECT 276.545 16.035 276.835 16.080 ;
        RECT 323.465 16.035 323.755 16.080 ;
        RECT 373.145 15.200 373.435 15.245 ;
        RECT 420.065 15.200 420.355 15.245 ;
        RECT 373.145 15.060 420.355 15.200 ;
        RECT 373.145 15.015 373.435 15.060 ;
        RECT 420.065 15.015 420.355 15.060 ;
        RECT 469.745 14.860 470.035 14.905 ;
        RECT 516.665 14.860 516.955 14.905 ;
        RECT 469.745 14.720 516.955 14.860 ;
        RECT 469.745 14.675 470.035 14.720 ;
        RECT 516.665 14.675 516.955 14.720 ;
        RECT 566.345 14.520 566.635 14.565 ;
        RECT 566.345 14.380 590.940 14.520 ;
        RECT 566.345 14.335 566.635 14.380 ;
        RECT 590.800 13.840 590.940 14.380 ;
        RECT 613.265 14.180 613.555 14.225 ;
        RECT 601.380 14.040 613.555 14.180 ;
        RECT 601.380 13.840 601.520 14.040 ;
        RECT 613.265 13.995 613.555 14.040 ;
        RECT 590.800 13.700 601.520 13.840 ;
      LAYER via ;
        RECT 121.540 18.400 121.800 18.660 ;
        RECT 759.560 17.720 759.820 17.980 ;
        RECT 806.480 17.720 806.740 17.980 ;
        RECT 1180.460 17.720 1180.720 17.980 ;
      LAYER met2 ;
        RECT 1182.290 1700.410 1182.570 1704.000 ;
        RECT 1181.440 1700.270 1182.570 1700.410 ;
        RECT 1181.440 1677.290 1181.580 1700.270 ;
        RECT 1182.290 1700.000 1182.570 1700.270 ;
        RECT 1180.520 1677.150 1181.580 1677.290 ;
        RECT 121.540 18.370 121.800 18.690 ;
        RECT 121.600 2.400 121.740 18.370 ;
        RECT 1180.520 18.010 1180.660 1677.150 ;
        RECT 759.560 17.690 759.820 18.010 ;
        RECT 806.480 17.690 806.740 18.010 ;
        RECT 1180.460 17.690 1180.720 18.010 ;
        RECT 759.620 16.165 759.760 17.690 ;
        RECT 806.540 16.165 806.680 17.690 ;
        RECT 759.550 15.795 759.830 16.165 ;
        RECT 806.470 15.795 806.750 16.165 ;
        RECT 121.390 -4.800 121.950 2.400 ;
      LAYER via2 ;
        RECT 759.550 15.840 759.830 16.120 ;
        RECT 806.470 15.840 806.750 16.120 ;
      LAYER met3 ;
        RECT 759.525 16.130 759.855 16.145 ;
        RECT 806.445 16.130 806.775 16.145 ;
        RECT 759.525 15.830 806.775 16.130 ;
        RECT 759.525 15.815 759.855 15.830 ;
        RECT 806.445 15.815 806.775 15.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 0.300 ;
=======
      LAYER li1 ;
        RECT 276.605 18.445 276.775 20.655 ;
        RECT 323.525 18.445 323.695 20.655 ;
        RECT 373.205 18.445 373.835 18.615 ;
        RECT 373.665 16.405 373.835 18.445 ;
        RECT 419.665 18.445 420.295 18.615 ;
        RECT 469.805 18.445 470.435 18.615 ;
        RECT 419.665 16.405 419.835 18.445 ;
        RECT 470.265 14.365 470.435 18.445 ;
        RECT 516.265 18.445 516.895 18.615 ;
        RECT 566.405 18.445 566.575 20.995 ;
        RECT 613.325 18.445 613.495 20.995 ;
        RECT 759.605 18.445 759.775 21.675 ;
        RECT 806.525 18.445 806.695 21.675 ;
        RECT 1049.865 18.445 1050.035 21.675 ;
        RECT 516.265 14.365 516.435 18.445 ;
      LAYER mcon ;
        RECT 759.605 21.505 759.775 21.675 ;
        RECT 566.405 20.825 566.575 20.995 ;
        RECT 276.605 20.485 276.775 20.655 ;
        RECT 323.525 20.485 323.695 20.655 ;
        RECT 420.125 18.445 420.295 18.615 ;
        RECT 516.725 18.445 516.895 18.615 ;
        RECT 613.325 20.825 613.495 20.995 ;
        RECT 806.525 21.505 806.695 21.675 ;
        RECT 1049.865 21.505 1050.035 21.675 ;
      LAYER met1 ;
        RECT 759.545 21.660 759.835 21.705 ;
        RECT 806.465 21.660 806.755 21.705 ;
        RECT 759.545 21.520 806.755 21.660 ;
        RECT 759.545 21.475 759.835 21.520 ;
        RECT 806.465 21.475 806.755 21.520 ;
        RECT 1049.805 21.660 1050.095 21.705 ;
        RECT 1095.790 21.660 1096.110 21.720 ;
        RECT 1049.805 21.520 1096.110 21.660 ;
        RECT 1049.805 21.475 1050.095 21.520 ;
        RECT 1095.790 21.460 1096.110 21.520 ;
        RECT 566.345 20.980 566.635 21.025 ;
        RECT 613.265 20.980 613.555 21.025 ;
        RECT 566.345 20.840 613.555 20.980 ;
        RECT 566.345 20.795 566.635 20.840 ;
        RECT 613.265 20.795 613.555 20.840 ;
        RECT 276.545 20.640 276.835 20.685 ;
        RECT 323.465 20.640 323.755 20.685 ;
        RECT 276.545 20.500 323.755 20.640 ;
        RECT 276.545 20.455 276.835 20.500 ;
        RECT 323.465 20.455 323.755 20.500 ;
        RECT 145.430 18.600 145.750 18.660 ;
        RECT 276.545 18.600 276.835 18.645 ;
        RECT 145.430 18.460 276.835 18.600 ;
        RECT 145.430 18.400 145.750 18.460 ;
        RECT 276.545 18.415 276.835 18.460 ;
        RECT 323.465 18.600 323.755 18.645 ;
        RECT 373.145 18.600 373.435 18.645 ;
        RECT 323.465 18.460 373.435 18.600 ;
        RECT 323.465 18.415 323.755 18.460 ;
        RECT 373.145 18.415 373.435 18.460 ;
        RECT 420.065 18.600 420.355 18.645 ;
        RECT 469.745 18.600 470.035 18.645 ;
        RECT 420.065 18.460 470.035 18.600 ;
        RECT 420.065 18.415 420.355 18.460 ;
        RECT 469.745 18.415 470.035 18.460 ;
        RECT 516.665 18.600 516.955 18.645 ;
        RECT 566.345 18.600 566.635 18.645 ;
        RECT 516.665 18.460 566.635 18.600 ;
        RECT 516.665 18.415 516.955 18.460 ;
        RECT 566.345 18.415 566.635 18.460 ;
        RECT 613.265 18.600 613.555 18.645 ;
        RECT 663.390 18.600 663.710 18.660 ;
        RECT 613.265 18.460 663.710 18.600 ;
        RECT 613.265 18.415 613.555 18.460 ;
        RECT 663.390 18.400 663.710 18.460 ;
        RECT 709.390 18.600 709.710 18.660 ;
        RECT 759.545 18.600 759.835 18.645 ;
        RECT 709.390 18.460 759.835 18.600 ;
        RECT 709.390 18.400 709.710 18.460 ;
        RECT 759.545 18.415 759.835 18.460 ;
        RECT 806.465 18.600 806.755 18.645 ;
        RECT 856.130 18.600 856.450 18.660 ;
        RECT 806.465 18.460 856.450 18.600 ;
        RECT 806.465 18.415 806.755 18.460 ;
        RECT 856.130 18.400 856.450 18.460 ;
        RECT 903.050 18.600 903.370 18.660 ;
        RECT 952.730 18.600 953.050 18.660 ;
        RECT 903.050 18.460 953.050 18.600 ;
        RECT 903.050 18.400 903.370 18.460 ;
        RECT 952.730 18.400 953.050 18.460 ;
        RECT 999.650 18.600 999.970 18.660 ;
        RECT 1049.805 18.600 1050.095 18.645 ;
        RECT 999.650 18.460 1050.095 18.600 ;
        RECT 999.650 18.400 999.970 18.460 ;
        RECT 1049.805 18.415 1050.095 18.460 ;
        RECT 1096.250 18.600 1096.570 18.660 ;
        RECT 1188.710 18.600 1189.030 18.660 ;
        RECT 1096.250 18.460 1189.030 18.600 ;
        RECT 1096.250 18.400 1096.570 18.460 ;
        RECT 1188.710 18.400 1189.030 18.460 ;
        RECT 373.605 16.560 373.895 16.605 ;
        RECT 419.605 16.560 419.895 16.605 ;
        RECT 373.605 16.420 419.895 16.560 ;
        RECT 373.605 16.375 373.895 16.420 ;
        RECT 419.605 16.375 419.895 16.420 ;
        RECT 470.205 14.520 470.495 14.565 ;
        RECT 516.205 14.520 516.495 14.565 ;
        RECT 470.205 14.380 516.495 14.520 ;
        RECT 470.205 14.335 470.495 14.380 ;
        RECT 516.205 14.335 516.495 14.380 ;
      LAYER via ;
        RECT 1095.820 21.460 1096.080 21.720 ;
        RECT 145.460 18.400 145.720 18.660 ;
        RECT 663.420 18.400 663.680 18.660 ;
        RECT 709.420 18.400 709.680 18.660 ;
        RECT 856.160 18.400 856.420 18.660 ;
        RECT 903.080 18.400 903.340 18.660 ;
        RECT 952.760 18.400 953.020 18.660 ;
        RECT 999.680 18.400 999.940 18.660 ;
        RECT 1096.280 18.400 1096.540 18.660 ;
        RECT 1188.740 18.400 1189.000 18.660 ;
      LAYER met2 ;
        RECT 1188.730 1700.000 1189.010 1704.000 ;
        RECT 1095.820 21.490 1096.080 21.750 ;
        RECT 1095.820 21.430 1096.480 21.490 ;
        RECT 1095.880 21.350 1096.480 21.430 ;
        RECT 663.410 20.555 663.690 20.925 ;
        RECT 709.410 20.555 709.690 20.925 ;
        RECT 856.150 20.555 856.430 20.925 ;
        RECT 903.070 20.555 903.350 20.925 ;
        RECT 952.750 20.555 953.030 20.925 ;
        RECT 999.670 20.555 999.950 20.925 ;
        RECT 663.480 18.690 663.620 20.555 ;
        RECT 709.480 18.690 709.620 20.555 ;
        RECT 856.220 18.690 856.360 20.555 ;
        RECT 903.140 18.690 903.280 20.555 ;
        RECT 952.820 18.690 952.960 20.555 ;
        RECT 999.740 18.690 999.880 20.555 ;
        RECT 1096.340 18.690 1096.480 21.350 ;
        RECT 1188.800 18.690 1188.940 1700.000 ;
        RECT 145.460 18.370 145.720 18.690 ;
        RECT 663.420 18.370 663.680 18.690 ;
        RECT 709.420 18.370 709.680 18.690 ;
        RECT 856.160 18.370 856.420 18.690 ;
        RECT 903.080 18.370 903.340 18.690 ;
        RECT 952.760 18.370 953.020 18.690 ;
        RECT 999.680 18.370 999.940 18.690 ;
        RECT 1096.280 18.370 1096.540 18.690 ;
        RECT 1188.740 18.370 1189.000 18.690 ;
        RECT 145.520 2.400 145.660 18.370 ;
        RECT 145.310 -4.800 145.870 2.400 ;
      LAYER via2 ;
        RECT 663.410 20.600 663.690 20.880 ;
        RECT 709.410 20.600 709.690 20.880 ;
        RECT 856.150 20.600 856.430 20.880 ;
        RECT 903.070 20.600 903.350 20.880 ;
        RECT 952.750 20.600 953.030 20.880 ;
        RECT 999.670 20.600 999.950 20.880 ;
      LAYER met3 ;
        RECT 663.385 20.890 663.715 20.905 ;
        RECT 709.385 20.890 709.715 20.905 ;
        RECT 663.385 20.590 709.715 20.890 ;
        RECT 663.385 20.575 663.715 20.590 ;
        RECT 709.385 20.575 709.715 20.590 ;
        RECT 856.125 20.890 856.455 20.905 ;
        RECT 903.045 20.890 903.375 20.905 ;
        RECT 856.125 20.590 903.375 20.890 ;
        RECT 856.125 20.575 856.455 20.590 ;
        RECT 903.045 20.575 903.375 20.590 ;
        RECT 952.725 20.890 953.055 20.905 ;
        RECT 999.645 20.890 999.975 20.905 ;
        RECT 952.725 20.590 999.975 20.890 ;
        RECT 952.725 20.575 953.055 20.590 ;
        RECT 999.645 20.575 999.975 20.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 0.300 ;
=======
      LAYER met1 ;
        RECT 163.370 14.180 163.690 14.240 ;
        RECT 165.210 14.180 165.530 14.240 ;
        RECT 163.370 14.040 165.530 14.180 ;
        RECT 163.370 13.980 163.690 14.040 ;
        RECT 165.210 13.980 165.530 14.040 ;
      LAYER via ;
        RECT 163.400 13.980 163.660 14.240 ;
        RECT 165.240 13.980 165.500 14.240 ;
      LAYER met2 ;
        RECT 1193.790 1700.000 1194.070 1704.000 ;
        RECT 1193.860 1689.645 1194.000 1700.000 ;
        RECT 165.230 1689.275 165.510 1689.645 ;
        RECT 1193.790 1689.275 1194.070 1689.645 ;
        RECT 165.300 14.270 165.440 1689.275 ;
        RECT 163.400 13.950 163.660 14.270 ;
        RECT 165.240 13.950 165.500 14.270 ;
        RECT 163.460 2.400 163.600 13.950 ;
        RECT 163.250 -4.800 163.810 2.400 ;
      LAYER via2 ;
        RECT 165.230 1689.320 165.510 1689.600 ;
        RECT 1193.790 1689.320 1194.070 1689.600 ;
      LAYER met3 ;
        RECT 165.205 1689.610 165.535 1689.625 ;
        RECT 1193.765 1689.610 1194.095 1689.625 ;
        RECT 165.205 1689.310 1194.095 1689.610 ;
        RECT 165.205 1689.295 165.535 1689.310 ;
        RECT 1193.765 1689.295 1194.095 1689.310 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 0.300 ;
=======
      LAYER li1 ;
        RECT 1149.225 17.425 1149.395 19.295 ;
      LAYER mcon ;
        RECT 1149.225 19.125 1149.395 19.295 ;
      LAYER met1 ;
        RECT 180.850 19.280 181.170 19.340 ;
        RECT 1149.165 19.280 1149.455 19.325 ;
        RECT 180.850 19.140 1149.455 19.280 ;
        RECT 180.850 19.080 181.170 19.140 ;
        RECT 1149.165 19.095 1149.455 19.140 ;
        RECT 1149.165 17.580 1149.455 17.625 ;
        RECT 1195.610 17.580 1195.930 17.640 ;
        RECT 1149.165 17.440 1195.930 17.580 ;
        RECT 1149.165 17.395 1149.455 17.440 ;
        RECT 1195.610 17.380 1195.930 17.440 ;
      LAYER via ;
        RECT 180.880 19.080 181.140 19.340 ;
        RECT 1195.640 17.380 1195.900 17.640 ;
      LAYER met2 ;
        RECT 1198.390 1700.410 1198.670 1704.000 ;
        RECT 1197.540 1700.270 1198.670 1700.410 ;
        RECT 1197.540 1678.140 1197.680 1700.270 ;
        RECT 1198.390 1700.000 1198.670 1700.270 ;
        RECT 1195.700 1678.000 1197.680 1678.140 ;
        RECT 180.880 19.050 181.140 19.370 ;
        RECT 180.940 2.400 181.080 19.050 ;
        RECT 1195.700 17.670 1195.840 1678.000 ;
        RECT 1195.640 17.350 1195.900 17.670 ;
        RECT 180.730 -4.800 181.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 0.300 ;
=======
      LAYER met1 ;
        RECT 1203.430 1688.000 1203.750 1688.060 ;
        RECT 1178.220 1687.860 1203.750 1688.000 ;
        RECT 199.710 1687.660 200.030 1687.720 ;
        RECT 1178.220 1687.660 1178.360 1687.860 ;
        RECT 1203.430 1687.800 1203.750 1687.860 ;
        RECT 199.710 1687.520 1178.360 1687.660 ;
        RECT 199.710 1687.460 200.030 1687.520 ;
      LAYER via ;
        RECT 199.740 1687.460 200.000 1687.720 ;
        RECT 1203.460 1687.800 1203.720 1688.060 ;
      LAYER met2 ;
        RECT 1203.450 1700.000 1203.730 1704.000 ;
        RECT 1203.520 1688.090 1203.660 1700.000 ;
        RECT 1203.460 1687.770 1203.720 1688.090 ;
        RECT 199.740 1687.430 200.000 1687.750 ;
        RECT 199.800 14.690 199.940 1687.430 ;
        RECT 199.340 14.550 199.940 14.690 ;
        RECT 199.340 14.010 199.480 14.550 ;
        RECT 198.880 13.870 199.480 14.010 ;
        RECT 198.880 2.400 199.020 13.870 ;
        RECT 198.670 -4.800 199.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 0.300 ;
=======
      LAYER met1 ;
        RECT 216.730 19.960 217.050 20.020 ;
        RECT 1208.490 19.960 1208.810 20.020 ;
        RECT 216.730 19.820 1208.810 19.960 ;
        RECT 216.730 19.760 217.050 19.820 ;
        RECT 1208.490 19.760 1208.810 19.820 ;
      LAYER via ;
        RECT 216.760 19.760 217.020 20.020 ;
        RECT 1208.520 19.760 1208.780 20.020 ;
      LAYER met2 ;
        RECT 1208.050 1700.410 1208.330 1704.000 ;
        RECT 1208.050 1700.270 1208.720 1700.410 ;
        RECT 1208.050 1700.000 1208.330 1700.270 ;
        RECT 1208.580 20.050 1208.720 1700.270 ;
        RECT 216.760 19.730 217.020 20.050 ;
        RECT 1208.520 19.730 1208.780 20.050 ;
        RECT 216.820 2.400 216.960 19.730 ;
        RECT 216.610 -4.800 217.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1213.090 1688.340 1213.410 1688.400 ;
        RECT 1177.760 1688.200 1213.410 1688.340 ;
        RECT 241.110 1688.000 241.430 1688.060 ;
        RECT 1177.760 1688.000 1177.900 1688.200 ;
        RECT 1213.090 1688.140 1213.410 1688.200 ;
        RECT 241.110 1687.860 1177.900 1688.000 ;
        RECT 241.110 1687.800 241.430 1687.860 ;
        RECT 234.670 16.900 234.990 16.960 ;
        RECT 241.110 16.900 241.430 16.960 ;
        RECT 234.670 16.760 241.430 16.900 ;
        RECT 234.670 16.700 234.990 16.760 ;
        RECT 241.110 16.700 241.430 16.760 ;
      LAYER via ;
        RECT 241.140 1687.800 241.400 1688.060 ;
        RECT 1213.120 1688.140 1213.380 1688.400 ;
        RECT 234.700 16.700 234.960 16.960 ;
        RECT 241.140 16.700 241.400 16.960 ;
      LAYER met2 ;
        RECT 1213.110 1700.000 1213.390 1704.000 ;
        RECT 1213.180 1688.430 1213.320 1700.000 ;
        RECT 1213.120 1688.110 1213.380 1688.430 ;
        RECT 241.140 1687.770 241.400 1688.090 ;
        RECT 241.200 16.990 241.340 1687.770 ;
        RECT 234.700 16.670 234.960 16.990 ;
        RECT 241.140 16.670 241.400 16.990 ;
        RECT 234.760 2.400 234.900 16.670 ;
        RECT 234.550 -4.800 235.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 0.300 ;
=======
      LAYER met1 ;
        RECT 1159.270 1690.720 1159.590 1690.780 ;
        RECT 1163.410 1690.720 1163.730 1690.780 ;
        RECT 1159.270 1690.580 1163.730 1690.720 ;
        RECT 1159.270 1690.520 1159.590 1690.580 ;
        RECT 1163.410 1690.520 1163.730 1690.580 ;
      LAYER via ;
        RECT 1159.300 1690.520 1159.560 1690.780 ;
        RECT 1163.440 1690.520 1163.700 1690.780 ;
      LAYER met2 ;
        RECT 1164.810 1700.410 1165.090 1704.000 ;
        RECT 1163.500 1700.270 1165.090 1700.410 ;
        RECT 1163.500 1690.810 1163.640 1700.270 ;
        RECT 1164.810 1700.000 1165.090 1700.270 ;
        RECT 1159.300 1690.490 1159.560 1690.810 ;
        RECT 1163.440 1690.490 1163.700 1690.810 ;
        RECT 1159.360 18.205 1159.500 1690.490 ;
        RECT 56.210 17.835 56.490 18.205 ;
        RECT 1159.290 17.835 1159.570 18.205 ;
        RECT 56.280 2.400 56.420 17.835 ;
        RECT 56.070 -4.800 56.630 2.400 ;
      LAYER via2 ;
        RECT 56.210 17.880 56.490 18.160 ;
        RECT 1159.290 17.880 1159.570 18.160 ;
      LAYER met3 ;
        RECT 56.185 18.170 56.515 18.185 ;
        RECT 1159.265 18.170 1159.595 18.185 ;
        RECT 56.185 17.870 1159.595 18.170 ;
        RECT 56.185 17.855 56.515 17.870 ;
        RECT 1159.265 17.855 1159.595 17.870 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 0.300 ;
=======
      LAYER met1 ;
        RECT 80.110 17.580 80.430 17.640 ;
        RECT 82.410 17.580 82.730 17.640 ;
        RECT 80.110 17.440 82.730 17.580 ;
        RECT 80.110 17.380 80.430 17.440 ;
        RECT 82.410 17.380 82.730 17.440 ;
      LAYER via ;
        RECT 80.140 17.380 80.400 17.640 ;
        RECT 82.440 17.380 82.700 17.640 ;
      LAYER met2 ;
        RECT 1171.250 1700.000 1171.530 1704.000 ;
        RECT 1171.320 1687.605 1171.460 1700.000 ;
        RECT 82.430 1687.235 82.710 1687.605 ;
        RECT 1171.250 1687.235 1171.530 1687.605 ;
        RECT 82.500 17.670 82.640 1687.235 ;
        RECT 80.140 17.350 80.400 17.670 ;
        RECT 82.440 17.350 82.700 17.670 ;
        RECT 80.200 2.400 80.340 17.350 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 82.430 1687.280 82.710 1687.560 ;
        RECT 1171.250 1687.280 1171.530 1687.560 ;
      LAYER met3 ;
        RECT 82.405 1687.570 82.735 1687.585 ;
        RECT 1171.225 1687.570 1171.555 1687.585 ;
        RECT 82.405 1687.270 1171.555 1687.570 ;
        RECT 82.405 1687.255 82.735 1687.270 ;
        RECT 1171.225 1687.255 1171.555 1687.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 0.300 ;
=======
      LAYER li1 ;
        RECT 1149.685 17.255 1149.855 19.295 ;
        RECT 1148.305 17.085 1149.855 17.255 ;
      LAYER mcon ;
        RECT 1149.685 19.125 1149.855 19.295 ;
      LAYER met1 ;
        RECT 1149.625 19.280 1149.915 19.325 ;
        RECT 1173.990 19.280 1174.310 19.340 ;
        RECT 1149.625 19.140 1174.310 19.280 ;
        RECT 1149.625 19.095 1149.915 19.140 ;
        RECT 1173.990 19.080 1174.310 19.140 ;
        RECT 103.570 17.240 103.890 17.300 ;
        RECT 1148.245 17.240 1148.535 17.285 ;
        RECT 103.570 17.100 1148.535 17.240 ;
        RECT 103.570 17.040 103.890 17.100 ;
        RECT 1148.245 17.055 1148.535 17.100 ;
      LAYER via ;
        RECT 1174.020 19.080 1174.280 19.340 ;
        RECT 103.600 17.040 103.860 17.300 ;
      LAYER met2 ;
        RECT 1177.690 1700.410 1177.970 1704.000 ;
        RECT 1176.380 1700.270 1177.970 1700.410 ;
        RECT 1176.380 1677.290 1176.520 1700.270 ;
        RECT 1177.690 1700.000 1177.970 1700.270 ;
        RECT 1174.080 1677.150 1176.520 1677.290 ;
        RECT 1174.080 19.370 1174.220 1677.150 ;
        RECT 1174.020 19.050 1174.280 19.370 ;
        RECT 103.600 17.010 103.860 17.330 ;
        RECT 103.660 2.400 103.800 17.010 ;
        RECT 103.450 -4.800 104.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 0.300 ;
=======
      LAYER met1 ;
        RECT 127.490 16.900 127.810 16.960 ;
        RECT 130.710 16.900 131.030 16.960 ;
        RECT 127.490 16.760 131.030 16.900 ;
        RECT 127.490 16.700 127.810 16.760 ;
        RECT 130.710 16.700 131.030 16.760 ;
      LAYER via ;
        RECT 127.520 16.700 127.780 16.960 ;
        RECT 130.740 16.700 131.000 16.960 ;
      LAYER met2 ;
        RECT 1184.130 1700.000 1184.410 1704.000 ;
        RECT 1184.200 1688.285 1184.340 1700.000 ;
        RECT 130.730 1687.915 131.010 1688.285 ;
        RECT 1184.130 1687.915 1184.410 1688.285 ;
        RECT 130.800 16.990 130.940 1687.915 ;
        RECT 127.520 16.670 127.780 16.990 ;
        RECT 130.740 16.670 131.000 16.990 ;
        RECT 127.580 2.400 127.720 16.670 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 130.730 1687.960 131.010 1688.240 ;
        RECT 1184.130 1687.960 1184.410 1688.240 ;
      LAYER met3 ;
        RECT 130.705 1688.250 131.035 1688.265 ;
        RECT 1184.105 1688.250 1184.435 1688.265 ;
        RECT 130.705 1687.950 1184.435 1688.250 ;
        RECT 130.705 1687.935 131.035 1687.950 ;
        RECT 1184.105 1687.935 1184.435 1687.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1153.750 1690.720 1154.070 1690.780 ;
        RECT 1155.590 1690.720 1155.910 1690.780 ;
        RECT 1153.750 1690.580 1155.910 1690.720 ;
        RECT 1153.750 1690.520 1154.070 1690.580 ;
        RECT 1155.590 1690.520 1155.910 1690.580 ;
      LAYER via ;
        RECT 1153.780 1690.520 1154.040 1690.780 ;
        RECT 1155.620 1690.520 1155.880 1690.780 ;
      LAYER met2 ;
        RECT 1156.530 1700.410 1156.810 1704.000 ;
        RECT 1155.680 1700.270 1156.810 1700.410 ;
        RECT 1155.680 1690.810 1155.820 1700.270 ;
        RECT 1156.530 1700.000 1156.810 1700.270 ;
        RECT 1153.780 1690.490 1154.040 1690.810 ;
        RECT 1155.620 1690.490 1155.880 1690.810 ;
        RECT 1153.840 16.845 1153.980 1690.490 ;
        RECT 26.310 16.475 26.590 16.845 ;
        RECT 1153.770 16.475 1154.050 16.845 ;
        RECT 26.380 2.400 26.520 16.475 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 26.310 16.520 26.590 16.800 ;
        RECT 1153.770 16.520 1154.050 16.800 ;
      LAYER met3 ;
        RECT 26.285 16.810 26.615 16.825 ;
        RECT 1153.745 16.810 1154.075 16.825 ;
        RECT 26.285 16.510 1154.075 16.810 ;
        RECT 26.285 16.495 26.615 16.510 ;
        RECT 1153.745 16.495 1154.075 16.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 32.150 -4.800 32.710 0.300 ;
=======
        RECT 1158.370 1700.000 1158.650 1704.000 ;
        RECT 1158.440 1686.925 1158.580 1700.000 ;
        RECT 34.130 1686.555 34.410 1686.925 ;
        RECT 1158.370 1686.555 1158.650 1686.925 ;
        RECT 34.200 3.130 34.340 1686.555 ;
        RECT 32.360 2.990 34.340 3.130 ;
        RECT 32.360 2.400 32.500 2.990 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 34.130 1686.600 34.410 1686.880 ;
        RECT 1158.370 1686.600 1158.650 1686.880 ;
      LAYER met3 ;
        RECT 34.105 1686.890 34.435 1686.905 ;
        RECT 1158.345 1686.890 1158.675 1686.905 ;
        RECT 34.105 1686.590 1158.675 1686.890 ;
        RECT 34.105 1686.575 34.435 1686.590 ;
        RECT 1158.345 1686.575 1158.675 1686.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
<<<<<<< HEAD
        RECT 4.020 3519.700 7.020 3529.000 ;
        RECT 184.020 3519.700 187.020 3529.000 ;
        RECT 364.020 3519.700 367.020 3529.000 ;
        RECT 544.020 3519.700 547.020 3529.000 ;
        RECT 724.020 3519.700 727.020 3529.000 ;
        RECT 904.020 3519.700 907.020 3529.000 ;
        RECT 1084.020 3519.700 1087.020 3529.000 ;
        RECT 1264.020 3519.700 1267.020 3529.000 ;
        RECT 1444.020 3519.700 1447.020 3529.000 ;
        RECT 1624.020 3519.700 1627.020 3529.000 ;
        RECT 1804.020 3519.700 1807.020 3529.000 ;
        RECT 1984.020 3519.700 1987.020 3529.000 ;
        RECT 2164.020 3519.700 2167.020 3529.000 ;
        RECT 2344.020 3519.700 2347.020 3529.000 ;
        RECT 2524.020 3519.700 2527.020 3529.000 ;
        RECT 2704.020 3519.700 2707.020 3529.000 ;
        RECT 2884.020 3519.700 2887.020 3529.000 ;
        RECT 4.020 -9.320 7.020 0.300 ;
        RECT 184.020 -9.320 187.020 0.300 ;
        RECT 364.020 -9.320 367.020 0.300 ;
        RECT 544.020 -9.320 547.020 0.300 ;
        RECT 724.020 -9.320 727.020 0.300 ;
        RECT 904.020 -9.320 907.020 0.300 ;
        RECT 1084.020 -9.320 1087.020 0.300 ;
        RECT 1264.020 -9.320 1267.020 0.300 ;
        RECT 1444.020 -9.320 1447.020 0.300 ;
        RECT 1624.020 -9.320 1627.020 0.300 ;
        RECT 1804.020 -9.320 1807.020 0.300 ;
        RECT 1984.020 -9.320 1987.020 0.300 ;
        RECT 2164.020 -9.320 2167.020 0.300 ;
        RECT 2344.020 -9.320 2347.020 0.300 ;
        RECT 2524.020 -9.320 2527.020 0.300 ;
        RECT 2704.020 -9.320 2707.020 0.300 ;
        RECT 2884.020 -9.320 2887.020 0.300 ;
=======
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 -9.220 547.020 3528.900 ;
        RECT 724.020 -9.220 727.020 3528.900 ;
        RECT 904.020 -9.220 907.020 3528.900 ;
        RECT 1084.020 -9.220 1087.020 3528.900 ;
        RECT 1264.020 -9.220 1267.020 3528.900 ;
        RECT 1444.020 -9.220 1447.020 3528.900 ;
        RECT 1624.020 -9.220 1627.020 3528.900 ;
        RECT 1804.020 -9.220 1807.020 3528.900 ;
        RECT 1984.020 -9.220 1987.020 3528.900 ;
        RECT 2164.020 -9.220 2167.020 3528.900 ;
        RECT 2344.020 -9.220 2347.020 3528.900 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
>>>>>>> Latest run - not LVS matched yet
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
<<<<<<< HEAD
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT -9.070 3430.850 -7.890 3432.030 ;
        RECT -9.070 3429.250 -7.890 3430.430 ;
        RECT -9.070 3250.850 -7.890 3252.030 ;
        RECT -9.070 3249.250 -7.890 3250.430 ;
        RECT -9.070 3070.850 -7.890 3072.030 ;
        RECT -9.070 3069.250 -7.890 3070.430 ;
        RECT -9.070 2890.850 -7.890 2892.030 ;
        RECT -9.070 2889.250 -7.890 2890.430 ;
        RECT -9.070 2710.850 -7.890 2712.030 ;
        RECT -9.070 2709.250 -7.890 2710.430 ;
        RECT -9.070 2530.850 -7.890 2532.030 ;
        RECT -9.070 2529.250 -7.890 2530.430 ;
        RECT -9.070 2350.850 -7.890 2352.030 ;
        RECT -9.070 2349.250 -7.890 2350.430 ;
        RECT -9.070 2170.850 -7.890 2172.030 ;
        RECT -9.070 2169.250 -7.890 2170.430 ;
        RECT -9.070 1990.850 -7.890 1992.030 ;
        RECT -9.070 1989.250 -7.890 1990.430 ;
        RECT -9.070 1810.850 -7.890 1812.030 ;
        RECT -9.070 1809.250 -7.890 1810.430 ;
        RECT -9.070 1630.850 -7.890 1632.030 ;
        RECT -9.070 1629.250 -7.890 1630.430 ;
        RECT -9.070 1450.850 -7.890 1452.030 ;
        RECT -9.070 1449.250 -7.890 1450.430 ;
        RECT -9.070 1270.850 -7.890 1272.030 ;
        RECT -9.070 1269.250 -7.890 1270.430 ;
        RECT -9.070 1090.850 -7.890 1092.030 ;
        RECT -9.070 1089.250 -7.890 1090.430 ;
        RECT -9.070 910.850 -7.890 912.030 ;
        RECT -9.070 909.250 -7.890 910.430 ;
        RECT -9.070 730.850 -7.890 732.030 ;
        RECT -9.070 729.250 -7.890 730.430 ;
        RECT -9.070 550.850 -7.890 552.030 ;
        RECT -9.070 549.250 -7.890 550.430 ;
        RECT -9.070 370.850 -7.890 372.030 ;
        RECT -9.070 369.250 -7.890 370.430 ;
        RECT -9.070 190.850 -7.890 192.030 ;
        RECT -9.070 189.250 -7.890 190.430 ;
        RECT -9.070 10.850 -7.890 12.030 ;
        RECT -9.070 9.250 -7.890 10.430 ;
        RECT 2927.510 3430.850 2928.690 3432.030 ;
        RECT 2927.510 3429.250 2928.690 3430.430 ;
        RECT 2927.510 3250.850 2928.690 3252.030 ;
        RECT 2927.510 3249.250 2928.690 3250.430 ;
        RECT 2927.510 3070.850 2928.690 3072.030 ;
        RECT 2927.510 3069.250 2928.690 3070.430 ;
        RECT 2927.510 2890.850 2928.690 2892.030 ;
        RECT 2927.510 2889.250 2928.690 2890.430 ;
        RECT 2927.510 2710.850 2928.690 2712.030 ;
        RECT 2927.510 2709.250 2928.690 2710.430 ;
        RECT 2927.510 2530.850 2928.690 2532.030 ;
        RECT 2927.510 2529.250 2928.690 2530.430 ;
        RECT 2927.510 2350.850 2928.690 2352.030 ;
        RECT 2927.510 2349.250 2928.690 2350.430 ;
        RECT 2927.510 2170.850 2928.690 2172.030 ;
        RECT 2927.510 2169.250 2928.690 2170.430 ;
        RECT 2927.510 1990.850 2928.690 1992.030 ;
        RECT 2927.510 1989.250 2928.690 1990.430 ;
        RECT 2927.510 1810.850 2928.690 1812.030 ;
        RECT 2927.510 1809.250 2928.690 1810.430 ;
        RECT 2927.510 1630.850 2928.690 1632.030 ;
        RECT 2927.510 1629.250 2928.690 1630.430 ;
        RECT 2927.510 1450.850 2928.690 1452.030 ;
        RECT 2927.510 1449.250 2928.690 1450.430 ;
        RECT 2927.510 1270.850 2928.690 1272.030 ;
        RECT 2927.510 1269.250 2928.690 1270.430 ;
        RECT 2927.510 1090.850 2928.690 1092.030 ;
        RECT 2927.510 1089.250 2928.690 1090.430 ;
        RECT 2927.510 910.850 2928.690 912.030 ;
        RECT 2927.510 909.250 2928.690 910.430 ;
        RECT 2927.510 730.850 2928.690 732.030 ;
        RECT 2927.510 729.250 2928.690 730.430 ;
        RECT 2927.510 550.850 2928.690 552.030 ;
        RECT 2927.510 549.250 2928.690 550.430 ;
        RECT 2927.510 370.850 2928.690 372.030 ;
        RECT 2927.510 369.250 2928.690 370.430 ;
        RECT 2927.510 190.850 2928.690 192.030 ;
        RECT 2927.510 189.250 2928.690 190.430 ;
        RECT 2927.510 10.850 2928.690 12.030 ;
        RECT 2927.510 9.250 2928.690 10.430 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
=======
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
>>>>>>> Latest run - not LVS matched yet
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
<<<<<<< HEAD
        RECT -9.980 3432.140 -6.980 3432.150 ;
        RECT 2926.600 3432.140 2929.600 3432.150 ;
        RECT -14.680 3429.140 0.300 3432.140 ;
        RECT 2919.700 3429.140 2934.300 3432.140 ;
        RECT -9.980 3429.130 -6.980 3429.140 ;
        RECT 2926.600 3429.130 2929.600 3429.140 ;
        RECT -9.980 3252.140 -6.980 3252.150 ;
        RECT 2926.600 3252.140 2929.600 3252.150 ;
        RECT -14.680 3249.140 0.300 3252.140 ;
        RECT 2919.700 3249.140 2934.300 3252.140 ;
        RECT -9.980 3249.130 -6.980 3249.140 ;
        RECT 2926.600 3249.130 2929.600 3249.140 ;
        RECT -9.980 3072.140 -6.980 3072.150 ;
        RECT 2926.600 3072.140 2929.600 3072.150 ;
        RECT -14.680 3069.140 0.300 3072.140 ;
        RECT 2919.700 3069.140 2934.300 3072.140 ;
        RECT -9.980 3069.130 -6.980 3069.140 ;
        RECT 2926.600 3069.130 2929.600 3069.140 ;
        RECT -9.980 2892.140 -6.980 2892.150 ;
        RECT 2926.600 2892.140 2929.600 2892.150 ;
        RECT -14.680 2889.140 0.300 2892.140 ;
        RECT 2919.700 2889.140 2934.300 2892.140 ;
        RECT -9.980 2889.130 -6.980 2889.140 ;
        RECT 2926.600 2889.130 2929.600 2889.140 ;
        RECT -9.980 2712.140 -6.980 2712.150 ;
        RECT 2926.600 2712.140 2929.600 2712.150 ;
        RECT -14.680 2709.140 0.300 2712.140 ;
        RECT 2919.700 2709.140 2934.300 2712.140 ;
        RECT -9.980 2709.130 -6.980 2709.140 ;
        RECT 2926.600 2709.130 2929.600 2709.140 ;
        RECT -9.980 2532.140 -6.980 2532.150 ;
        RECT 2926.600 2532.140 2929.600 2532.150 ;
        RECT -14.680 2529.140 0.300 2532.140 ;
        RECT 2919.700 2529.140 2934.300 2532.140 ;
        RECT -9.980 2529.130 -6.980 2529.140 ;
        RECT 2926.600 2529.130 2929.600 2529.140 ;
        RECT -9.980 2352.140 -6.980 2352.150 ;
        RECT 2926.600 2352.140 2929.600 2352.150 ;
        RECT -14.680 2349.140 0.300 2352.140 ;
        RECT 2919.700 2349.140 2934.300 2352.140 ;
        RECT -9.980 2349.130 -6.980 2349.140 ;
        RECT 2926.600 2349.130 2929.600 2349.140 ;
        RECT -9.980 2172.140 -6.980 2172.150 ;
        RECT 2926.600 2172.140 2929.600 2172.150 ;
        RECT -14.680 2169.140 0.300 2172.140 ;
        RECT 2919.700 2169.140 2934.300 2172.140 ;
        RECT -9.980 2169.130 -6.980 2169.140 ;
        RECT 2926.600 2169.130 2929.600 2169.140 ;
        RECT -9.980 1992.140 -6.980 1992.150 ;
        RECT 2926.600 1992.140 2929.600 1992.150 ;
        RECT -14.680 1989.140 0.300 1992.140 ;
        RECT 2919.700 1989.140 2934.300 1992.140 ;
        RECT -9.980 1989.130 -6.980 1989.140 ;
        RECT 2926.600 1989.130 2929.600 1989.140 ;
        RECT -9.980 1812.140 -6.980 1812.150 ;
        RECT 2926.600 1812.140 2929.600 1812.150 ;
        RECT -14.680 1809.140 0.300 1812.140 ;
        RECT 2919.700 1809.140 2934.300 1812.140 ;
        RECT -9.980 1809.130 -6.980 1809.140 ;
        RECT 2926.600 1809.130 2929.600 1809.140 ;
        RECT -9.980 1632.140 -6.980 1632.150 ;
        RECT 2926.600 1632.140 2929.600 1632.150 ;
        RECT -14.680 1629.140 0.300 1632.140 ;
        RECT 2919.700 1629.140 2934.300 1632.140 ;
        RECT -9.980 1629.130 -6.980 1629.140 ;
        RECT 2926.600 1629.130 2929.600 1629.140 ;
        RECT -9.980 1452.140 -6.980 1452.150 ;
        RECT 2926.600 1452.140 2929.600 1452.150 ;
        RECT -14.680 1449.140 0.300 1452.140 ;
        RECT 2919.700 1449.140 2934.300 1452.140 ;
        RECT -9.980 1449.130 -6.980 1449.140 ;
        RECT 2926.600 1449.130 2929.600 1449.140 ;
        RECT -9.980 1272.140 -6.980 1272.150 ;
        RECT 2926.600 1272.140 2929.600 1272.150 ;
        RECT -14.680 1269.140 0.300 1272.140 ;
        RECT 2919.700 1269.140 2934.300 1272.140 ;
        RECT -9.980 1269.130 -6.980 1269.140 ;
        RECT 2926.600 1269.130 2929.600 1269.140 ;
        RECT -9.980 1092.140 -6.980 1092.150 ;
        RECT 2926.600 1092.140 2929.600 1092.150 ;
        RECT -14.680 1089.140 0.300 1092.140 ;
        RECT 2919.700 1089.140 2934.300 1092.140 ;
        RECT -9.980 1089.130 -6.980 1089.140 ;
        RECT 2926.600 1089.130 2929.600 1089.140 ;
        RECT -9.980 912.140 -6.980 912.150 ;
        RECT 2926.600 912.140 2929.600 912.150 ;
        RECT -14.680 909.140 0.300 912.140 ;
        RECT 2919.700 909.140 2934.300 912.140 ;
        RECT -9.980 909.130 -6.980 909.140 ;
        RECT 2926.600 909.130 2929.600 909.140 ;
        RECT -9.980 732.140 -6.980 732.150 ;
        RECT 2926.600 732.140 2929.600 732.150 ;
        RECT -14.680 729.140 0.300 732.140 ;
        RECT 2919.700 729.140 2934.300 732.140 ;
        RECT -9.980 729.130 -6.980 729.140 ;
        RECT 2926.600 729.130 2929.600 729.140 ;
        RECT -9.980 552.140 -6.980 552.150 ;
        RECT 2926.600 552.140 2929.600 552.150 ;
        RECT -14.680 549.140 0.300 552.140 ;
        RECT 2919.700 549.140 2934.300 552.140 ;
        RECT -9.980 549.130 -6.980 549.140 ;
        RECT 2926.600 549.130 2929.600 549.140 ;
        RECT -9.980 372.140 -6.980 372.150 ;
        RECT 2926.600 372.140 2929.600 372.150 ;
        RECT -14.680 369.140 0.300 372.140 ;
        RECT 2919.700 369.140 2934.300 372.140 ;
        RECT -9.980 369.130 -6.980 369.140 ;
        RECT 2926.600 369.130 2929.600 369.140 ;
        RECT -9.980 192.140 -6.980 192.150 ;
        RECT 2926.600 192.140 2929.600 192.150 ;
        RECT -14.680 189.140 0.300 192.140 ;
        RECT 2919.700 189.140 2934.300 192.140 ;
        RECT -9.980 189.130 -6.980 189.140 ;
        RECT 2926.600 189.130 2929.600 189.140 ;
        RECT -9.980 12.140 -6.980 12.150 ;
        RECT 2926.600 12.140 2929.600 12.150 ;
        RECT -14.680 9.140 0.300 12.140 ;
        RECT 2919.700 9.140 2934.300 12.140 ;
        RECT -9.980 9.130 -6.980 9.140 ;
        RECT 2926.600 9.130 2929.600 9.140 ;
=======
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
>>>>>>> Latest run - not LVS matched yet
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 3519.700 97.020 3529.000 ;
        RECT 274.020 3519.700 277.020 3529.000 ;
        RECT 454.020 3519.700 457.020 3529.000 ;
        RECT 634.020 3519.700 637.020 3529.000 ;
        RECT 814.020 3519.700 817.020 3529.000 ;
        RECT 994.020 3519.700 997.020 3529.000 ;
        RECT 1174.020 3519.700 1177.020 3529.000 ;
        RECT 1354.020 3519.700 1357.020 3529.000 ;
        RECT 1534.020 3519.700 1537.020 3529.000 ;
        RECT 1714.020 3519.700 1717.020 3529.000 ;
        RECT 1894.020 3519.700 1897.020 3529.000 ;
        RECT 2074.020 3519.700 2077.020 3529.000 ;
        RECT 2254.020 3519.700 2257.020 3529.000 ;
        RECT 2434.020 3519.700 2437.020 3529.000 ;
        RECT 2614.020 3519.700 2617.020 3529.000 ;
        RECT 2794.020 3519.700 2797.020 3529.000 ;
        RECT 94.020 -9.320 97.020 0.300 ;
        RECT 274.020 -9.320 277.020 0.300 ;
        RECT 454.020 -9.320 457.020 0.300 ;
        RECT 634.020 -9.320 637.020 0.300 ;
        RECT 814.020 -9.320 817.020 0.300 ;
        RECT 994.020 -9.320 997.020 0.300 ;
        RECT 1174.020 -9.320 1177.020 0.300 ;
        RECT 1354.020 -9.320 1357.020 0.300 ;
        RECT 1534.020 -9.320 1537.020 0.300 ;
        RECT 1714.020 -9.320 1717.020 0.300 ;
        RECT 1894.020 -9.320 1897.020 0.300 ;
        RECT 2074.020 -9.320 2077.020 0.300 ;
        RECT 2254.020 -9.320 2257.020 0.300 ;
        RECT 2434.020 -9.320 2437.020 0.300 ;
        RECT 2614.020 -9.320 2617.020 0.300 ;
        RECT 2794.020 -9.320 2797.020 0.300 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT -13.770 3340.850 -12.590 3342.030 ;
        RECT -13.770 3339.250 -12.590 3340.430 ;
        RECT -13.770 3160.850 -12.590 3162.030 ;
        RECT -13.770 3159.250 -12.590 3160.430 ;
        RECT -13.770 2980.850 -12.590 2982.030 ;
        RECT -13.770 2979.250 -12.590 2980.430 ;
        RECT -13.770 2800.850 -12.590 2802.030 ;
        RECT -13.770 2799.250 -12.590 2800.430 ;
        RECT -13.770 2620.850 -12.590 2622.030 ;
        RECT -13.770 2619.250 -12.590 2620.430 ;
        RECT -13.770 2440.850 -12.590 2442.030 ;
        RECT -13.770 2439.250 -12.590 2440.430 ;
        RECT -13.770 2260.850 -12.590 2262.030 ;
        RECT -13.770 2259.250 -12.590 2260.430 ;
        RECT -13.770 2080.850 -12.590 2082.030 ;
        RECT -13.770 2079.250 -12.590 2080.430 ;
        RECT -13.770 1900.850 -12.590 1902.030 ;
        RECT -13.770 1899.250 -12.590 1900.430 ;
        RECT -13.770 1720.850 -12.590 1722.030 ;
        RECT -13.770 1719.250 -12.590 1720.430 ;
        RECT -13.770 1540.850 -12.590 1542.030 ;
        RECT -13.770 1539.250 -12.590 1540.430 ;
        RECT -13.770 1360.850 -12.590 1362.030 ;
        RECT -13.770 1359.250 -12.590 1360.430 ;
        RECT -13.770 1180.850 -12.590 1182.030 ;
        RECT -13.770 1179.250 -12.590 1180.430 ;
        RECT -13.770 1000.850 -12.590 1002.030 ;
        RECT -13.770 999.250 -12.590 1000.430 ;
        RECT -13.770 820.850 -12.590 822.030 ;
        RECT -13.770 819.250 -12.590 820.430 ;
        RECT -13.770 640.850 -12.590 642.030 ;
        RECT -13.770 639.250 -12.590 640.430 ;
        RECT -13.770 460.850 -12.590 462.030 ;
        RECT -13.770 459.250 -12.590 460.430 ;
        RECT -13.770 280.850 -12.590 282.030 ;
        RECT -13.770 279.250 -12.590 280.430 ;
        RECT -13.770 100.850 -12.590 102.030 ;
        RECT -13.770 99.250 -12.590 100.430 ;
        RECT 2932.210 3340.850 2933.390 3342.030 ;
        RECT 2932.210 3339.250 2933.390 3340.430 ;
        RECT 2932.210 3160.850 2933.390 3162.030 ;
        RECT 2932.210 3159.250 2933.390 3160.430 ;
        RECT 2932.210 2980.850 2933.390 2982.030 ;
        RECT 2932.210 2979.250 2933.390 2980.430 ;
        RECT 2932.210 2800.850 2933.390 2802.030 ;
        RECT 2932.210 2799.250 2933.390 2800.430 ;
        RECT 2932.210 2620.850 2933.390 2622.030 ;
        RECT 2932.210 2619.250 2933.390 2620.430 ;
        RECT 2932.210 2440.850 2933.390 2442.030 ;
        RECT 2932.210 2439.250 2933.390 2440.430 ;
        RECT 2932.210 2260.850 2933.390 2262.030 ;
        RECT 2932.210 2259.250 2933.390 2260.430 ;
        RECT 2932.210 2080.850 2933.390 2082.030 ;
        RECT 2932.210 2079.250 2933.390 2080.430 ;
        RECT 2932.210 1900.850 2933.390 1902.030 ;
        RECT 2932.210 1899.250 2933.390 1900.430 ;
        RECT 2932.210 1720.850 2933.390 1722.030 ;
        RECT 2932.210 1719.250 2933.390 1720.430 ;
        RECT 2932.210 1540.850 2933.390 1542.030 ;
        RECT 2932.210 1539.250 2933.390 1540.430 ;
        RECT 2932.210 1360.850 2933.390 1362.030 ;
        RECT 2932.210 1359.250 2933.390 1360.430 ;
        RECT 2932.210 1180.850 2933.390 1182.030 ;
        RECT 2932.210 1179.250 2933.390 1180.430 ;
        RECT 2932.210 1000.850 2933.390 1002.030 ;
        RECT 2932.210 999.250 2933.390 1000.430 ;
        RECT 2932.210 820.850 2933.390 822.030 ;
        RECT 2932.210 819.250 2933.390 820.430 ;
        RECT 2932.210 640.850 2933.390 642.030 ;
        RECT 2932.210 639.250 2933.390 640.430 ;
        RECT 2932.210 460.850 2933.390 462.030 ;
        RECT 2932.210 459.250 2933.390 460.430 ;
        RECT 2932.210 280.850 2933.390 282.030 ;
        RECT 2932.210 279.250 2933.390 280.430 ;
        RECT 2932.210 100.850 2933.390 102.030 ;
        RECT 2932.210 99.250 2933.390 100.430 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.140 -11.680 3342.150 ;
        RECT 2931.300 3342.140 2934.300 3342.150 ;
        RECT -14.680 3339.140 0.300 3342.140 ;
        RECT 2919.700 3339.140 2934.300 3342.140 ;
        RECT -14.680 3339.130 -11.680 3339.140 ;
        RECT 2931.300 3339.130 2934.300 3339.140 ;
        RECT -14.680 3162.140 -11.680 3162.150 ;
        RECT 2931.300 3162.140 2934.300 3162.150 ;
        RECT -14.680 3159.140 0.300 3162.140 ;
        RECT 2919.700 3159.140 2934.300 3162.140 ;
        RECT -14.680 3159.130 -11.680 3159.140 ;
        RECT 2931.300 3159.130 2934.300 3159.140 ;
        RECT -14.680 2982.140 -11.680 2982.150 ;
        RECT 2931.300 2982.140 2934.300 2982.150 ;
        RECT -14.680 2979.140 0.300 2982.140 ;
        RECT 2919.700 2979.140 2934.300 2982.140 ;
        RECT -14.680 2979.130 -11.680 2979.140 ;
        RECT 2931.300 2979.130 2934.300 2979.140 ;
        RECT -14.680 2802.140 -11.680 2802.150 ;
        RECT 2931.300 2802.140 2934.300 2802.150 ;
        RECT -14.680 2799.140 0.300 2802.140 ;
        RECT 2919.700 2799.140 2934.300 2802.140 ;
        RECT -14.680 2799.130 -11.680 2799.140 ;
        RECT 2931.300 2799.130 2934.300 2799.140 ;
        RECT -14.680 2622.140 -11.680 2622.150 ;
        RECT 2931.300 2622.140 2934.300 2622.150 ;
        RECT -14.680 2619.140 0.300 2622.140 ;
        RECT 2919.700 2619.140 2934.300 2622.140 ;
        RECT -14.680 2619.130 -11.680 2619.140 ;
        RECT 2931.300 2619.130 2934.300 2619.140 ;
        RECT -14.680 2442.140 -11.680 2442.150 ;
        RECT 2931.300 2442.140 2934.300 2442.150 ;
        RECT -14.680 2439.140 0.300 2442.140 ;
        RECT 2919.700 2439.140 2934.300 2442.140 ;
        RECT -14.680 2439.130 -11.680 2439.140 ;
        RECT 2931.300 2439.130 2934.300 2439.140 ;
        RECT -14.680 2262.140 -11.680 2262.150 ;
        RECT 2931.300 2262.140 2934.300 2262.150 ;
        RECT -14.680 2259.140 0.300 2262.140 ;
        RECT 2919.700 2259.140 2934.300 2262.140 ;
        RECT -14.680 2259.130 -11.680 2259.140 ;
        RECT 2931.300 2259.130 2934.300 2259.140 ;
        RECT -14.680 2082.140 -11.680 2082.150 ;
        RECT 2931.300 2082.140 2934.300 2082.150 ;
        RECT -14.680 2079.140 0.300 2082.140 ;
        RECT 2919.700 2079.140 2934.300 2082.140 ;
        RECT -14.680 2079.130 -11.680 2079.140 ;
        RECT 2931.300 2079.130 2934.300 2079.140 ;
        RECT -14.680 1902.140 -11.680 1902.150 ;
        RECT 2931.300 1902.140 2934.300 1902.150 ;
        RECT -14.680 1899.140 0.300 1902.140 ;
        RECT 2919.700 1899.140 2934.300 1902.140 ;
        RECT -14.680 1899.130 -11.680 1899.140 ;
        RECT 2931.300 1899.130 2934.300 1899.140 ;
        RECT -14.680 1722.140 -11.680 1722.150 ;
        RECT 2931.300 1722.140 2934.300 1722.150 ;
        RECT -14.680 1719.140 0.300 1722.140 ;
        RECT 2919.700 1719.140 2934.300 1722.140 ;
        RECT -14.680 1719.130 -11.680 1719.140 ;
        RECT 2931.300 1719.130 2934.300 1719.140 ;
        RECT -14.680 1542.140 -11.680 1542.150 ;
        RECT 2931.300 1542.140 2934.300 1542.150 ;
        RECT -14.680 1539.140 0.300 1542.140 ;
        RECT 2919.700 1539.140 2934.300 1542.140 ;
        RECT -14.680 1539.130 -11.680 1539.140 ;
        RECT 2931.300 1539.130 2934.300 1539.140 ;
        RECT -14.680 1362.140 -11.680 1362.150 ;
        RECT 2931.300 1362.140 2934.300 1362.150 ;
        RECT -14.680 1359.140 0.300 1362.140 ;
        RECT 2919.700 1359.140 2934.300 1362.140 ;
        RECT -14.680 1359.130 -11.680 1359.140 ;
        RECT 2931.300 1359.130 2934.300 1359.140 ;
        RECT -14.680 1182.140 -11.680 1182.150 ;
        RECT 2931.300 1182.140 2934.300 1182.150 ;
        RECT -14.680 1179.140 0.300 1182.140 ;
        RECT 2919.700 1179.140 2934.300 1182.140 ;
        RECT -14.680 1179.130 -11.680 1179.140 ;
        RECT 2931.300 1179.130 2934.300 1179.140 ;
        RECT -14.680 1002.140 -11.680 1002.150 ;
        RECT 2931.300 1002.140 2934.300 1002.150 ;
        RECT -14.680 999.140 0.300 1002.140 ;
        RECT 2919.700 999.140 2934.300 1002.140 ;
        RECT -14.680 999.130 -11.680 999.140 ;
        RECT 2931.300 999.130 2934.300 999.140 ;
        RECT -14.680 822.140 -11.680 822.150 ;
        RECT 2931.300 822.140 2934.300 822.150 ;
        RECT -14.680 819.140 0.300 822.140 ;
        RECT 2919.700 819.140 2934.300 822.140 ;
        RECT -14.680 819.130 -11.680 819.140 ;
        RECT 2931.300 819.130 2934.300 819.140 ;
        RECT -14.680 642.140 -11.680 642.150 ;
        RECT 2931.300 642.140 2934.300 642.150 ;
        RECT -14.680 639.140 0.300 642.140 ;
        RECT 2919.700 639.140 2934.300 642.140 ;
        RECT -14.680 639.130 -11.680 639.140 ;
        RECT 2931.300 639.130 2934.300 639.140 ;
        RECT -14.680 462.140 -11.680 462.150 ;
        RECT 2931.300 462.140 2934.300 462.150 ;
        RECT -14.680 459.140 0.300 462.140 ;
        RECT 2919.700 459.140 2934.300 462.140 ;
        RECT -14.680 459.130 -11.680 459.140 ;
        RECT 2931.300 459.130 2934.300 459.140 ;
        RECT -14.680 282.140 -11.680 282.150 ;
        RECT 2931.300 282.140 2934.300 282.150 ;
        RECT -14.680 279.140 0.300 282.140 ;
        RECT 2919.700 279.140 2934.300 282.140 ;
        RECT -14.680 279.130 -11.680 279.140 ;
        RECT 2931.300 279.130 2934.300 279.140 ;
        RECT -14.680 102.140 -11.680 102.150 ;
        RECT 2931.300 102.140 2934.300 102.150 ;
        RECT -14.680 99.140 0.300 102.140 ;
        RECT 2919.700 99.140 2934.300 102.140 ;
        RECT -14.680 99.130 -11.680 99.140 ;
        RECT 2931.300 99.130 2934.300 99.140 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
=======
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 -9.220 457.020 3528.900 ;
        RECT 634.020 -9.220 637.020 3528.900 ;
        RECT 814.020 -9.220 817.020 3528.900 ;
        RECT 994.020 -9.220 997.020 3528.900 ;
        RECT 1174.020 -9.220 1177.020 3528.900 ;
        RECT 1354.020 -9.220 1357.020 3528.900 ;
        RECT 1534.020 -9.220 1537.020 3528.900 ;
        RECT 1714.020 -9.220 1717.020 3528.900 ;
        RECT 1894.020 -9.220 1897.020 3528.900 ;
        RECT 2074.020 -9.220 2077.020 3528.900 ;
        RECT 2254.020 -9.220 2257.020 3528.900 ;
        RECT 2434.020 -9.220 2437.020 3528.900 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 3519.700 25.020 3538.400 ;
        RECT 202.020 3519.700 205.020 3538.400 ;
        RECT 382.020 3519.700 385.020 3538.400 ;
        RECT 562.020 3519.700 565.020 3538.400 ;
        RECT 742.020 3519.700 745.020 3538.400 ;
        RECT 922.020 3519.700 925.020 3538.400 ;
        RECT 1102.020 3519.700 1105.020 3538.400 ;
        RECT 1282.020 3519.700 1285.020 3538.400 ;
        RECT 1462.020 3519.700 1465.020 3538.400 ;
        RECT 1642.020 3519.700 1645.020 3538.400 ;
        RECT 1822.020 3519.700 1825.020 3538.400 ;
        RECT 2002.020 3519.700 2005.020 3538.400 ;
        RECT 2182.020 3519.700 2185.020 3538.400 ;
        RECT 2362.020 3519.700 2365.020 3538.400 ;
        RECT 2542.020 3519.700 2545.020 3538.400 ;
        RECT 2722.020 3519.700 2725.020 3538.400 ;
        RECT 2902.020 3519.700 2905.020 3538.400 ;
        RECT 22.020 -18.720 25.020 0.300 ;
        RECT 202.020 -18.720 205.020 0.300 ;
        RECT 382.020 -18.720 385.020 0.300 ;
        RECT 562.020 -18.720 565.020 0.300 ;
        RECT 742.020 -18.720 745.020 0.300 ;
        RECT 922.020 -18.720 925.020 0.300 ;
        RECT 1102.020 -18.720 1105.020 0.300 ;
        RECT 1282.020 -18.720 1285.020 0.300 ;
        RECT 1462.020 -18.720 1465.020 0.300 ;
        RECT 1642.020 -18.720 1645.020 0.300 ;
        RECT 1822.020 -18.720 1825.020 0.300 ;
        RECT 2002.020 -18.720 2005.020 0.300 ;
        RECT 2182.020 -18.720 2185.020 0.300 ;
        RECT 2362.020 -18.720 2365.020 0.300 ;
        RECT 2542.020 -18.720 2545.020 0.300 ;
        RECT 2722.020 -18.720 2725.020 0.300 ;
        RECT 2902.020 -18.720 2905.020 0.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 0.300 3450.380 ;
        RECT 2919.700 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 0.300 3270.380 ;
        RECT 2919.700 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 0.300 3090.380 ;
        RECT 2919.700 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 0.300 2910.380 ;
        RECT 2919.700 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 0.300 2730.380 ;
        RECT 2919.700 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 0.300 2550.380 ;
        RECT 2919.700 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 0.300 2370.380 ;
        RECT 2919.700 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 0.300 2190.380 ;
        RECT 2919.700 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 0.300 2010.380 ;
        RECT 2919.700 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 0.300 1830.380 ;
        RECT 2919.700 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 0.300 1650.380 ;
        RECT 2919.700 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 0.300 1470.380 ;
        RECT 2919.700 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 0.300 1290.380 ;
        RECT 2919.700 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 0.300 1110.380 ;
        RECT 2919.700 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 0.300 930.380 ;
        RECT 2919.700 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 0.300 750.380 ;
        RECT 2919.700 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 0.300 570.380 ;
        RECT 2919.700 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 0.300 390.380 ;
        RECT 2919.700 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 0.300 210.380 ;
        RECT 2919.700 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 0.300 30.380 ;
        RECT 2919.700 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
=======
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 -18.420 565.020 3538.100 ;
        RECT 742.020 -18.420 745.020 3538.100 ;
        RECT 922.020 -18.420 925.020 3538.100 ;
        RECT 1102.020 -18.420 1105.020 3538.100 ;
        RECT 1282.020 -18.420 1285.020 3538.100 ;
        RECT 1462.020 -18.420 1465.020 3538.100 ;
        RECT 1642.020 -18.420 1645.020 3538.100 ;
        RECT 1822.020 -18.420 1825.020 3538.100 ;
        RECT 2002.020 -18.420 2005.020 3538.100 ;
        RECT 2182.020 -18.420 2185.020 3538.100 ;
        RECT 2362.020 -18.420 2365.020 3538.100 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 3519.700 115.020 3538.400 ;
        RECT 292.020 3519.700 295.020 3538.400 ;
        RECT 472.020 3519.700 475.020 3538.400 ;
        RECT 652.020 3519.700 655.020 3538.400 ;
        RECT 832.020 3519.700 835.020 3538.400 ;
        RECT 1012.020 3519.700 1015.020 3538.400 ;
        RECT 1192.020 3519.700 1195.020 3538.400 ;
        RECT 1372.020 3519.700 1375.020 3538.400 ;
        RECT 1552.020 3519.700 1555.020 3538.400 ;
        RECT 1732.020 3519.700 1735.020 3538.400 ;
        RECT 1912.020 3519.700 1915.020 3538.400 ;
        RECT 2092.020 3519.700 2095.020 3538.400 ;
        RECT 2272.020 3519.700 2275.020 3538.400 ;
        RECT 2452.020 3519.700 2455.020 3538.400 ;
        RECT 2632.020 3519.700 2635.020 3538.400 ;
        RECT 2812.020 3519.700 2815.020 3538.400 ;
        RECT 112.020 -18.720 115.020 0.300 ;
        RECT 292.020 -18.720 295.020 0.300 ;
        RECT 472.020 -18.720 475.020 0.300 ;
        RECT 652.020 -18.720 655.020 0.300 ;
        RECT 832.020 -18.720 835.020 0.300 ;
        RECT 1012.020 -18.720 1015.020 0.300 ;
        RECT 1192.020 -18.720 1195.020 0.300 ;
        RECT 1372.020 -18.720 1375.020 0.300 ;
        RECT 1552.020 -18.720 1555.020 0.300 ;
        RECT 1732.020 -18.720 1735.020 0.300 ;
        RECT 1912.020 -18.720 1915.020 0.300 ;
        RECT 2092.020 -18.720 2095.020 0.300 ;
        RECT 2272.020 -18.720 2275.020 0.300 ;
        RECT 2452.020 -18.720 2455.020 0.300 ;
        RECT 2632.020 -18.720 2635.020 0.300 ;
        RECT 2812.020 -18.720 2815.020 0.300 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 0.300 3360.380 ;
        RECT 2919.700 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 0.300 3180.380 ;
        RECT 2919.700 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 0.300 3000.380 ;
        RECT 2919.700 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 0.300 2820.380 ;
        RECT 2919.700 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 0.300 2640.380 ;
        RECT 2919.700 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 0.300 2460.380 ;
        RECT 2919.700 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 0.300 2280.380 ;
        RECT 2919.700 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 0.300 2100.380 ;
        RECT 2919.700 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 0.300 1920.380 ;
        RECT 2919.700 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 0.300 1740.380 ;
        RECT 2919.700 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 0.300 1560.380 ;
        RECT 2919.700 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 0.300 1380.380 ;
        RECT 2919.700 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 0.300 1200.380 ;
        RECT 2919.700 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 0.300 1020.380 ;
        RECT 2919.700 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 0.300 840.380 ;
        RECT 2919.700 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 0.300 660.380 ;
        RECT 2919.700 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 0.300 480.380 ;
        RECT 2919.700 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 0.300 300.380 ;
        RECT 2919.700 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 0.300 120.380 ;
        RECT 2919.700 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
=======
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 -18.420 475.020 3538.100 ;
        RECT 652.020 -18.420 655.020 3538.100 ;
        RECT 832.020 -18.420 835.020 3538.100 ;
        RECT 1012.020 -18.420 1015.020 3538.100 ;
        RECT 1192.020 -18.420 1195.020 3538.100 ;
        RECT 1372.020 -18.420 1375.020 3538.100 ;
        RECT 1552.020 -18.420 1555.020 3538.100 ;
        RECT 1732.020 -18.420 1735.020 3538.100 ;
        RECT 1912.020 -18.420 1915.020 3538.100 ;
        RECT 2092.020 -18.420 2095.020 3538.100 ;
        RECT 2272.020 -18.420 2275.020 3538.100 ;
        RECT 2452.020 -18.420 2455.020 3538.100 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 3519.700 43.020 3547.800 ;
        RECT 220.020 3519.700 223.020 3547.800 ;
        RECT 400.020 3519.700 403.020 3547.800 ;
        RECT 580.020 3519.700 583.020 3547.800 ;
        RECT 760.020 3519.700 763.020 3547.800 ;
        RECT 940.020 3519.700 943.020 3547.800 ;
        RECT 1120.020 3519.700 1123.020 3547.800 ;
        RECT 1300.020 3519.700 1303.020 3547.800 ;
        RECT 1480.020 3519.700 1483.020 3547.800 ;
        RECT 1660.020 3519.700 1663.020 3547.800 ;
        RECT 1840.020 3519.700 1843.020 3547.800 ;
        RECT 2020.020 3519.700 2023.020 3547.800 ;
        RECT 2200.020 3519.700 2203.020 3547.800 ;
        RECT 2380.020 3519.700 2383.020 3547.800 ;
        RECT 2560.020 3519.700 2563.020 3547.800 ;
        RECT 2740.020 3519.700 2743.020 3547.800 ;
        RECT 40.020 -28.120 43.020 0.300 ;
        RECT 220.020 -28.120 223.020 0.300 ;
        RECT 400.020 -28.120 403.020 0.300 ;
        RECT 580.020 -28.120 583.020 0.300 ;
        RECT 760.020 -28.120 763.020 0.300 ;
        RECT 940.020 -28.120 943.020 0.300 ;
        RECT 1120.020 -28.120 1123.020 0.300 ;
        RECT 1300.020 -28.120 1303.020 0.300 ;
        RECT 1480.020 -28.120 1483.020 0.300 ;
        RECT 1660.020 -28.120 1663.020 0.300 ;
        RECT 1840.020 -28.120 1843.020 0.300 ;
        RECT 2020.020 -28.120 2023.020 0.300 ;
        RECT 2200.020 -28.120 2203.020 0.300 ;
        RECT 2380.020 -28.120 2383.020 0.300 ;
        RECT 2560.020 -28.120 2563.020 0.300 ;
        RECT 2740.020 -28.120 2743.020 0.300 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 0.300 3468.380 ;
        RECT 2919.700 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 0.300 3288.380 ;
        RECT 2919.700 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 0.300 3108.380 ;
        RECT 2919.700 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 0.300 2928.380 ;
        RECT 2919.700 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 0.300 2748.380 ;
        RECT 2919.700 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 0.300 2568.380 ;
        RECT 2919.700 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 0.300 2388.380 ;
        RECT 2919.700 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 0.300 2208.380 ;
        RECT 2919.700 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 0.300 2028.380 ;
        RECT 2919.700 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 0.300 1848.380 ;
        RECT 2919.700 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 0.300 1668.380 ;
        RECT 2919.700 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 0.300 1488.380 ;
        RECT 2919.700 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 0.300 1308.380 ;
        RECT 2919.700 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 0.300 1128.380 ;
        RECT 2919.700 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 0.300 948.380 ;
        RECT 2919.700 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 0.300 768.380 ;
        RECT 2919.700 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 0.300 588.380 ;
        RECT 2919.700 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 0.300 408.380 ;
        RECT 2919.700 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 0.300 228.380 ;
        RECT 2919.700 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 0.300 48.380 ;
        RECT 2919.700 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
=======
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 -27.620 583.020 3547.300 ;
        RECT 760.020 -27.620 763.020 3547.300 ;
        RECT 940.020 -27.620 943.020 3547.300 ;
        RECT 1120.020 -27.620 1123.020 3547.300 ;
        RECT 1300.020 -27.620 1303.020 3547.300 ;
        RECT 1480.020 -27.620 1483.020 3547.300 ;
        RECT 1660.020 -27.620 1663.020 3547.300 ;
        RECT 1840.020 -27.620 1843.020 3547.300 ;
        RECT 2020.020 -27.620 2023.020 3547.300 ;
        RECT 2200.020 -27.620 2203.020 3547.300 ;
        RECT 2380.020 -27.620 2383.020 3547.300 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 3519.700 133.020 3547.800 ;
        RECT 310.020 3519.700 313.020 3547.800 ;
        RECT 490.020 3519.700 493.020 3547.800 ;
        RECT 670.020 3519.700 673.020 3547.800 ;
        RECT 850.020 3519.700 853.020 3547.800 ;
        RECT 1030.020 3519.700 1033.020 3547.800 ;
        RECT 1210.020 3519.700 1213.020 3547.800 ;
        RECT 1390.020 3519.700 1393.020 3547.800 ;
        RECT 1570.020 3519.700 1573.020 3547.800 ;
        RECT 1750.020 3519.700 1753.020 3547.800 ;
        RECT 1930.020 3519.700 1933.020 3547.800 ;
        RECT 2110.020 3519.700 2113.020 3547.800 ;
        RECT 2290.020 3519.700 2293.020 3547.800 ;
        RECT 2470.020 3519.700 2473.020 3547.800 ;
        RECT 2650.020 3519.700 2653.020 3547.800 ;
        RECT 2830.020 3519.700 2833.020 3547.800 ;
        RECT 130.020 -28.120 133.020 0.300 ;
        RECT 310.020 -28.120 313.020 0.300 ;
        RECT 490.020 -28.120 493.020 0.300 ;
        RECT 670.020 -28.120 673.020 0.300 ;
        RECT 850.020 -28.120 853.020 0.300 ;
        RECT 1030.020 -28.120 1033.020 0.300 ;
        RECT 1210.020 -28.120 1213.020 0.300 ;
        RECT 1390.020 -28.120 1393.020 0.300 ;
        RECT 1570.020 -28.120 1573.020 0.300 ;
        RECT 1750.020 -28.120 1753.020 0.300 ;
        RECT 1930.020 -28.120 1933.020 0.300 ;
        RECT 2110.020 -28.120 2113.020 0.300 ;
        RECT 2290.020 -28.120 2293.020 0.300 ;
        RECT 2470.020 -28.120 2473.020 0.300 ;
        RECT 2650.020 -28.120 2653.020 0.300 ;
        RECT 2830.020 -28.120 2833.020 0.300 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 0.300 3378.380 ;
        RECT 2919.700 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 0.300 3198.380 ;
        RECT 2919.700 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 0.300 3018.380 ;
        RECT 2919.700 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 0.300 2838.380 ;
        RECT 2919.700 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 0.300 2658.380 ;
        RECT 2919.700 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 0.300 2478.380 ;
        RECT 2919.700 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 0.300 2298.380 ;
        RECT 2919.700 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 0.300 2118.380 ;
        RECT 2919.700 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 0.300 1938.380 ;
        RECT 2919.700 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 0.300 1758.380 ;
        RECT 2919.700 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 0.300 1578.380 ;
        RECT 2919.700 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 0.300 1398.380 ;
        RECT 2919.700 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 0.300 1218.380 ;
        RECT 2919.700 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 0.300 1038.380 ;
        RECT 2919.700 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 0.300 858.380 ;
        RECT 2919.700 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 0.300 678.380 ;
        RECT 2919.700 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 0.300 498.380 ;
        RECT 2919.700 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 0.300 318.380 ;
        RECT 2919.700 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 0.300 138.380 ;
        RECT 2919.700 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 3519.700 61.020 3557.200 ;
        RECT 238.020 3519.700 241.020 3557.200 ;
        RECT 418.020 3519.700 421.020 3557.200 ;
        RECT 598.020 3519.700 601.020 3557.200 ;
        RECT 778.020 3519.700 781.020 3557.200 ;
        RECT 958.020 3519.700 961.020 3557.200 ;
        RECT 1138.020 3519.700 1141.020 3557.200 ;
        RECT 1318.020 3519.700 1321.020 3557.200 ;
        RECT 1498.020 3519.700 1501.020 3557.200 ;
        RECT 1678.020 3519.700 1681.020 3557.200 ;
        RECT 1858.020 3519.700 1861.020 3557.200 ;
        RECT 2038.020 3519.700 2041.020 3557.200 ;
        RECT 2218.020 3519.700 2221.020 3557.200 ;
        RECT 2398.020 3519.700 2401.020 3557.200 ;
        RECT 2578.020 3519.700 2581.020 3557.200 ;
        RECT 2758.020 3519.700 2761.020 3557.200 ;
        RECT 58.020 -37.520 61.020 0.300 ;
        RECT 238.020 -37.520 241.020 0.300 ;
        RECT 418.020 -37.520 421.020 0.300 ;
        RECT 598.020 -37.520 601.020 0.300 ;
        RECT 778.020 -37.520 781.020 0.300 ;
        RECT 958.020 -37.520 961.020 0.300 ;
        RECT 1138.020 -37.520 1141.020 0.300 ;
        RECT 1318.020 -37.520 1321.020 0.300 ;
        RECT 1498.020 -37.520 1501.020 0.300 ;
        RECT 1678.020 -37.520 1681.020 0.300 ;
        RECT 1858.020 -37.520 1861.020 0.300 ;
        RECT 2038.020 -37.520 2041.020 0.300 ;
        RECT 2218.020 -37.520 2221.020 0.300 ;
        RECT 2398.020 -37.520 2401.020 0.300 ;
        RECT 2578.020 -37.520 2581.020 0.300 ;
        RECT 2758.020 -37.520 2761.020 0.300 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 0.300 3486.380 ;
        RECT 2919.700 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 0.300 3306.380 ;
        RECT 2919.700 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 0.300 3126.380 ;
        RECT 2919.700 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 0.300 2946.380 ;
        RECT 2919.700 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 0.300 2766.380 ;
        RECT 2919.700 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 0.300 2586.380 ;
        RECT 2919.700 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 0.300 2406.380 ;
        RECT 2919.700 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 0.300 2226.380 ;
        RECT 2919.700 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 0.300 2046.380 ;
        RECT 2919.700 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 0.300 1866.380 ;
        RECT 2919.700 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 0.300 1686.380 ;
        RECT 2919.700 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 0.300 1506.380 ;
        RECT 2919.700 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 0.300 1326.380 ;
        RECT 2919.700 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 0.300 1146.380 ;
        RECT 2919.700 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 0.300 966.380 ;
        RECT 2919.700 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 0.300 786.380 ;
        RECT 2919.700 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 0.300 606.380 ;
        RECT 2919.700 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 0.300 426.380 ;
        RECT 2919.700 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 0.300 246.380 ;
        RECT 2919.700 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 0.300 66.380 ;
        RECT 2919.700 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
=======
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 -27.620 493.020 3547.300 ;
        RECT 670.020 -27.620 673.020 3547.300 ;
        RECT 850.020 -27.620 853.020 3547.300 ;
        RECT 1030.020 -27.620 1033.020 3547.300 ;
        RECT 1210.020 -27.620 1213.020 3547.300 ;
        RECT 1390.020 -27.620 1393.020 3547.300 ;
        RECT 1570.020 -27.620 1573.020 3547.300 ;
        RECT 1750.020 -27.620 1753.020 3547.300 ;
        RECT 1930.020 -27.620 1933.020 3547.300 ;
        RECT 2110.020 -27.620 2113.020 3547.300 ;
        RECT 2290.020 -27.620 2293.020 3547.300 ;
        RECT 2470.020 -27.620 2473.020 3547.300 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 -36.820 421.020 3556.500 ;
        RECT 598.020 -36.820 601.020 3556.500 ;
        RECT 778.020 -36.820 781.020 3556.500 ;
        RECT 958.020 -36.820 961.020 3556.500 ;
        RECT 1138.020 -36.820 1141.020 3556.500 ;
        RECT 1318.020 -36.820 1321.020 3556.500 ;
        RECT 1498.020 -36.820 1501.020 3556.500 ;
        RECT 1678.020 -36.820 1681.020 3556.500 ;
        RECT 1858.020 -36.820 1861.020 3556.500 ;
        RECT 2038.020 -36.820 2041.020 3556.500 ;
        RECT 2218.020 -36.820 2221.020 3556.500 ;
        RECT 2398.020 -36.820 2401.020 3556.500 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 3519.700 151.020 3557.200 ;
        RECT 328.020 3519.700 331.020 3557.200 ;
        RECT 508.020 3519.700 511.020 3557.200 ;
        RECT 688.020 3519.700 691.020 3557.200 ;
        RECT 868.020 3519.700 871.020 3557.200 ;
        RECT 1048.020 3519.700 1051.020 3557.200 ;
        RECT 1228.020 3519.700 1231.020 3557.200 ;
        RECT 1408.020 3519.700 1411.020 3557.200 ;
        RECT 1588.020 3519.700 1591.020 3557.200 ;
        RECT 1768.020 3519.700 1771.020 3557.200 ;
        RECT 1948.020 3519.700 1951.020 3557.200 ;
        RECT 2128.020 3519.700 2131.020 3557.200 ;
        RECT 2308.020 3519.700 2311.020 3557.200 ;
        RECT 2488.020 3519.700 2491.020 3557.200 ;
        RECT 2668.020 3519.700 2671.020 3557.200 ;
        RECT 2848.020 3519.700 2851.020 3557.200 ;
        RECT 148.020 -37.520 151.020 0.300 ;
        RECT 328.020 -37.520 331.020 0.300 ;
        RECT 508.020 -37.520 511.020 0.300 ;
        RECT 688.020 -37.520 691.020 0.300 ;
        RECT 868.020 -37.520 871.020 0.300 ;
        RECT 1048.020 -37.520 1051.020 0.300 ;
        RECT 1228.020 -37.520 1231.020 0.300 ;
        RECT 1408.020 -37.520 1411.020 0.300 ;
        RECT 1588.020 -37.520 1591.020 0.300 ;
        RECT 1768.020 -37.520 1771.020 0.300 ;
        RECT 1948.020 -37.520 1951.020 0.300 ;
        RECT 2128.020 -37.520 2131.020 0.300 ;
        RECT 2308.020 -37.520 2311.020 0.300 ;
        RECT 2488.020 -37.520 2491.020 0.300 ;
        RECT 2668.020 -37.520 2671.020 0.300 ;
        RECT 2848.020 -37.520 2851.020 0.300 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 0.300 3396.380 ;
        RECT 2919.700 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 0.300 3216.380 ;
        RECT 2919.700 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 0.300 3036.380 ;
        RECT 2919.700 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 0.300 2856.380 ;
        RECT 2919.700 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 0.300 2676.380 ;
        RECT 2919.700 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 0.300 2496.380 ;
        RECT 2919.700 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 0.300 2316.380 ;
        RECT 2919.700 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 0.300 2136.380 ;
        RECT 2919.700 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 0.300 1956.380 ;
        RECT 2919.700 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 0.300 1776.380 ;
        RECT 2919.700 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 0.300 1596.380 ;
        RECT 2919.700 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 0.300 1416.380 ;
        RECT 2919.700 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 0.300 1236.380 ;
        RECT 2919.700 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 0.300 1056.380 ;
        RECT 2919.700 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 0.300 876.380 ;
        RECT 2919.700 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 0.300 696.380 ;
        RECT 2919.700 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 0.300 516.380 ;
        RECT 2919.700 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 0.300 336.380 ;
        RECT 2919.700 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 0.300 156.380 ;
        RECT 2919.700 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
=======
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 -36.820 511.020 3556.500 ;
        RECT 688.020 -36.820 691.020 3556.500 ;
        RECT 868.020 -36.820 871.020 3556.500 ;
        RECT 1048.020 -36.820 1051.020 3556.500 ;
        RECT 1228.020 -36.820 1231.020 3556.500 ;
        RECT 1408.020 -36.820 1411.020 3556.500 ;
        RECT 1588.020 -36.820 1591.020 3556.500 ;
        RECT 1768.020 -36.820 1771.020 3556.500 ;
        RECT 1948.020 -36.820 1951.020 3556.500 ;
        RECT 2128.020 -36.820 2131.020 3556.500 ;
        RECT 2308.020 -36.820 2311.020 3556.500 ;
        RECT 2488.020 -36.820 2491.020 3556.500 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vssa2
  OBS
      LAYER li1 ;
<<<<<<< HEAD
        RECT 276.145 2.805 2799.415 3477.435 ;
      LAYER met1 ;
        RECT 2.830 2.760 2914.100 3512.160 ;
      LAYER met2 ;
        RECT 2.710 0.300 2917.370 3519.700 ;
      LAYER met3 ;
        RECT 0.300 10.715 2919.700 3508.965 ;
      LAYER met4 ;
        RECT 4.020 0.300 2905.020 3519.700 ;
      LAYER met5 ;
        RECT 0.300 9.130 2919.700 3486.390 ;
=======
        RECT 1155.520 1710.795 1944.420 2488.885 ;
      LAYER met1 ;
        RECT 1153.290 1709.220 1946.650 2489.780 ;
      LAYER met2 ;
        RECT 1150.550 2495.720 1153.030 2496.010 ;
        RECT 1153.870 2495.720 1159.470 2496.010 ;
        RECT 1160.310 2495.720 1165.910 2496.010 ;
        RECT 1166.750 2495.720 1172.810 2496.010 ;
        RECT 1173.650 2495.720 1179.250 2496.010 ;
        RECT 1180.090 2495.720 1185.690 2496.010 ;
        RECT 1186.530 2495.720 1192.590 2496.010 ;
        RECT 1193.430 2495.720 1199.030 2496.010 ;
        RECT 1199.870 2495.720 1205.470 2496.010 ;
        RECT 1206.310 2495.720 1212.370 2496.010 ;
        RECT 1213.210 2495.720 1218.810 2496.010 ;
        RECT 1219.650 2495.720 1225.710 2496.010 ;
        RECT 1226.550 2495.720 1232.150 2496.010 ;
        RECT 1232.990 2495.720 1238.590 2496.010 ;
        RECT 1239.430 2495.720 1245.490 2496.010 ;
        RECT 1246.330 2495.720 1251.930 2496.010 ;
        RECT 1252.770 2495.720 1258.370 2496.010 ;
        RECT 1259.210 2495.720 1265.270 2496.010 ;
        RECT 1266.110 2495.720 1271.710 2496.010 ;
        RECT 1272.550 2495.720 1278.610 2496.010 ;
        RECT 1279.450 2495.720 1285.050 2496.010 ;
        RECT 1285.890 2495.720 1291.490 2496.010 ;
        RECT 1292.330 2495.720 1298.390 2496.010 ;
        RECT 1299.230 2495.720 1304.830 2496.010 ;
        RECT 1305.670 2495.720 1311.270 2496.010 ;
        RECT 1312.110 2495.720 1318.170 2496.010 ;
        RECT 1319.010 2495.720 1324.610 2496.010 ;
        RECT 1325.450 2495.720 1331.510 2496.010 ;
        RECT 1332.350 2495.720 1337.950 2496.010 ;
        RECT 1338.790 2495.720 1344.390 2496.010 ;
        RECT 1345.230 2495.720 1351.290 2496.010 ;
        RECT 1352.130 2495.720 1357.730 2496.010 ;
        RECT 1358.570 2495.720 1364.170 2496.010 ;
        RECT 1365.010 2495.720 1371.070 2496.010 ;
        RECT 1371.910 2495.720 1377.510 2496.010 ;
        RECT 1378.350 2495.720 1384.410 2496.010 ;
        RECT 1385.250 2495.720 1390.850 2496.010 ;
        RECT 1391.690 2495.720 1397.290 2496.010 ;
        RECT 1398.130 2495.720 1404.190 2496.010 ;
        RECT 1405.030 2495.720 1410.630 2496.010 ;
        RECT 1411.470 2495.720 1417.070 2496.010 ;
        RECT 1417.910 2495.720 1423.970 2496.010 ;
        RECT 1424.810 2495.720 1430.410 2496.010 ;
        RECT 1431.250 2495.720 1436.850 2496.010 ;
        RECT 1437.690 2495.720 1443.750 2496.010 ;
        RECT 1444.590 2495.720 1450.190 2496.010 ;
        RECT 1451.030 2495.720 1457.090 2496.010 ;
        RECT 1457.930 2495.720 1463.530 2496.010 ;
        RECT 1464.370 2495.720 1469.970 2496.010 ;
        RECT 1470.810 2495.720 1476.870 2496.010 ;
        RECT 1477.710 2495.720 1483.310 2496.010 ;
        RECT 1484.150 2495.720 1489.750 2496.010 ;
        RECT 1490.590 2495.720 1496.650 2496.010 ;
        RECT 1497.490 2495.720 1503.090 2496.010 ;
        RECT 1503.930 2495.720 1509.990 2496.010 ;
        RECT 1510.830 2495.720 1516.430 2496.010 ;
        RECT 1517.270 2495.720 1522.870 2496.010 ;
        RECT 1523.710 2495.720 1529.770 2496.010 ;
        RECT 1530.610 2495.720 1536.210 2496.010 ;
        RECT 1537.050 2495.720 1542.650 2496.010 ;
        RECT 1543.490 2495.720 1549.550 2496.010 ;
        RECT 1550.390 2495.720 1555.990 2496.010 ;
        RECT 1556.830 2495.720 1562.890 2496.010 ;
        RECT 1563.730 2495.720 1569.330 2496.010 ;
        RECT 1570.170 2495.720 1575.770 2496.010 ;
        RECT 1576.610 2495.720 1582.670 2496.010 ;
        RECT 1583.510 2495.720 1589.110 2496.010 ;
        RECT 1589.950 2495.720 1595.550 2496.010 ;
        RECT 1596.390 2495.720 1602.450 2496.010 ;
        RECT 1603.290 2495.720 1608.890 2496.010 ;
        RECT 1609.730 2495.720 1615.790 2496.010 ;
        RECT 1616.630 2495.720 1622.230 2496.010 ;
        RECT 1623.070 2495.720 1628.670 2496.010 ;
        RECT 1629.510 2495.720 1635.570 2496.010 ;
        RECT 1636.410 2495.720 1642.010 2496.010 ;
        RECT 1642.850 2495.720 1648.450 2496.010 ;
        RECT 1649.290 2495.720 1655.350 2496.010 ;
        RECT 1656.190 2495.720 1661.790 2496.010 ;
        RECT 1662.630 2495.720 1668.690 2496.010 ;
        RECT 1669.530 2495.720 1675.130 2496.010 ;
        RECT 1675.970 2495.720 1681.570 2496.010 ;
        RECT 1682.410 2495.720 1688.470 2496.010 ;
        RECT 1689.310 2495.720 1694.910 2496.010 ;
        RECT 1695.750 2495.720 1701.350 2496.010 ;
        RECT 1702.190 2495.720 1708.250 2496.010 ;
        RECT 1709.090 2495.720 1714.690 2496.010 ;
        RECT 1715.530 2495.720 1721.130 2496.010 ;
        RECT 1721.970 2495.720 1728.030 2496.010 ;
        RECT 1728.870 2495.720 1734.470 2496.010 ;
        RECT 1735.310 2495.720 1741.370 2496.010 ;
        RECT 1742.210 2495.720 1747.810 2496.010 ;
        RECT 1748.650 2495.720 1754.250 2496.010 ;
        RECT 1755.090 2495.720 1761.150 2496.010 ;
        RECT 1761.990 2495.720 1767.590 2496.010 ;
        RECT 1768.430 2495.720 1774.030 2496.010 ;
        RECT 1774.870 2495.720 1780.930 2496.010 ;
        RECT 1781.770 2495.720 1787.370 2496.010 ;
        RECT 1788.210 2495.720 1794.270 2496.010 ;
        RECT 1795.110 2495.720 1800.710 2496.010 ;
        RECT 1801.550 2495.720 1807.150 2496.010 ;
        RECT 1807.990 2495.720 1814.050 2496.010 ;
        RECT 1814.890 2495.720 1820.490 2496.010 ;
        RECT 1821.330 2495.720 1826.930 2496.010 ;
        RECT 1827.770 2495.720 1833.830 2496.010 ;
        RECT 1834.670 2495.720 1840.270 2496.010 ;
        RECT 1841.110 2495.720 1847.170 2496.010 ;
        RECT 1848.010 2495.720 1853.610 2496.010 ;
        RECT 1854.450 2495.720 1860.050 2496.010 ;
        RECT 1860.890 2495.720 1866.950 2496.010 ;
        RECT 1867.790 2495.720 1873.390 2496.010 ;
        RECT 1874.230 2495.720 1879.830 2496.010 ;
        RECT 1880.670 2495.720 1886.730 2496.010 ;
        RECT 1887.570 2495.720 1893.170 2496.010 ;
        RECT 1894.010 2495.720 1900.070 2496.010 ;
        RECT 1900.910 2495.720 1906.510 2496.010 ;
        RECT 1907.350 2495.720 1912.950 2496.010 ;
        RECT 1913.790 2495.720 1919.850 2496.010 ;
        RECT 1920.690 2495.720 1926.290 2496.010 ;
        RECT 1927.130 2495.720 1932.730 2496.010 ;
        RECT 1933.570 2495.720 1939.630 2496.010 ;
        RECT 1940.470 2495.720 1946.070 2496.010 ;
        RECT 1150.550 1704.280 1946.620 2495.720 ;
        RECT 1151.110 1704.000 1151.650 1704.280 ;
        RECT 1152.490 1704.000 1153.030 1704.280 ;
        RECT 1153.870 1704.000 1154.870 1704.280 ;
        RECT 1155.710 1704.000 1156.250 1704.280 ;
        RECT 1157.090 1704.000 1158.090 1704.280 ;
        RECT 1158.930 1704.000 1159.470 1704.280 ;
        RECT 1160.310 1704.000 1161.310 1704.280 ;
        RECT 1162.150 1704.000 1162.690 1704.280 ;
        RECT 1163.530 1704.000 1164.530 1704.280 ;
        RECT 1165.370 1704.000 1165.910 1704.280 ;
        RECT 1166.750 1704.000 1167.750 1704.280 ;
        RECT 1168.590 1704.000 1169.130 1704.280 ;
        RECT 1169.970 1704.000 1170.970 1704.280 ;
        RECT 1171.810 1704.000 1172.350 1704.280 ;
        RECT 1173.190 1704.000 1174.190 1704.280 ;
        RECT 1175.030 1704.000 1175.570 1704.280 ;
        RECT 1176.410 1704.000 1177.410 1704.280 ;
        RECT 1178.250 1704.000 1178.790 1704.280 ;
        RECT 1179.630 1704.000 1180.630 1704.280 ;
        RECT 1181.470 1704.000 1182.010 1704.280 ;
        RECT 1182.850 1704.000 1183.850 1704.280 ;
        RECT 1184.690 1704.000 1185.230 1704.280 ;
        RECT 1186.070 1704.000 1187.070 1704.280 ;
        RECT 1187.910 1704.000 1188.450 1704.280 ;
        RECT 1189.290 1704.000 1190.290 1704.280 ;
        RECT 1191.130 1704.000 1191.670 1704.280 ;
        RECT 1192.510 1704.000 1193.510 1704.280 ;
        RECT 1194.350 1704.000 1194.890 1704.280 ;
        RECT 1195.730 1704.000 1196.730 1704.280 ;
        RECT 1197.570 1704.000 1198.110 1704.280 ;
        RECT 1198.950 1704.000 1199.950 1704.280 ;
        RECT 1200.790 1704.000 1201.330 1704.280 ;
        RECT 1202.170 1704.000 1203.170 1704.280 ;
        RECT 1204.010 1704.000 1204.550 1704.280 ;
        RECT 1205.390 1704.000 1206.390 1704.280 ;
        RECT 1207.230 1704.000 1207.770 1704.280 ;
        RECT 1208.610 1704.000 1209.610 1704.280 ;
        RECT 1210.450 1704.000 1210.990 1704.280 ;
        RECT 1211.830 1704.000 1212.830 1704.280 ;
        RECT 1213.670 1704.000 1214.210 1704.280 ;
        RECT 1215.050 1704.000 1216.050 1704.280 ;
        RECT 1216.890 1704.000 1217.430 1704.280 ;
        RECT 1218.270 1704.000 1219.270 1704.280 ;
        RECT 1220.110 1704.000 1220.650 1704.280 ;
        RECT 1221.490 1704.000 1222.490 1704.280 ;
        RECT 1223.330 1704.000 1223.870 1704.280 ;
        RECT 1224.710 1704.000 1225.710 1704.280 ;
        RECT 1226.550 1704.000 1227.090 1704.280 ;
        RECT 1227.930 1704.000 1228.930 1704.280 ;
        RECT 1229.770 1704.000 1230.310 1704.280 ;
        RECT 1231.150 1704.000 1232.150 1704.280 ;
        RECT 1232.990 1704.000 1233.530 1704.280 ;
        RECT 1234.370 1704.000 1235.370 1704.280 ;
        RECT 1236.210 1704.000 1236.750 1704.280 ;
        RECT 1237.590 1704.000 1238.590 1704.280 ;
        RECT 1239.430 1704.000 1239.970 1704.280 ;
        RECT 1240.810 1704.000 1241.810 1704.280 ;
        RECT 1242.650 1704.000 1243.190 1704.280 ;
        RECT 1244.030 1704.000 1245.030 1704.280 ;
        RECT 1245.870 1704.000 1246.410 1704.280 ;
        RECT 1247.250 1704.000 1248.250 1704.280 ;
        RECT 1249.090 1704.000 1249.630 1704.280 ;
        RECT 1250.470 1704.000 1251.010 1704.280 ;
        RECT 1251.850 1704.000 1252.850 1704.280 ;
        RECT 1253.690 1704.000 1254.230 1704.280 ;
        RECT 1255.070 1704.000 1256.070 1704.280 ;
        RECT 1256.910 1704.000 1257.450 1704.280 ;
        RECT 1258.290 1704.000 1259.290 1704.280 ;
        RECT 1260.130 1704.000 1260.670 1704.280 ;
        RECT 1261.510 1704.000 1262.510 1704.280 ;
        RECT 1263.350 1704.000 1263.890 1704.280 ;
        RECT 1264.730 1704.000 1265.730 1704.280 ;
        RECT 1266.570 1704.000 1267.110 1704.280 ;
        RECT 1267.950 1704.000 1268.950 1704.280 ;
        RECT 1269.790 1704.000 1270.330 1704.280 ;
        RECT 1271.170 1704.000 1272.170 1704.280 ;
        RECT 1273.010 1704.000 1273.550 1704.280 ;
        RECT 1274.390 1704.000 1275.390 1704.280 ;
        RECT 1276.230 1704.000 1276.770 1704.280 ;
        RECT 1277.610 1704.000 1278.610 1704.280 ;
        RECT 1279.450 1704.000 1279.990 1704.280 ;
        RECT 1280.830 1704.000 1281.830 1704.280 ;
        RECT 1282.670 1704.000 1283.210 1704.280 ;
        RECT 1284.050 1704.000 1285.050 1704.280 ;
        RECT 1285.890 1704.000 1286.430 1704.280 ;
        RECT 1287.270 1704.000 1288.270 1704.280 ;
        RECT 1289.110 1704.000 1289.650 1704.280 ;
        RECT 1290.490 1704.000 1291.490 1704.280 ;
        RECT 1292.330 1704.000 1292.870 1704.280 ;
        RECT 1293.710 1704.000 1294.710 1704.280 ;
        RECT 1295.550 1704.000 1296.090 1704.280 ;
        RECT 1296.930 1704.000 1297.930 1704.280 ;
        RECT 1298.770 1704.000 1299.310 1704.280 ;
        RECT 1300.150 1704.000 1301.150 1704.280 ;
        RECT 1301.990 1704.000 1302.530 1704.280 ;
        RECT 1303.370 1704.000 1304.370 1704.280 ;
        RECT 1305.210 1704.000 1305.750 1704.280 ;
        RECT 1306.590 1704.000 1307.590 1704.280 ;
        RECT 1308.430 1704.000 1308.970 1704.280 ;
        RECT 1309.810 1704.000 1310.810 1704.280 ;
        RECT 1311.650 1704.000 1312.190 1704.280 ;
        RECT 1313.030 1704.000 1314.030 1704.280 ;
        RECT 1314.870 1704.000 1315.410 1704.280 ;
        RECT 1316.250 1704.000 1317.250 1704.280 ;
        RECT 1318.090 1704.000 1318.630 1704.280 ;
        RECT 1319.470 1704.000 1320.470 1704.280 ;
        RECT 1321.310 1704.000 1321.850 1704.280 ;
        RECT 1322.690 1704.000 1323.690 1704.280 ;
        RECT 1324.530 1704.000 1325.070 1704.280 ;
        RECT 1325.910 1704.000 1326.910 1704.280 ;
        RECT 1327.750 1704.000 1328.290 1704.280 ;
        RECT 1329.130 1704.000 1330.130 1704.280 ;
        RECT 1330.970 1704.000 1331.510 1704.280 ;
        RECT 1332.350 1704.000 1333.350 1704.280 ;
        RECT 1334.190 1704.000 1334.730 1704.280 ;
        RECT 1335.570 1704.000 1336.570 1704.280 ;
        RECT 1337.410 1704.000 1337.950 1704.280 ;
        RECT 1338.790 1704.000 1339.790 1704.280 ;
        RECT 1340.630 1704.000 1341.170 1704.280 ;
        RECT 1342.010 1704.000 1343.010 1704.280 ;
        RECT 1343.850 1704.000 1344.390 1704.280 ;
        RECT 1345.230 1704.000 1346.230 1704.280 ;
        RECT 1347.070 1704.000 1347.610 1704.280 ;
        RECT 1348.450 1704.000 1349.450 1704.280 ;
        RECT 1350.290 1704.000 1350.830 1704.280 ;
        RECT 1351.670 1704.000 1352.210 1704.280 ;
        RECT 1353.050 1704.000 1354.050 1704.280 ;
        RECT 1354.890 1704.000 1355.430 1704.280 ;
        RECT 1356.270 1704.000 1357.270 1704.280 ;
        RECT 1358.110 1704.000 1358.650 1704.280 ;
        RECT 1359.490 1704.000 1360.490 1704.280 ;
        RECT 1361.330 1704.000 1361.870 1704.280 ;
        RECT 1362.710 1704.000 1363.710 1704.280 ;
        RECT 1364.550 1704.000 1365.090 1704.280 ;
        RECT 1365.930 1704.000 1366.930 1704.280 ;
        RECT 1367.770 1704.000 1368.310 1704.280 ;
        RECT 1369.150 1704.000 1370.150 1704.280 ;
        RECT 1370.990 1704.000 1371.530 1704.280 ;
        RECT 1372.370 1704.000 1373.370 1704.280 ;
        RECT 1374.210 1704.000 1374.750 1704.280 ;
        RECT 1375.590 1704.000 1376.590 1704.280 ;
        RECT 1377.430 1704.000 1377.970 1704.280 ;
        RECT 1378.810 1704.000 1379.810 1704.280 ;
        RECT 1380.650 1704.000 1381.190 1704.280 ;
        RECT 1382.030 1704.000 1383.030 1704.280 ;
        RECT 1383.870 1704.000 1384.410 1704.280 ;
        RECT 1385.250 1704.000 1386.250 1704.280 ;
        RECT 1387.090 1704.000 1387.630 1704.280 ;
        RECT 1388.470 1704.000 1389.470 1704.280 ;
        RECT 1390.310 1704.000 1390.850 1704.280 ;
        RECT 1391.690 1704.000 1392.690 1704.280 ;
        RECT 1393.530 1704.000 1394.070 1704.280 ;
        RECT 1394.910 1704.000 1395.910 1704.280 ;
        RECT 1396.750 1704.000 1397.290 1704.280 ;
        RECT 1398.130 1704.000 1399.130 1704.280 ;
        RECT 1399.970 1704.000 1400.510 1704.280 ;
        RECT 1401.350 1704.000 1402.350 1704.280 ;
        RECT 1403.190 1704.000 1403.730 1704.280 ;
        RECT 1404.570 1704.000 1405.570 1704.280 ;
        RECT 1406.410 1704.000 1406.950 1704.280 ;
        RECT 1407.790 1704.000 1408.790 1704.280 ;
        RECT 1409.630 1704.000 1410.170 1704.280 ;
        RECT 1411.010 1704.000 1412.010 1704.280 ;
        RECT 1412.850 1704.000 1413.390 1704.280 ;
        RECT 1414.230 1704.000 1415.230 1704.280 ;
        RECT 1416.070 1704.000 1416.610 1704.280 ;
        RECT 1417.450 1704.000 1418.450 1704.280 ;
        RECT 1419.290 1704.000 1419.830 1704.280 ;
        RECT 1420.670 1704.000 1421.670 1704.280 ;
        RECT 1422.510 1704.000 1423.050 1704.280 ;
        RECT 1423.890 1704.000 1424.890 1704.280 ;
        RECT 1425.730 1704.000 1426.270 1704.280 ;
        RECT 1427.110 1704.000 1428.110 1704.280 ;
        RECT 1428.950 1704.000 1429.490 1704.280 ;
        RECT 1430.330 1704.000 1431.330 1704.280 ;
        RECT 1432.170 1704.000 1432.710 1704.280 ;
        RECT 1433.550 1704.000 1434.550 1704.280 ;
        RECT 1435.390 1704.000 1435.930 1704.280 ;
        RECT 1436.770 1704.000 1437.770 1704.280 ;
        RECT 1438.610 1704.000 1439.150 1704.280 ;
        RECT 1439.990 1704.000 1440.990 1704.280 ;
        RECT 1441.830 1704.000 1442.370 1704.280 ;
        RECT 1443.210 1704.000 1444.210 1704.280 ;
        RECT 1445.050 1704.000 1445.590 1704.280 ;
        RECT 1446.430 1704.000 1447.430 1704.280 ;
        RECT 1448.270 1704.000 1448.810 1704.280 ;
        RECT 1449.650 1704.000 1450.190 1704.280 ;
        RECT 1451.030 1704.000 1452.030 1704.280 ;
        RECT 1452.870 1704.000 1453.410 1704.280 ;
        RECT 1454.250 1704.000 1455.250 1704.280 ;
        RECT 1456.090 1704.000 1456.630 1704.280 ;
        RECT 1457.470 1704.000 1458.470 1704.280 ;
        RECT 1459.310 1704.000 1459.850 1704.280 ;
        RECT 1460.690 1704.000 1461.690 1704.280 ;
        RECT 1462.530 1704.000 1463.070 1704.280 ;
        RECT 1463.910 1704.000 1464.910 1704.280 ;
        RECT 1465.750 1704.000 1466.290 1704.280 ;
        RECT 1467.130 1704.000 1468.130 1704.280 ;
        RECT 1468.970 1704.000 1469.510 1704.280 ;
        RECT 1470.350 1704.000 1471.350 1704.280 ;
        RECT 1472.190 1704.000 1472.730 1704.280 ;
        RECT 1473.570 1704.000 1474.570 1704.280 ;
        RECT 1475.410 1704.000 1475.950 1704.280 ;
        RECT 1476.790 1704.000 1477.790 1704.280 ;
        RECT 1478.630 1704.000 1479.170 1704.280 ;
        RECT 1480.010 1704.000 1481.010 1704.280 ;
        RECT 1481.850 1704.000 1482.390 1704.280 ;
        RECT 1483.230 1704.000 1484.230 1704.280 ;
        RECT 1485.070 1704.000 1485.610 1704.280 ;
        RECT 1486.450 1704.000 1487.450 1704.280 ;
        RECT 1488.290 1704.000 1488.830 1704.280 ;
        RECT 1489.670 1704.000 1490.670 1704.280 ;
        RECT 1491.510 1704.000 1492.050 1704.280 ;
        RECT 1492.890 1704.000 1493.890 1704.280 ;
        RECT 1494.730 1704.000 1495.270 1704.280 ;
        RECT 1496.110 1704.000 1497.110 1704.280 ;
        RECT 1497.950 1704.000 1498.490 1704.280 ;
        RECT 1499.330 1704.000 1500.330 1704.280 ;
        RECT 1501.170 1704.000 1501.710 1704.280 ;
        RECT 1502.550 1704.000 1503.550 1704.280 ;
        RECT 1504.390 1704.000 1504.930 1704.280 ;
        RECT 1505.770 1704.000 1506.770 1704.280 ;
        RECT 1507.610 1704.000 1508.150 1704.280 ;
        RECT 1508.990 1704.000 1509.990 1704.280 ;
        RECT 1510.830 1704.000 1511.370 1704.280 ;
        RECT 1512.210 1704.000 1513.210 1704.280 ;
        RECT 1514.050 1704.000 1514.590 1704.280 ;
        RECT 1515.430 1704.000 1516.430 1704.280 ;
        RECT 1517.270 1704.000 1517.810 1704.280 ;
        RECT 1518.650 1704.000 1519.650 1704.280 ;
        RECT 1520.490 1704.000 1521.030 1704.280 ;
        RECT 1521.870 1704.000 1522.870 1704.280 ;
        RECT 1523.710 1704.000 1524.250 1704.280 ;
        RECT 1525.090 1704.000 1526.090 1704.280 ;
        RECT 1526.930 1704.000 1527.470 1704.280 ;
        RECT 1528.310 1704.000 1529.310 1704.280 ;
        RECT 1530.150 1704.000 1530.690 1704.280 ;
        RECT 1531.530 1704.000 1532.530 1704.280 ;
        RECT 1533.370 1704.000 1533.910 1704.280 ;
        RECT 1534.750 1704.000 1535.750 1704.280 ;
        RECT 1536.590 1704.000 1537.130 1704.280 ;
        RECT 1537.970 1704.000 1538.970 1704.280 ;
        RECT 1539.810 1704.000 1540.350 1704.280 ;
        RECT 1541.190 1704.000 1542.190 1704.280 ;
        RECT 1543.030 1704.000 1543.570 1704.280 ;
        RECT 1544.410 1704.000 1545.410 1704.280 ;
        RECT 1546.250 1704.000 1546.790 1704.280 ;
        RECT 1547.630 1704.000 1548.630 1704.280 ;
        RECT 1549.470 1704.000 1550.010 1704.280 ;
        RECT 1550.850 1704.000 1551.390 1704.280 ;
        RECT 1552.230 1704.000 1553.230 1704.280 ;
        RECT 1554.070 1704.000 1554.610 1704.280 ;
        RECT 1555.450 1704.000 1556.450 1704.280 ;
        RECT 1557.290 1704.000 1557.830 1704.280 ;
        RECT 1558.670 1704.000 1559.670 1704.280 ;
        RECT 1560.510 1704.000 1561.050 1704.280 ;
        RECT 1561.890 1704.000 1562.890 1704.280 ;
        RECT 1563.730 1704.000 1564.270 1704.280 ;
        RECT 1565.110 1704.000 1566.110 1704.280 ;
        RECT 1566.950 1704.000 1567.490 1704.280 ;
        RECT 1568.330 1704.000 1569.330 1704.280 ;
        RECT 1570.170 1704.000 1570.710 1704.280 ;
        RECT 1571.550 1704.000 1572.550 1704.280 ;
        RECT 1573.390 1704.000 1573.930 1704.280 ;
        RECT 1574.770 1704.000 1575.770 1704.280 ;
        RECT 1576.610 1704.000 1577.150 1704.280 ;
        RECT 1577.990 1704.000 1578.990 1704.280 ;
        RECT 1579.830 1704.000 1580.370 1704.280 ;
        RECT 1581.210 1704.000 1582.210 1704.280 ;
        RECT 1583.050 1704.000 1583.590 1704.280 ;
        RECT 1584.430 1704.000 1585.430 1704.280 ;
        RECT 1586.270 1704.000 1586.810 1704.280 ;
        RECT 1587.650 1704.000 1588.650 1704.280 ;
        RECT 1589.490 1704.000 1590.030 1704.280 ;
        RECT 1590.870 1704.000 1591.870 1704.280 ;
        RECT 1592.710 1704.000 1593.250 1704.280 ;
        RECT 1594.090 1704.000 1595.090 1704.280 ;
        RECT 1595.930 1704.000 1596.470 1704.280 ;
        RECT 1597.310 1704.000 1598.310 1704.280 ;
        RECT 1599.150 1704.000 1599.690 1704.280 ;
        RECT 1600.530 1704.000 1601.530 1704.280 ;
        RECT 1602.370 1704.000 1602.910 1704.280 ;
        RECT 1603.750 1704.000 1604.750 1704.280 ;
        RECT 1605.590 1704.000 1606.130 1704.280 ;
        RECT 1606.970 1704.000 1607.970 1704.280 ;
        RECT 1608.810 1704.000 1609.350 1704.280 ;
        RECT 1610.190 1704.000 1611.190 1704.280 ;
        RECT 1612.030 1704.000 1612.570 1704.280 ;
        RECT 1613.410 1704.000 1614.410 1704.280 ;
        RECT 1615.250 1704.000 1615.790 1704.280 ;
        RECT 1616.630 1704.000 1617.630 1704.280 ;
        RECT 1618.470 1704.000 1619.010 1704.280 ;
        RECT 1619.850 1704.000 1620.850 1704.280 ;
        RECT 1621.690 1704.000 1622.230 1704.280 ;
        RECT 1623.070 1704.000 1624.070 1704.280 ;
        RECT 1624.910 1704.000 1625.450 1704.280 ;
        RECT 1626.290 1704.000 1627.290 1704.280 ;
        RECT 1628.130 1704.000 1628.670 1704.280 ;
        RECT 1629.510 1704.000 1630.510 1704.280 ;
        RECT 1631.350 1704.000 1631.890 1704.280 ;
        RECT 1632.730 1704.000 1633.730 1704.280 ;
        RECT 1634.570 1704.000 1635.110 1704.280 ;
        RECT 1635.950 1704.000 1636.950 1704.280 ;
        RECT 1637.790 1704.000 1638.330 1704.280 ;
        RECT 1639.170 1704.000 1640.170 1704.280 ;
        RECT 1641.010 1704.000 1641.550 1704.280 ;
        RECT 1642.390 1704.000 1643.390 1704.280 ;
        RECT 1644.230 1704.000 1644.770 1704.280 ;
        RECT 1645.610 1704.000 1646.610 1704.280 ;
        RECT 1647.450 1704.000 1647.990 1704.280 ;
        RECT 1648.830 1704.000 1649.830 1704.280 ;
        RECT 1650.670 1704.000 1651.210 1704.280 ;
        RECT 1652.050 1704.000 1652.590 1704.280 ;
        RECT 1653.430 1704.000 1654.430 1704.280 ;
        RECT 1655.270 1704.000 1655.810 1704.280 ;
        RECT 1656.650 1704.000 1657.650 1704.280 ;
        RECT 1658.490 1704.000 1659.030 1704.280 ;
        RECT 1659.870 1704.000 1660.870 1704.280 ;
        RECT 1661.710 1704.000 1662.250 1704.280 ;
        RECT 1663.090 1704.000 1664.090 1704.280 ;
        RECT 1664.930 1704.000 1665.470 1704.280 ;
        RECT 1666.310 1704.000 1667.310 1704.280 ;
        RECT 1668.150 1704.000 1668.690 1704.280 ;
        RECT 1669.530 1704.000 1670.530 1704.280 ;
        RECT 1671.370 1704.000 1671.910 1704.280 ;
        RECT 1672.750 1704.000 1673.750 1704.280 ;
        RECT 1674.590 1704.000 1675.130 1704.280 ;
        RECT 1675.970 1704.000 1676.970 1704.280 ;
        RECT 1677.810 1704.000 1678.350 1704.280 ;
        RECT 1679.190 1704.000 1680.190 1704.280 ;
        RECT 1681.030 1704.000 1681.570 1704.280 ;
        RECT 1682.410 1704.000 1683.410 1704.280 ;
        RECT 1684.250 1704.000 1684.790 1704.280 ;
        RECT 1685.630 1704.000 1686.630 1704.280 ;
        RECT 1687.470 1704.000 1688.010 1704.280 ;
        RECT 1688.850 1704.000 1689.850 1704.280 ;
        RECT 1690.690 1704.000 1691.230 1704.280 ;
        RECT 1692.070 1704.000 1693.070 1704.280 ;
        RECT 1693.910 1704.000 1694.450 1704.280 ;
        RECT 1695.290 1704.000 1696.290 1704.280 ;
        RECT 1697.130 1704.000 1697.670 1704.280 ;
        RECT 1698.510 1704.000 1699.510 1704.280 ;
        RECT 1700.350 1704.000 1700.890 1704.280 ;
        RECT 1701.730 1704.000 1702.730 1704.280 ;
        RECT 1703.570 1704.000 1704.110 1704.280 ;
        RECT 1704.950 1704.000 1705.950 1704.280 ;
        RECT 1706.790 1704.000 1707.330 1704.280 ;
        RECT 1708.170 1704.000 1709.170 1704.280 ;
        RECT 1710.010 1704.000 1710.550 1704.280 ;
        RECT 1711.390 1704.000 1712.390 1704.280 ;
        RECT 1713.230 1704.000 1713.770 1704.280 ;
        RECT 1714.610 1704.000 1715.610 1704.280 ;
        RECT 1716.450 1704.000 1716.990 1704.280 ;
        RECT 1717.830 1704.000 1718.830 1704.280 ;
        RECT 1719.670 1704.000 1720.210 1704.280 ;
        RECT 1721.050 1704.000 1722.050 1704.280 ;
        RECT 1722.890 1704.000 1723.430 1704.280 ;
        RECT 1724.270 1704.000 1725.270 1704.280 ;
        RECT 1726.110 1704.000 1726.650 1704.280 ;
        RECT 1727.490 1704.000 1728.490 1704.280 ;
        RECT 1729.330 1704.000 1729.870 1704.280 ;
        RECT 1730.710 1704.000 1731.710 1704.280 ;
        RECT 1732.550 1704.000 1733.090 1704.280 ;
        RECT 1733.930 1704.000 1734.930 1704.280 ;
        RECT 1735.770 1704.000 1736.310 1704.280 ;
        RECT 1737.150 1704.000 1738.150 1704.280 ;
        RECT 1738.990 1704.000 1739.530 1704.280 ;
        RECT 1740.370 1704.000 1741.370 1704.280 ;
        RECT 1742.210 1704.000 1742.750 1704.280 ;
        RECT 1743.590 1704.000 1744.590 1704.280 ;
        RECT 1745.430 1704.000 1745.970 1704.280 ;
        RECT 1746.810 1704.000 1747.810 1704.280 ;
        RECT 1748.650 1704.000 1749.190 1704.280 ;
        RECT 1750.030 1704.000 1750.570 1704.280 ;
        RECT 1751.410 1704.000 1752.410 1704.280 ;
        RECT 1753.250 1704.000 1753.790 1704.280 ;
        RECT 1754.630 1704.000 1755.630 1704.280 ;
        RECT 1756.470 1704.000 1757.010 1704.280 ;
        RECT 1757.850 1704.000 1758.850 1704.280 ;
        RECT 1759.690 1704.000 1760.230 1704.280 ;
        RECT 1761.070 1704.000 1762.070 1704.280 ;
        RECT 1762.910 1704.000 1763.450 1704.280 ;
        RECT 1764.290 1704.000 1765.290 1704.280 ;
        RECT 1766.130 1704.000 1766.670 1704.280 ;
        RECT 1767.510 1704.000 1768.510 1704.280 ;
        RECT 1769.350 1704.000 1769.890 1704.280 ;
        RECT 1770.730 1704.000 1771.730 1704.280 ;
        RECT 1772.570 1704.000 1773.110 1704.280 ;
        RECT 1773.950 1704.000 1774.950 1704.280 ;
        RECT 1775.790 1704.000 1776.330 1704.280 ;
        RECT 1777.170 1704.000 1778.170 1704.280 ;
        RECT 1779.010 1704.000 1779.550 1704.280 ;
        RECT 1780.390 1704.000 1781.390 1704.280 ;
        RECT 1782.230 1704.000 1782.770 1704.280 ;
        RECT 1783.610 1704.000 1784.610 1704.280 ;
        RECT 1785.450 1704.000 1785.990 1704.280 ;
        RECT 1786.830 1704.000 1787.830 1704.280 ;
        RECT 1788.670 1704.000 1789.210 1704.280 ;
        RECT 1790.050 1704.000 1791.050 1704.280 ;
        RECT 1791.890 1704.000 1792.430 1704.280 ;
        RECT 1793.270 1704.000 1794.270 1704.280 ;
        RECT 1795.110 1704.000 1795.650 1704.280 ;
        RECT 1796.490 1704.000 1797.490 1704.280 ;
        RECT 1798.330 1704.000 1798.870 1704.280 ;
        RECT 1799.710 1704.000 1800.710 1704.280 ;
        RECT 1801.550 1704.000 1802.090 1704.280 ;
        RECT 1802.930 1704.000 1803.930 1704.280 ;
        RECT 1804.770 1704.000 1805.310 1704.280 ;
        RECT 1806.150 1704.000 1807.150 1704.280 ;
        RECT 1807.990 1704.000 1808.530 1704.280 ;
        RECT 1809.370 1704.000 1810.370 1704.280 ;
        RECT 1811.210 1704.000 1811.750 1704.280 ;
        RECT 1812.590 1704.000 1813.590 1704.280 ;
        RECT 1814.430 1704.000 1814.970 1704.280 ;
        RECT 1815.810 1704.000 1816.810 1704.280 ;
        RECT 1817.650 1704.000 1818.190 1704.280 ;
        RECT 1819.030 1704.000 1820.030 1704.280 ;
        RECT 1820.870 1704.000 1821.410 1704.280 ;
        RECT 1822.250 1704.000 1823.250 1704.280 ;
        RECT 1824.090 1704.000 1824.630 1704.280 ;
        RECT 1825.470 1704.000 1826.470 1704.280 ;
        RECT 1827.310 1704.000 1827.850 1704.280 ;
        RECT 1828.690 1704.000 1829.690 1704.280 ;
        RECT 1830.530 1704.000 1831.070 1704.280 ;
        RECT 1831.910 1704.000 1832.910 1704.280 ;
        RECT 1833.750 1704.000 1834.290 1704.280 ;
        RECT 1835.130 1704.000 1836.130 1704.280 ;
        RECT 1836.970 1704.000 1837.510 1704.280 ;
        RECT 1838.350 1704.000 1839.350 1704.280 ;
        RECT 1840.190 1704.000 1840.730 1704.280 ;
        RECT 1841.570 1704.000 1842.570 1704.280 ;
        RECT 1843.410 1704.000 1843.950 1704.280 ;
        RECT 1844.790 1704.000 1845.790 1704.280 ;
        RECT 1846.630 1704.000 1847.170 1704.280 ;
        RECT 1848.010 1704.000 1849.010 1704.280 ;
        RECT 1849.850 1704.000 1850.390 1704.280 ;
        RECT 1851.230 1704.000 1851.770 1704.280 ;
        RECT 1852.610 1704.000 1853.610 1704.280 ;
        RECT 1854.450 1704.000 1854.990 1704.280 ;
        RECT 1855.830 1704.000 1856.830 1704.280 ;
        RECT 1857.670 1704.000 1858.210 1704.280 ;
        RECT 1859.050 1704.000 1860.050 1704.280 ;
        RECT 1860.890 1704.000 1861.430 1704.280 ;
        RECT 1862.270 1704.000 1863.270 1704.280 ;
        RECT 1864.110 1704.000 1864.650 1704.280 ;
        RECT 1865.490 1704.000 1866.490 1704.280 ;
        RECT 1867.330 1704.000 1867.870 1704.280 ;
        RECT 1868.710 1704.000 1869.710 1704.280 ;
        RECT 1870.550 1704.000 1871.090 1704.280 ;
        RECT 1871.930 1704.000 1872.930 1704.280 ;
        RECT 1873.770 1704.000 1874.310 1704.280 ;
        RECT 1875.150 1704.000 1876.150 1704.280 ;
        RECT 1876.990 1704.000 1877.530 1704.280 ;
        RECT 1878.370 1704.000 1879.370 1704.280 ;
        RECT 1880.210 1704.000 1880.750 1704.280 ;
        RECT 1881.590 1704.000 1882.590 1704.280 ;
        RECT 1883.430 1704.000 1883.970 1704.280 ;
        RECT 1884.810 1704.000 1885.810 1704.280 ;
        RECT 1886.650 1704.000 1887.190 1704.280 ;
        RECT 1888.030 1704.000 1889.030 1704.280 ;
        RECT 1889.870 1704.000 1890.410 1704.280 ;
        RECT 1891.250 1704.000 1892.250 1704.280 ;
        RECT 1893.090 1704.000 1893.630 1704.280 ;
        RECT 1894.470 1704.000 1895.470 1704.280 ;
        RECT 1896.310 1704.000 1896.850 1704.280 ;
        RECT 1897.690 1704.000 1898.690 1704.280 ;
        RECT 1899.530 1704.000 1900.070 1704.280 ;
        RECT 1900.910 1704.000 1901.910 1704.280 ;
        RECT 1902.750 1704.000 1903.290 1704.280 ;
        RECT 1904.130 1704.000 1905.130 1704.280 ;
        RECT 1905.970 1704.000 1906.510 1704.280 ;
        RECT 1907.350 1704.000 1908.350 1704.280 ;
        RECT 1909.190 1704.000 1909.730 1704.280 ;
        RECT 1910.570 1704.000 1911.570 1704.280 ;
        RECT 1912.410 1704.000 1912.950 1704.280 ;
        RECT 1913.790 1704.000 1914.790 1704.280 ;
        RECT 1915.630 1704.000 1916.170 1704.280 ;
        RECT 1917.010 1704.000 1918.010 1704.280 ;
        RECT 1918.850 1704.000 1919.390 1704.280 ;
        RECT 1920.230 1704.000 1921.230 1704.280 ;
        RECT 1922.070 1704.000 1922.610 1704.280 ;
        RECT 1923.450 1704.000 1924.450 1704.280 ;
        RECT 1925.290 1704.000 1925.830 1704.280 ;
        RECT 1926.670 1704.000 1927.670 1704.280 ;
        RECT 1928.510 1704.000 1929.050 1704.280 ;
        RECT 1929.890 1704.000 1930.890 1704.280 ;
        RECT 1931.730 1704.000 1932.270 1704.280 ;
        RECT 1933.110 1704.000 1934.110 1704.280 ;
        RECT 1934.950 1704.000 1935.490 1704.280 ;
        RECT 1936.330 1704.000 1937.330 1704.280 ;
        RECT 1938.170 1704.000 1938.710 1704.280 ;
        RECT 1939.550 1704.000 1940.550 1704.280 ;
        RECT 1941.390 1704.000 1941.930 1704.280 ;
        RECT 1942.770 1704.000 1943.770 1704.280 ;
        RECT 1944.610 1704.000 1945.150 1704.280 ;
        RECT 1945.990 1704.000 1946.620 1704.280 ;
      LAYER met3 ;
        RECT 1150.525 2459.920 1946.000 2488.965 ;
        RECT 1154.400 2458.520 1946.000 2459.920 ;
        RECT 1150.525 2434.080 1946.000 2458.520 ;
        RECT 1150.525 2432.680 1945.600 2434.080 ;
        RECT 1150.525 2379.680 1946.000 2432.680 ;
        RECT 1154.400 2378.280 1946.000 2379.680 ;
        RECT 1150.525 2300.800 1946.000 2378.280 ;
        RECT 1150.525 2300.120 1945.600 2300.800 ;
        RECT 1154.400 2299.400 1945.600 2300.120 ;
        RECT 1154.400 2298.720 1946.000 2299.400 ;
        RECT 1150.525 2219.880 1946.000 2298.720 ;
        RECT 1154.400 2218.480 1946.000 2219.880 ;
        RECT 1150.525 2167.520 1946.000 2218.480 ;
        RECT 1150.525 2166.120 1945.600 2167.520 ;
        RECT 1150.525 2140.320 1946.000 2166.120 ;
        RECT 1154.400 2138.920 1946.000 2140.320 ;
        RECT 1150.525 2060.080 1946.000 2138.920 ;
        RECT 1154.400 2058.680 1946.000 2060.080 ;
        RECT 1150.525 2034.240 1946.000 2058.680 ;
        RECT 1150.525 2032.840 1945.600 2034.240 ;
        RECT 1150.525 1979.840 1946.000 2032.840 ;
        RECT 1154.400 1978.440 1946.000 1979.840 ;
        RECT 1150.525 1900.960 1946.000 1978.440 ;
        RECT 1150.525 1900.280 1945.600 1900.960 ;
        RECT 1154.400 1899.560 1945.600 1900.280 ;
        RECT 1154.400 1898.880 1946.000 1899.560 ;
        RECT 1150.525 1820.040 1946.000 1898.880 ;
        RECT 1154.400 1818.640 1946.000 1820.040 ;
        RECT 1150.525 1767.680 1946.000 1818.640 ;
        RECT 1150.525 1766.280 1945.600 1767.680 ;
        RECT 1150.525 1740.480 1946.000 1766.280 ;
        RECT 1154.400 1739.080 1946.000 1740.480 ;
        RECT 1150.525 1710.715 1946.000 1739.080 ;
      LAYER met4 ;
        RECT 1171.040 1710.640 1172.640 2489.040 ;
        RECT 1247.840 1710.640 1249.440 2489.040 ;
      LAYER met4 ;
        RECT 1281.855 1710.640 1282.020 2489.040 ;
        RECT 1285.020 1710.640 1300.020 2489.040 ;
        RECT 1303.020 1710.640 1318.020 2489.040 ;
        RECT 1321.020 1710.640 1354.020 2489.040 ;
        RECT 1357.020 1710.640 1372.020 2489.040 ;
        RECT 1375.020 1710.640 1390.020 2489.040 ;
        RECT 1393.020 1710.640 1408.020 2489.040 ;
        RECT 1411.020 1710.640 1444.020 2489.040 ;
        RECT 1447.020 1710.640 1462.020 2489.040 ;
        RECT 1465.020 1710.640 1480.020 2489.040 ;
        RECT 1483.020 1710.640 1498.020 2489.040 ;
        RECT 1501.020 1710.640 1534.020 2489.040 ;
        RECT 1537.020 1710.640 1552.020 2489.040 ;
        RECT 1555.020 1710.640 1570.020 2489.040 ;
        RECT 1573.020 1710.640 1588.020 2489.040 ;
        RECT 1591.020 1710.640 1624.020 2489.040 ;
        RECT 1627.020 1710.640 1642.020 2489.040 ;
        RECT 1645.020 1710.640 1660.020 2489.040 ;
        RECT 1663.020 1710.640 1678.020 2489.040 ;
        RECT 1681.020 1710.640 1714.020 2489.040 ;
        RECT 1717.020 1710.640 1732.020 2489.040 ;
        RECT 1735.020 1710.640 1750.020 2489.040 ;
        RECT 1753.020 1710.640 1768.020 2489.040 ;
        RECT 1771.020 1710.640 1804.020 2489.040 ;
        RECT 1807.020 1710.640 1822.020 2489.040 ;
        RECT 1825.020 1710.640 1840.020 2489.040 ;
        RECT 1843.020 1710.640 1858.020 2489.040 ;
        RECT 1861.020 1710.640 1894.020 2489.040 ;
        RECT 1897.020 1710.640 1912.020 2489.040 ;
        RECT 1915.020 1710.640 1930.020 2489.040 ;
        RECT 1933.020 1710.640 1940.640 2489.040 ;
>>>>>>> Latest run - not LVS matched yet
  END
END user_project_wrapper
END LIBRARY

