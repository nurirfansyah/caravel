VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1297.270 30.840 1297.590 30.900 ;
        RECT 1386.050 30.840 1386.370 30.900 ;
        RECT 1297.270 30.700 1386.370 30.840 ;
        RECT 1297.270 30.640 1297.590 30.700 ;
        RECT 1386.050 30.640 1386.370 30.700 ;
        RECT 2801.470 29.480 2801.790 29.540 ;
        RECT 2849.310 29.480 2849.630 29.540 ;
        RECT 2801.470 29.340 2849.630 29.480 ;
        RECT 2801.470 29.280 2801.790 29.340 ;
        RECT 2849.310 29.280 2849.630 29.340 ;
        RECT 1435.730 28.460 1436.050 28.520 ;
        RECT 1454.590 28.460 1454.910 28.520 ;
        RECT 1435.730 28.320 1454.910 28.460 ;
        RECT 1435.730 28.260 1436.050 28.320 ;
        RECT 1454.590 28.260 1454.910 28.320 ;
        RECT 1653.770 28.460 1654.090 28.520 ;
        RECT 1656.990 28.460 1657.310 28.520 ;
        RECT 1653.770 28.320 1657.310 28.460 ;
        RECT 1653.770 28.260 1654.090 28.320 ;
        RECT 1656.990 28.260 1657.310 28.320 ;
        RECT 2401.270 28.460 2401.590 28.520 ;
        RECT 2415.070 28.460 2415.390 28.520 ;
        RECT 2401.270 28.320 2415.390 28.460 ;
        RECT 2401.270 28.260 2401.590 28.320 ;
        RECT 2415.070 28.260 2415.390 28.320 ;
        RECT 2553.070 28.460 2553.390 28.520 ;
        RECT 2600.910 28.460 2601.230 28.520 ;
        RECT 2553.070 28.320 2601.230 28.460 ;
        RECT 2553.070 28.260 2553.390 28.320 ;
        RECT 2600.910 28.260 2601.230 28.320 ;
        RECT 2705.330 28.460 2705.650 28.520 ;
        RECT 2752.710 28.460 2753.030 28.520 ;
        RECT 2705.330 28.320 2753.030 28.460 ;
        RECT 2705.330 28.260 2705.650 28.320 ;
        RECT 2752.710 28.260 2753.030 28.320 ;
      LAYER via ;
        RECT 1297.300 30.640 1297.560 30.900 ;
        RECT 1386.080 30.640 1386.340 30.900 ;
        RECT 2801.500 29.280 2801.760 29.540 ;
        RECT 2849.340 29.280 2849.600 29.540 ;
        RECT 1435.760 28.260 1436.020 28.520 ;
        RECT 1454.620 28.260 1454.880 28.520 ;
        RECT 1653.800 28.260 1654.060 28.520 ;
        RECT 1657.020 28.260 1657.280 28.520 ;
        RECT 2401.300 28.260 2401.560 28.520 ;
        RECT 2415.100 28.260 2415.360 28.520 ;
        RECT 2553.100 28.260 2553.360 28.520 ;
        RECT 2600.940 28.260 2601.200 28.520 ;
        RECT 2705.360 28.260 2705.620 28.520 ;
        RECT 2752.740 28.260 2753.000 28.520 ;
      LAYER met2 ;
        RECT 1138.130 1744.355 1138.410 1744.725 ;
        RECT 1138.200 29.765 1138.340 1744.355 ;
        RECT 1248.530 30.755 1248.810 31.125 ;
        RECT 1248.600 30.445 1248.740 30.755 ;
        RECT 1297.300 30.610 1297.560 30.930 ;
        RECT 1386.080 30.610 1386.340 30.930 ;
        RECT 1201.150 30.075 1201.430 30.445 ;
        RECT 1248.530 30.075 1248.810 30.445 ;
        RECT 1138.130 29.395 1138.410 29.765 ;
        RECT 1200.690 29.395 1200.970 29.765 ;
        RECT 1200.760 28.970 1200.900 29.395 ;
        RECT 1201.220 28.970 1201.360 30.075 ;
        RECT 1297.360 29.085 1297.500 30.610 ;
        RECT 1200.760 28.830 1201.360 28.970 ;
        RECT 1297.290 28.715 1297.570 29.085 ;
        RECT 1386.140 28.405 1386.280 30.610 ;
        RECT 1617.450 30.075 1617.730 30.445 ;
        RECT 1683.690 30.075 1683.970 30.445 ;
        RECT 2070.090 30.075 2070.370 30.445 ;
        RECT 2117.930 30.075 2118.210 30.445 ;
        RECT 1386.070 28.035 1386.350 28.405 ;
        RECT 1435.290 28.290 1435.570 28.405 ;
        RECT 1435.760 28.290 1436.020 28.550 ;
        RECT 1454.620 28.405 1454.880 28.550 ;
        RECT 1617.520 28.405 1617.660 30.075 ;
        RECT 1683.760 29.085 1683.900 30.075 ;
        RECT 1657.010 28.715 1657.290 29.085 ;
        RECT 1683.690 28.715 1683.970 29.085 ;
        RECT 1973.030 28.715 1973.310 29.085 ;
        RECT 2021.330 28.715 2021.610 29.085 ;
        RECT 1657.080 28.550 1657.220 28.715 ;
        RECT 1653.800 28.405 1654.060 28.550 ;
        RECT 1435.290 28.230 1436.020 28.290 ;
        RECT 1435.290 28.150 1435.960 28.230 ;
        RECT 1435.290 28.035 1435.570 28.150 ;
        RECT 1454.610 28.035 1454.890 28.405 ;
        RECT 1617.450 28.035 1617.730 28.405 ;
        RECT 1653.790 28.035 1654.070 28.405 ;
        RECT 1657.020 28.230 1657.280 28.550 ;
        RECT 1852.510 28.035 1852.790 28.405 ;
        RECT 1852.580 25.685 1852.720 28.035 ;
        RECT 1973.100 27.045 1973.240 28.715 ;
        RECT 2021.400 27.725 2021.540 28.715 ;
        RECT 2070.160 28.405 2070.300 30.075 ;
        RECT 2118.000 29.085 2118.140 30.075 ;
        RECT 2801.490 29.395 2801.770 29.765 ;
        RECT 2801.500 29.250 2801.760 29.395 ;
        RECT 2849.340 29.250 2849.600 29.570 ;
        RECT 2117.930 28.715 2118.210 29.085 ;
        RECT 2138.630 28.970 2138.910 29.085 ;
        RECT 2187.850 28.970 2188.130 29.085 ;
        RECT 2284.450 28.970 2284.730 29.085 ;
        RECT 2138.630 28.830 2139.760 28.970 ;
        RECT 2138.630 28.715 2138.910 28.830 ;
        RECT 2139.620 28.405 2139.760 28.830 ;
        RECT 2187.000 28.830 2188.130 28.970 ;
        RECT 2187.000 28.405 2187.140 28.830 ;
        RECT 2187.850 28.715 2188.130 28.830 ;
        RECT 2283.600 28.830 2284.730 28.970 ;
        RECT 2283.600 28.405 2283.740 28.830 ;
        RECT 2284.450 28.715 2284.730 28.830 ;
        RECT 2304.690 28.715 2304.970 29.085 ;
        RECT 2600.930 28.715 2601.210 29.085 ;
        RECT 2304.760 28.405 2304.900 28.715 ;
        RECT 2601.000 28.550 2601.140 28.715 ;
        RECT 2401.300 28.405 2401.560 28.550 ;
        RECT 2415.100 28.405 2415.360 28.550 ;
        RECT 2553.100 28.405 2553.360 28.550 ;
        RECT 2070.090 28.035 2070.370 28.405 ;
        RECT 2139.550 28.035 2139.830 28.405 ;
        RECT 2186.930 28.035 2187.210 28.405 ;
        RECT 2283.530 28.035 2283.810 28.405 ;
        RECT 2304.690 28.035 2304.970 28.405 ;
        RECT 2401.290 28.035 2401.570 28.405 ;
        RECT 2415.090 28.035 2415.370 28.405 ;
        RECT 2528.710 28.035 2528.990 28.405 ;
        RECT 2553.090 28.035 2553.370 28.405 ;
        RECT 2600.940 28.230 2601.200 28.550 ;
        RECT 2705.360 28.405 2705.620 28.550 ;
        RECT 2752.740 28.405 2753.000 28.550 ;
        RECT 2849.400 28.405 2849.540 29.250 ;
        RECT 2680.510 28.035 2680.790 28.405 ;
        RECT 2705.350 28.035 2705.630 28.405 ;
        RECT 2752.730 28.035 2753.010 28.405 ;
        RECT 2849.330 28.035 2849.610 28.405 ;
        RECT 2021.330 27.355 2021.610 27.725 ;
        RECT 1973.030 26.675 1973.310 27.045 ;
        RECT 2528.780 26.365 2528.920 28.035 ;
        RECT 2680.580 27.045 2680.720 28.035 ;
        RECT 2680.510 26.675 2680.790 27.045 ;
        RECT 2528.710 25.995 2528.990 26.365 ;
        RECT 1852.510 25.315 1852.790 25.685 ;
      LAYER via2 ;
        RECT 1138.130 1744.400 1138.410 1744.680 ;
        RECT 1248.530 30.800 1248.810 31.080 ;
        RECT 1201.150 30.120 1201.430 30.400 ;
        RECT 1248.530 30.120 1248.810 30.400 ;
        RECT 1138.130 29.440 1138.410 29.720 ;
        RECT 1200.690 29.440 1200.970 29.720 ;
        RECT 1297.290 28.760 1297.570 29.040 ;
        RECT 1617.450 30.120 1617.730 30.400 ;
        RECT 1683.690 30.120 1683.970 30.400 ;
        RECT 2070.090 30.120 2070.370 30.400 ;
        RECT 2117.930 30.120 2118.210 30.400 ;
        RECT 1386.070 28.080 1386.350 28.360 ;
        RECT 1435.290 28.080 1435.570 28.360 ;
        RECT 1657.010 28.760 1657.290 29.040 ;
        RECT 1683.690 28.760 1683.970 29.040 ;
        RECT 1973.030 28.760 1973.310 29.040 ;
        RECT 2021.330 28.760 2021.610 29.040 ;
        RECT 1454.610 28.080 1454.890 28.360 ;
        RECT 1617.450 28.080 1617.730 28.360 ;
        RECT 1653.790 28.080 1654.070 28.360 ;
        RECT 1852.510 28.080 1852.790 28.360 ;
        RECT 2801.490 29.440 2801.770 29.720 ;
        RECT 2117.930 28.760 2118.210 29.040 ;
        RECT 2138.630 28.760 2138.910 29.040 ;
        RECT 2187.850 28.760 2188.130 29.040 ;
        RECT 2284.450 28.760 2284.730 29.040 ;
        RECT 2304.690 28.760 2304.970 29.040 ;
        RECT 2600.930 28.760 2601.210 29.040 ;
        RECT 2070.090 28.080 2070.370 28.360 ;
        RECT 2139.550 28.080 2139.830 28.360 ;
        RECT 2186.930 28.080 2187.210 28.360 ;
        RECT 2283.530 28.080 2283.810 28.360 ;
        RECT 2304.690 28.080 2304.970 28.360 ;
        RECT 2401.290 28.080 2401.570 28.360 ;
        RECT 2415.090 28.080 2415.370 28.360 ;
        RECT 2528.710 28.080 2528.990 28.360 ;
        RECT 2553.090 28.080 2553.370 28.360 ;
        RECT 2680.510 28.080 2680.790 28.360 ;
        RECT 2705.350 28.080 2705.630 28.360 ;
        RECT 2752.730 28.080 2753.010 28.360 ;
        RECT 2849.330 28.080 2849.610 28.360 ;
        RECT 2021.330 27.400 2021.610 27.680 ;
        RECT 1973.030 26.720 1973.310 27.000 ;
        RECT 2680.510 26.720 2680.790 27.000 ;
        RECT 2528.710 26.040 2528.990 26.320 ;
        RECT 1852.510 25.360 1852.790 25.640 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 28.980 2924.800 30.180 ;
=======
        RECT 2900.825 29.730 2901.155 29.745 ;
=======
        RECT 1138.105 1744.690 1138.435 1744.705 ;
        RECT 1150.000 1744.690 1154.000 1744.840 ;
        RECT 1138.105 1744.390 1154.000 1744.690 ;
        RECT 1138.105 1744.375 1138.435 1744.390 ;
        RECT 1150.000 1744.240 1154.000 1744.390 ;
        RECT 1248.505 31.100 1248.835 31.105 ;
        RECT 1248.505 31.090 1249.090 31.100 ;
        RECT 1248.300 30.790 1249.090 31.090 ;
        RECT 1248.505 30.780 1249.090 30.790 ;
        RECT 1248.505 30.775 1248.835 30.780 ;
        RECT 1201.125 30.410 1201.455 30.425 ;
        RECT 1248.505 30.410 1248.835 30.425 ;
        RECT 1617.425 30.410 1617.755 30.425 ;
        RECT 1201.125 30.110 1248.835 30.410 ;
        RECT 1201.125 30.095 1201.455 30.110 ;
        RECT 1248.505 30.095 1248.835 30.110 ;
        RECT 1593.750 30.110 1617.755 30.410 ;
        RECT 1138.105 29.730 1138.435 29.745 ;
        RECT 1200.665 29.730 1200.995 29.745 ;
        RECT 1138.105 29.430 1200.995 29.730 ;
        RECT 1138.105 29.415 1138.435 29.430 ;
        RECT 1200.665 29.415 1200.995 29.430 ;
        RECT 1497.110 29.730 1497.490 29.740 ;
        RECT 1538.510 29.730 1538.890 29.740 ;
        RECT 1497.110 29.430 1538.890 29.730 ;
        RECT 1497.110 29.420 1497.490 29.430 ;
        RECT 1538.510 29.420 1538.890 29.430 ;
        RECT 1248.710 29.050 1249.090 29.060 ;
        RECT 1297.265 29.050 1297.595 29.065 ;
        RECT 1248.710 28.750 1297.595 29.050 ;
        RECT 1248.710 28.740 1249.090 28.750 ;
        RECT 1297.265 28.735 1297.595 28.750 ;
        RECT 1586.350 29.050 1586.730 29.060 ;
        RECT 1593.750 29.050 1594.050 30.110 ;
        RECT 1617.425 30.095 1617.755 30.110 ;
        RECT 1683.665 30.410 1683.995 30.425 ;
        RECT 1730.790 30.410 1731.170 30.420 ;
        RECT 1683.665 30.110 1731.170 30.410 ;
        RECT 1683.665 30.095 1683.995 30.110 ;
        RECT 1730.790 30.100 1731.170 30.110 ;
        RECT 2070.065 30.410 2070.395 30.425 ;
        RECT 2117.905 30.410 2118.235 30.425 ;
        RECT 2070.065 30.110 2118.235 30.410 ;
        RECT 2070.065 30.095 2070.395 30.110 ;
        RECT 2117.905 30.095 2118.235 30.110 ;
        RECT 2801.465 29.730 2801.795 29.745 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 29.730 2924.800 30.180 ;
        RECT 2766.750 29.430 2801.795 29.730 ;
        RECT 1586.350 28.750 1594.050 29.050 ;
        RECT 1656.985 29.050 1657.315 29.065 ;
        RECT 1683.665 29.050 1683.995 29.065 ;
        RECT 1656.985 28.750 1683.995 29.050 ;
        RECT 1586.350 28.740 1586.730 28.750 ;
        RECT 1656.985 28.735 1657.315 28.750 ;
        RECT 1683.665 28.735 1683.995 28.750 ;
        RECT 1751.990 29.050 1753.210 29.220 ;
        RECT 1786.910 29.050 1787.290 29.060 ;
        RECT 1973.005 29.050 1973.335 29.065 ;
        RECT 2021.305 29.050 2021.635 29.065 ;
        RECT 2117.905 29.050 2118.235 29.065 ;
        RECT 2138.605 29.050 2138.935 29.065 ;
        RECT 1751.990 28.920 1787.290 29.050 ;
        RECT 1386.045 28.370 1386.375 28.385 ;
        RECT 1435.265 28.370 1435.595 28.385 ;
        RECT 1386.045 28.070 1435.595 28.370 ;
        RECT 1386.045 28.055 1386.375 28.070 ;
        RECT 1435.265 28.055 1435.595 28.070 ;
        RECT 1454.585 28.370 1454.915 28.385 ;
        RECT 1617.425 28.370 1617.755 28.385 ;
        RECT 1653.765 28.370 1654.095 28.385 ;
        RECT 1454.585 28.070 1497.450 28.370 ;
        RECT 1454.585 28.055 1454.915 28.070 ;
        RECT 1497.150 27.700 1497.450 28.070 ;
        RECT 1617.425 28.070 1654.095 28.370 ;
        RECT 1617.425 28.055 1617.755 28.070 ;
        RECT 1653.765 28.055 1654.095 28.070 ;
        RECT 1730.790 28.370 1731.170 28.380 ;
        RECT 1751.990 28.370 1752.290 28.920 ;
        RECT 1752.910 28.750 1787.290 28.920 ;
        RECT 1786.910 28.740 1787.290 28.750 ;
        RECT 1876.190 28.750 1907.770 29.050 ;
        RECT 1730.790 28.070 1752.290 28.370 ;
        RECT 1852.485 28.370 1852.815 28.385 ;
        RECT 1876.190 28.370 1876.490 28.750 ;
        RECT 1852.485 28.070 1876.490 28.370 ;
        RECT 1907.470 28.370 1907.770 28.750 ;
        RECT 1973.005 28.750 1974.010 29.050 ;
        RECT 1973.005 28.735 1973.335 28.750 ;
        RECT 1924.910 28.370 1925.290 28.380 ;
        RECT 1907.470 28.070 1925.290 28.370 ;
        RECT 1730.790 28.060 1731.170 28.070 ;
        RECT 1852.485 28.055 1852.815 28.070 ;
        RECT 1924.910 28.060 1925.290 28.070 ;
        RECT 1497.110 27.380 1497.490 27.700 ;
        RECT 1538.510 27.690 1538.890 27.700 ;
        RECT 1586.350 27.690 1586.730 27.700 ;
        RECT 1538.510 27.390 1586.730 27.690 ;
        RECT 1973.710 27.690 1974.010 28.750 ;
        RECT 2021.305 28.750 2028.290 29.050 ;
        RECT 2021.305 28.735 2021.635 28.750 ;
        RECT 2027.990 28.370 2028.290 28.750 ;
        RECT 2117.905 28.750 2138.935 29.050 ;
        RECT 2117.905 28.735 2118.235 28.750 ;
        RECT 2138.605 28.735 2138.935 28.750 ;
        RECT 2187.825 29.050 2188.155 29.065 ;
        RECT 2284.425 29.050 2284.755 29.065 ;
        RECT 2304.665 29.050 2304.995 29.065 ;
        RECT 2187.825 28.750 2235.290 29.050 ;
        RECT 2187.825 28.735 2188.155 28.750 ;
        RECT 2070.065 28.370 2070.395 28.385 ;
        RECT 2027.990 28.070 2070.395 28.370 ;
        RECT 2070.065 28.055 2070.395 28.070 ;
        RECT 2139.525 28.370 2139.855 28.385 ;
        RECT 2186.905 28.370 2187.235 28.385 ;
        RECT 2139.525 28.070 2187.235 28.370 ;
        RECT 2234.990 28.370 2235.290 28.750 ;
        RECT 2284.425 28.750 2304.995 29.050 ;
        RECT 2284.425 28.735 2284.755 28.750 ;
        RECT 2304.665 28.735 2304.995 28.750 ;
        RECT 2600.905 29.050 2601.235 29.065 ;
        RECT 2600.905 28.750 2621.690 29.050 ;
        RECT 2600.905 28.735 2601.235 28.750 ;
        RECT 2283.505 28.370 2283.835 28.385 ;
        RECT 2234.990 28.070 2283.835 28.370 ;
        RECT 2139.525 28.055 2139.855 28.070 ;
        RECT 2186.905 28.055 2187.235 28.070 ;
        RECT 2283.505 28.055 2283.835 28.070 ;
        RECT 2304.665 28.370 2304.995 28.385 ;
        RECT 2401.265 28.370 2401.595 28.385 ;
        RECT 2304.665 28.070 2401.595 28.370 ;
        RECT 2304.665 28.055 2304.995 28.070 ;
        RECT 2401.265 28.055 2401.595 28.070 ;
        RECT 2415.065 28.370 2415.395 28.385 ;
        RECT 2528.685 28.370 2529.015 28.385 ;
        RECT 2553.065 28.370 2553.395 28.385 ;
        RECT 2415.065 28.070 2487.370 28.370 ;
        RECT 2415.065 28.055 2415.395 28.070 ;
        RECT 2021.305 27.690 2021.635 27.705 ;
        RECT 1973.710 27.390 2021.635 27.690 ;
        RECT 2487.070 27.690 2487.370 28.070 ;
        RECT 2528.685 28.070 2553.395 28.370 ;
        RECT 2621.390 28.370 2621.690 28.750 ;
        RECT 2704.190 28.750 2705.410 29.050 ;
        RECT 2656.310 28.370 2656.690 28.380 ;
        RECT 2621.390 28.070 2656.690 28.370 ;
        RECT 2528.685 28.055 2529.015 28.070 ;
        RECT 2553.065 28.055 2553.395 28.070 ;
        RECT 2656.310 28.060 2656.690 28.070 ;
        RECT 2680.485 28.370 2680.815 28.385 ;
        RECT 2704.190 28.370 2704.490 28.750 ;
        RECT 2680.485 28.070 2704.490 28.370 ;
        RECT 2705.110 28.385 2705.410 28.750 ;
        RECT 2705.110 28.070 2705.655 28.385 ;
        RECT 2680.485 28.055 2680.815 28.070 ;
        RECT 2705.325 28.055 2705.655 28.070 ;
        RECT 2752.705 28.370 2753.035 28.385 ;
        RECT 2766.750 28.370 2767.050 29.430 ;
        RECT 2801.465 29.415 2801.795 29.430 ;
        RECT 2916.710 29.430 2924.800 29.730 ;
        RECT 2916.710 29.050 2917.010 29.430 ;
        RECT 2884.510 28.750 2917.010 29.050 ;
        RECT 2917.600 28.980 2924.800 29.430 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2752.705 28.070 2767.050 28.370 ;
        RECT 2849.305 28.370 2849.635 28.385 ;
        RECT 2884.510 28.370 2884.810 28.750 ;
        RECT 2849.305 28.070 2884.810 28.370 ;
        RECT 2752.705 28.055 2753.035 28.070 ;
        RECT 2849.305 28.055 2849.635 28.070 ;
        RECT 2504.510 27.690 2504.890 27.700 ;
        RECT 2487.070 27.390 2504.890 27.690 ;
        RECT 1538.510 27.380 1538.890 27.390 ;
        RECT 1586.350 27.380 1586.730 27.390 ;
        RECT 2021.305 27.375 2021.635 27.390 ;
        RECT 2504.510 27.380 2504.890 27.390 ;
        RECT 1786.910 27.010 1787.290 27.020 ;
        RECT 1828.310 27.010 1828.690 27.020 ;
        RECT 1786.910 26.710 1828.690 27.010 ;
        RECT 1786.910 26.700 1787.290 26.710 ;
        RECT 1828.310 26.700 1828.690 26.710 ;
        RECT 1924.910 27.010 1925.290 27.020 ;
        RECT 1973.005 27.010 1973.335 27.025 ;
        RECT 1924.910 26.710 1973.335 27.010 ;
        RECT 1924.910 26.700 1925.290 26.710 ;
        RECT 1973.005 26.695 1973.335 26.710 ;
        RECT 2656.310 27.010 2656.690 27.020 ;
        RECT 2680.485 27.010 2680.815 27.025 ;
        RECT 2656.310 26.710 2680.815 27.010 ;
        RECT 2656.310 26.700 2656.690 26.710 ;
        RECT 2680.485 26.695 2680.815 26.710 ;
        RECT 2504.510 26.330 2504.890 26.340 ;
        RECT 2528.685 26.330 2529.015 26.345 ;
        RECT 2504.510 26.030 2529.015 26.330 ;
        RECT 2504.510 26.020 2504.890 26.030 ;
        RECT 2528.685 26.015 2529.015 26.030 ;
        RECT 1828.310 25.650 1828.690 25.660 ;
        RECT 1852.485 25.650 1852.815 25.665 ;
        RECT 1828.310 25.350 1852.815 25.650 ;
        RECT 1828.310 25.340 1828.690 25.350 ;
        RECT 1852.485 25.335 1852.815 25.350 ;
      LAYER via3 ;
        RECT 1248.740 30.780 1249.060 31.100 ;
        RECT 1497.140 29.420 1497.460 29.740 ;
        RECT 1538.540 29.420 1538.860 29.740 ;
        RECT 1248.740 28.740 1249.060 29.060 ;
        RECT 1586.380 28.740 1586.700 29.060 ;
        RECT 1730.820 30.100 1731.140 30.420 ;
        RECT 1730.820 28.060 1731.140 28.380 ;
        RECT 1786.940 28.740 1787.260 29.060 ;
        RECT 1924.940 28.060 1925.260 28.380 ;
        RECT 1497.140 27.380 1497.460 27.700 ;
        RECT 1538.540 27.380 1538.860 27.700 ;
        RECT 1586.380 27.380 1586.700 27.700 ;
        RECT 2656.340 28.060 2656.660 28.380 ;
        RECT 2504.540 27.380 2504.860 27.700 ;
        RECT 1786.940 26.700 1787.260 27.020 ;
        RECT 1828.340 26.700 1828.660 27.020 ;
        RECT 1924.940 26.700 1925.260 27.020 ;
        RECT 2656.340 26.700 2656.660 27.020 ;
        RECT 2504.540 26.020 2504.860 26.340 ;
        RECT 1828.340 25.340 1828.660 25.660 ;
      LAYER met4 ;
        RECT 1248.735 30.775 1249.065 31.105 ;
        RECT 1248.750 29.065 1249.050 30.775 ;
        RECT 1730.815 30.095 1731.145 30.425 ;
        RECT 1497.135 29.415 1497.465 29.745 ;
        RECT 1538.535 29.415 1538.865 29.745 ;
        RECT 1248.735 28.735 1249.065 29.065 ;
        RECT 1497.150 27.705 1497.450 29.415 ;
        RECT 1538.550 27.705 1538.850 29.415 ;
        RECT 1586.375 28.735 1586.705 29.065 ;
        RECT 1586.390 27.705 1586.690 28.735 ;
        RECT 1730.830 28.385 1731.130 30.095 ;
        RECT 1786.935 28.735 1787.265 29.065 ;
        RECT 1730.815 28.055 1731.145 28.385 ;
        RECT 1497.135 27.375 1497.465 27.705 ;
        RECT 1538.535 27.375 1538.865 27.705 ;
        RECT 1586.375 27.375 1586.705 27.705 ;
        RECT 1786.950 27.025 1787.250 28.735 ;
        RECT 1924.935 28.055 1925.265 28.385 ;
        RECT 2656.335 28.055 2656.665 28.385 ;
        RECT 1924.950 27.025 1925.250 28.055 ;
        RECT 2504.535 27.375 2504.865 27.705 ;
        RECT 1786.935 26.695 1787.265 27.025 ;
        RECT 1828.335 26.695 1828.665 27.025 ;
        RECT 1924.935 26.695 1925.265 27.025 ;
        RECT 1828.350 25.665 1828.650 26.695 ;
        RECT 2504.550 26.345 2504.850 27.375 ;
        RECT 2656.350 27.025 2656.650 28.055 ;
        RECT 2656.335 26.695 2656.665 27.025 ;
        RECT 2504.535 26.015 2504.865 26.345 ;
        RECT 1828.335 25.335 1828.665 25.665 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1963.350 2373.780 1963.670 2373.840 ;
        RECT 2899.450 2373.780 2899.770 2373.840 ;
        RECT 1963.350 2373.640 2899.770 2373.780 ;
        RECT 1963.350 2373.580 1963.670 2373.640 ;
        RECT 2899.450 2373.580 2899.770 2373.640 ;
      LAYER via ;
        RECT 1963.380 2373.580 1963.640 2373.840 ;
        RECT 2899.480 2373.580 2899.740 2373.840 ;
      LAYER met2 ;
        RECT 2899.470 2375.395 2899.750 2375.765 ;
        RECT 2899.540 2373.870 2899.680 2375.395 ;
        RECT 1963.380 2373.550 1963.640 2373.870 ;
        RECT 2899.480 2373.550 2899.740 2373.870 ;
        RECT 1963.440 2033.725 1963.580 2373.550 ;
        RECT 1963.370 2033.355 1963.650 2033.725 ;
      LAYER via2 ;
        RECT 2899.470 2375.440 2899.750 2375.720 ;
        RECT 1963.370 2033.400 1963.650 2033.680 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 2374.980 2924.800 2376.180 ;
=======
        RECT 2901.745 2375.730 2902.075 2375.745 ;
=======
        RECT 2899.445 2375.730 2899.775 2375.745 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 2375.730 2924.800 2376.180 ;
        RECT 2899.445 2375.430 2924.800 2375.730 ;
        RECT 2899.445 2375.415 2899.775 2375.430 ;
        RECT 2917.600 2374.980 2924.800 2375.430 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1946.000 2033.690 1950.000 2033.840 ;
        RECT 1963.345 2033.690 1963.675 2033.705 ;
        RECT 1946.000 2033.390 1963.675 2033.690 ;
        RECT 1946.000 2033.240 1950.000 2033.390 ;
        RECT 1963.345 2033.375 1963.675 2033.390 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2147.425 2608.225 2148.515 2608.395 ;
        RECT 2230.225 2608.225 2231.315 2608.395 ;
        RECT 2796.025 2608.225 2797.115 2608.395 ;
      LAYER mcon ;
        RECT 2148.345 2608.225 2148.515 2608.395 ;
        RECT 2231.145 2608.225 2231.315 2608.395 ;
        RECT 2796.945 2608.225 2797.115 2608.395 ;
      LAYER met1 ;
        RECT 1904.010 2608.380 1904.330 2608.440 ;
        RECT 2147.365 2608.380 2147.655 2608.425 ;
        RECT 1904.010 2608.240 2147.655 2608.380 ;
        RECT 1904.010 2608.180 1904.330 2608.240 ;
        RECT 2147.365 2608.195 2147.655 2608.240 ;
        RECT 2148.285 2608.380 2148.575 2608.425 ;
        RECT 2230.165 2608.380 2230.455 2608.425 ;
        RECT 2148.285 2608.240 2230.455 2608.380 ;
        RECT 2148.285 2608.195 2148.575 2608.240 ;
        RECT 2230.165 2608.195 2230.455 2608.240 ;
        RECT 2231.085 2608.380 2231.375 2608.425 ;
        RECT 2795.965 2608.380 2796.255 2608.425 ;
        RECT 2231.085 2608.240 2796.255 2608.380 ;
        RECT 2231.085 2608.195 2231.375 2608.240 ;
        RECT 2795.965 2608.195 2796.255 2608.240 ;
        RECT 2796.885 2608.380 2797.175 2608.425 ;
        RECT 2899.450 2608.380 2899.770 2608.440 ;
        RECT 2796.885 2608.240 2899.770 2608.380 ;
        RECT 2796.885 2608.195 2797.175 2608.240 ;
        RECT 2899.450 2608.180 2899.770 2608.240 ;
      LAYER via ;
        RECT 1904.040 2608.180 1904.300 2608.440 ;
        RECT 2899.480 2608.180 2899.740 2608.440 ;
      LAYER met2 ;
        RECT 2899.470 2609.995 2899.750 2610.365 ;
        RECT 2899.540 2608.470 2899.680 2609.995 ;
        RECT 1904.040 2608.150 1904.300 2608.470 ;
        RECT 2899.480 2608.150 2899.740 2608.470 ;
        RECT 1904.100 2500.090 1904.240 2608.150 ;
        RECT 1901.270 2499.410 1901.550 2500.000 ;
        RECT 1903.180 2499.950 1904.240 2500.090 ;
        RECT 1903.180 2499.410 1903.320 2499.950 ;
        RECT 1901.270 2499.270 1903.320 2499.410 ;
        RECT 1901.270 2496.000 1901.550 2499.270 ;
      LAYER via2 ;
        RECT 2899.470 2610.040 2899.750 2610.320 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 2609.580 2924.800 2610.780 ;
=======
        RECT 2900.825 2610.330 2901.155 2610.345 ;
=======
        RECT 2899.445 2610.330 2899.775 2610.345 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 2610.330 2924.800 2610.780 ;
        RECT 2899.445 2610.030 2924.800 2610.330 ;
        RECT 2899.445 2610.015 2899.775 2610.030 ;
        RECT 2917.600 2609.580 2924.800 2610.030 ;
<<<<<<< HEAD
        RECT 1946.000 1900.410 1950.000 1900.560 ;
        RECT 1963.345 1900.410 1963.675 1900.425 ;
        RECT 1946.000 1900.110 1963.675 1900.410 ;
        RECT 1946.000 1899.960 1950.000 1900.110 ;
        RECT 1963.345 1900.095 1963.675 1900.110 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1910.910 2842.980 1911.230 2843.040 ;
        RECT 2899.450 2842.980 2899.770 2843.040 ;
        RECT 1910.910 2842.840 2899.770 2842.980 ;
        RECT 1910.910 2842.780 1911.230 2842.840 ;
        RECT 2899.450 2842.780 2899.770 2842.840 ;
      LAYER via ;
        RECT 1910.940 2842.780 1911.200 2843.040 ;
        RECT 2899.480 2842.780 2899.740 2843.040 ;
      LAYER met2 ;
        RECT 2899.470 2844.595 2899.750 2844.965 ;
        RECT 2899.540 2843.070 2899.680 2844.595 ;
        RECT 1910.940 2842.750 1911.200 2843.070 ;
        RECT 2899.480 2842.750 2899.740 2843.070 ;
        RECT 1911.000 2500.090 1911.140 2842.750 ;
        RECT 1907.710 2499.410 1907.990 2500.000 ;
        RECT 1909.620 2499.950 1911.140 2500.090 ;
        RECT 1909.620 2499.410 1909.760 2499.950 ;
        RECT 1907.710 2499.270 1909.760 2499.410 ;
        RECT 1907.710 2496.000 1907.990 2499.270 ;
      LAYER via2 ;
        RECT 2899.470 2844.640 2899.750 2844.920 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 2844.180 2924.800 2845.380 ;
=======
        RECT 2900.825 2844.930 2901.155 2844.945 ;
=======
        RECT 2899.445 2844.930 2899.775 2844.945 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 2844.930 2924.800 2845.380 ;
        RECT 2899.445 2844.630 2924.800 2844.930 ;
        RECT 2899.445 2844.615 2899.775 2844.630 ;
        RECT 2917.600 2844.180 2924.800 2844.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1962.890 3077.580 1963.210 3077.640 ;
        RECT 2899.450 3077.580 2899.770 3077.640 ;
        RECT 1962.890 3077.440 2899.770 3077.580 ;
        RECT 1962.890 3077.380 1963.210 3077.440 ;
        RECT 2899.450 3077.380 2899.770 3077.440 ;
      LAYER via ;
        RECT 1962.920 3077.380 1963.180 3077.640 ;
        RECT 2899.480 3077.380 2899.740 3077.640 ;
      LAYER met2 ;
        RECT 2899.470 3079.195 2899.750 3079.565 ;
        RECT 2899.540 3077.670 2899.680 3079.195 ;
        RECT 1962.920 3077.350 1963.180 3077.670 ;
        RECT 2899.480 3077.350 2899.740 3077.670 ;
        RECT 1962.980 2167.005 1963.120 3077.350 ;
        RECT 1962.910 2166.635 1963.190 2167.005 ;
      LAYER via2 ;
        RECT 2899.470 3079.240 2899.750 3079.520 ;
        RECT 1962.910 2166.680 1963.190 2166.960 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 3078.780 2924.800 3079.980 ;
=======
        RECT 1943.310 3079.530 1943.690 3079.540 ;
        RECT 2028.665 3079.530 2028.995 3079.545 ;
        RECT 1943.310 3079.230 1966.650 3079.530 ;
        RECT 1943.310 3079.220 1943.690 3079.230 ;
        RECT 1966.350 3078.850 1966.650 3079.230 ;
        RECT 2015.110 3079.230 2028.995 3079.530 ;
        RECT 1966.350 3078.550 2014.490 3078.850 ;
        RECT 2014.190 3078.170 2014.490 3078.550 ;
        RECT 2015.110 3078.170 2015.410 3079.230 ;
        RECT 2028.665 3079.215 2028.995 3079.230 ;
        RECT 2207.605 3079.530 2207.935 3079.545 ;
        RECT 2669.905 3079.530 2670.235 3079.545 ;
        RECT 2207.605 3079.230 2256.450 3079.530 ;
        RECT 2207.605 3079.215 2207.935 3079.230 ;
        RECT 2090.305 3078.850 2090.635 3078.865 ;
        RECT 2173.310 3078.850 2173.690 3078.860 ;
        RECT 2076.750 3078.550 2090.635 3078.850 ;
        RECT 2014.190 3077.870 2015.410 3078.170 ;
        RECT 2042.925 3078.170 2043.255 3078.185 ;
        RECT 2076.750 3078.170 2077.050 3078.550 ;
        RECT 2090.305 3078.535 2090.635 3078.550 ;
        RECT 2139.310 3078.550 2173.690 3078.850 ;
        RECT 2256.150 3078.850 2256.450 3079.230 ;
        RECT 2304.910 3079.230 2353.050 3079.530 ;
        RECT 2256.150 3078.550 2304.290 3078.850 ;
        RECT 2042.925 3077.870 2077.050 3078.170 ;
        RECT 2090.765 3078.170 2091.095 3078.185 ;
        RECT 2139.310 3078.170 2139.610 3078.550 ;
        RECT 2173.310 3078.540 2173.690 3078.550 ;
        RECT 2090.765 3077.870 2139.610 3078.170 ;
        RECT 2303.990 3078.170 2304.290 3078.550 ;
        RECT 2304.910 3078.170 2305.210 3079.230 ;
        RECT 2352.750 3078.850 2353.050 3079.230 ;
        RECT 2401.510 3079.230 2449.650 3079.530 ;
        RECT 2352.750 3078.550 2400.890 3078.850 ;
        RECT 2303.990 3077.870 2305.210 3078.170 ;
        RECT 2400.590 3078.170 2400.890 3078.550 ;
        RECT 2401.510 3078.170 2401.810 3079.230 ;
        RECT 2449.350 3078.850 2449.650 3079.230 ;
        RECT 2498.110 3079.230 2546.250 3079.530 ;
        RECT 2449.350 3078.550 2497.490 3078.850 ;
        RECT 2400.590 3077.870 2401.810 3078.170 ;
        RECT 2497.190 3078.170 2497.490 3078.550 ;
        RECT 2498.110 3078.170 2498.410 3079.230 ;
        RECT 2545.950 3078.850 2546.250 3079.230 ;
        RECT 2594.710 3079.230 2670.235 3079.530 ;
        RECT 2545.950 3078.550 2594.090 3078.850 ;
        RECT 2497.190 3077.870 2498.410 3078.170 ;
        RECT 2593.790 3078.170 2594.090 3078.550 ;
        RECT 2594.710 3078.170 2595.010 3079.230 ;
        RECT 2669.905 3079.215 2670.235 3079.230 ;
        RECT 2704.405 3079.530 2704.735 3079.545 ;
        RECT 2787.205 3079.530 2787.535 3079.545 ;
=======
        RECT 2899.445 3079.530 2899.775 3079.545 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 3079.530 2924.800 3079.980 ;
        RECT 2899.445 3079.230 2924.800 3079.530 ;
        RECT 2899.445 3079.215 2899.775 3079.230 ;
        RECT 2917.600 3078.780 2924.800 3079.230 ;
<<<<<<< HEAD
        RECT 2884.510 3078.170 2884.810 3078.550 ;
        RECT 2883.590 3077.870 2884.810 3078.170 ;
        RECT 2042.925 3077.855 2043.255 3077.870 ;
        RECT 2090.765 3077.855 2091.095 3077.870 ;
        RECT 2173.310 3077.490 2173.690 3077.500 ;
        RECT 2207.605 3077.490 2207.935 3077.505 ;
        RECT 2173.310 3077.190 2207.935 3077.490 ;
        RECT 2173.310 3077.180 2173.690 3077.190 ;
        RECT 2207.605 3077.175 2207.935 3077.190 ;
        RECT 2752.910 3077.490 2753.290 3077.500 ;
        RECT 2787.205 3077.490 2787.535 3077.505 ;
        RECT 2752.910 3077.190 2787.535 3077.490 ;
        RECT 2752.910 3077.180 2753.290 3077.190 ;
        RECT 2787.205 3077.175 2787.535 3077.190 ;
        RECT 1943.105 1703.220 1943.435 1703.225 ;
        RECT 1943.105 1703.210 1943.690 1703.220 ;
        RECT 1942.880 1702.910 1943.690 1703.210 ;
        RECT 1943.105 1702.900 1943.690 1702.910 ;
        RECT 1943.105 1702.895 1943.435 1702.900 ;
      LAYER via3 ;
        RECT 1943.340 3079.220 1943.660 3079.540 ;
        RECT 2173.340 3078.540 2173.660 3078.860 ;
        RECT 2752.940 3078.540 2753.260 3078.860 ;
        RECT 2173.340 3077.180 2173.660 3077.500 ;
        RECT 2752.940 3077.180 2753.260 3077.500 ;
        RECT 1943.340 1702.900 1943.660 1703.220 ;
      LAYER met4 ;
        RECT 1943.335 3079.215 1943.665 3079.545 ;
        RECT 1943.350 1703.225 1943.650 3079.215 ;
        RECT 2173.335 3078.535 2173.665 3078.865 ;
        RECT 2752.935 3078.535 2753.265 3078.865 ;
        RECT 2173.350 3077.505 2173.650 3078.535 ;
        RECT 2752.950 3077.505 2753.250 3078.535 ;
        RECT 2173.335 3077.175 2173.665 3077.505 ;
        RECT 2752.935 3077.175 2753.265 3077.505 ;
        RECT 1943.335 1702.895 1943.665 1703.225 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1946.000 2166.970 1950.000 2167.120 ;
        RECT 1962.885 2166.970 1963.215 2166.985 ;
        RECT 1946.000 2166.670 1963.215 2166.970 ;
        RECT 1946.000 2166.520 1950.000 2166.670 ;
        RECT 1962.885 2166.655 1963.215 2166.670 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2230.685 1690.225 2231.775 1690.395 ;
      LAYER mcon ;
        RECT 2231.605 1690.225 2231.775 1690.395 ;
      LAYER met1 ;
        RECT 1943.200 1690.580 1946.560 1690.720 ;
        RECT 1943.200 1690.440 1943.340 1690.580 ;
        RECT 1943.110 1690.180 1943.430 1690.440 ;
        RECT 1946.420 1690.380 1946.560 1690.580 ;
        RECT 2230.625 1690.380 2230.915 1690.425 ;
        RECT 1946.420 1690.240 2230.915 1690.380 ;
        RECT 2230.625 1690.195 2230.915 1690.240 ;
        RECT 2231.545 1690.380 2231.835 1690.425 ;
        RECT 2901.290 1690.380 2901.610 1690.440 ;
        RECT 2231.545 1690.240 2901.610 1690.380 ;
        RECT 2231.545 1690.195 2231.835 1690.240 ;
        RECT 2901.290 1690.180 2901.610 1690.240 ;
      LAYER via ;
        RECT 1943.140 1690.180 1943.400 1690.440 ;
        RECT 2901.320 1690.180 2901.580 1690.440 ;
      LAYER met2 ;
        RECT 2901.310 3313.795 2901.590 3314.165 ;
        RECT 1942.210 1700.410 1942.490 1704.000 ;
        RECT 1942.210 1700.270 1943.340 1700.410 ;
        RECT 1942.210 1700.000 1942.490 1700.270 ;
        RECT 1943.200 1690.470 1943.340 1700.270 ;
        RECT 2901.380 1690.470 2901.520 3313.795 ;
        RECT 1943.140 1690.150 1943.400 1690.470 ;
        RECT 2901.320 1690.150 2901.580 1690.470 ;
      LAYER via2 ;
        RECT 2901.310 3313.840 2901.590 3314.120 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 3313.380 2924.800 3314.580 ;
=======
        RECT 2900.825 3314.130 2901.155 3314.145 ;
=======
        RECT 2901.285 3314.130 2901.615 3314.145 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 3314.130 2924.800 3314.580 ;
        RECT 2901.285 3313.830 2924.800 3314.130 ;
        RECT 2901.285 3313.815 2901.615 3313.830 ;
        RECT 2917.600 3313.380 2924.800 3313.830 ;
<<<<<<< HEAD
        RECT 1946.000 2033.690 1950.000 2033.840 ;
        RECT 1962.885 2033.690 1963.215 2033.705 ;
        RECT 1946.000 2033.390 1963.215 2033.690 ;
        RECT 1946.000 2033.240 1950.000 2033.390 ;
        RECT 1962.885 2033.375 1963.215 2033.390 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1917.810 3501.560 1918.130 3501.620 ;
        RECT 2879.210 3501.560 2879.530 3501.620 ;
        RECT 1917.810 3501.420 2879.530 3501.560 ;
        RECT 1917.810 3501.360 1918.130 3501.420 ;
        RECT 2879.210 3501.360 2879.530 3501.420 ;
      LAYER via ;
        RECT 1917.840 3501.360 1918.100 3501.620 ;
        RECT 2879.240 3501.360 2879.500 3501.620 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2879.090 3519.700 2879.650 3524.800 ;
=======
        RECT 2879.090 3517.600 2879.650 3524.800 ;
<<<<<<< HEAD
        RECT 2879.300 3501.845 2879.440 3517.600 ;
        RECT 2879.230 3501.475 2879.510 3501.845 ;
        RECT 1944.050 1703.130 1944.330 1704.000 ;
        RECT 1944.510 1703.130 1944.790 1703.245 ;
        RECT 1944.050 1702.990 1944.790 1703.130 ;
        RECT 1944.050 1700.000 1944.330 1702.990 ;
        RECT 1944.510 1702.875 1944.790 1702.990 ;
      LAYER via2 ;
        RECT 2879.230 3501.520 2879.510 3501.800 ;
        RECT 1944.510 1702.920 1944.790 1703.200 ;
      LAYER met3 ;
        RECT 1944.230 3501.810 1944.610 3501.820 ;
        RECT 2879.205 3501.810 2879.535 3501.825 ;
        RECT 1944.230 3501.510 2879.535 3501.810 ;
        RECT 1944.230 3501.500 1944.610 3501.510 ;
        RECT 2879.205 3501.495 2879.535 3501.510 ;
        RECT 1944.485 1703.220 1944.815 1703.225 ;
        RECT 1944.230 1703.210 1944.815 1703.220 ;
        RECT 1944.230 1702.910 1945.040 1703.210 ;
        RECT 1944.230 1702.900 1944.815 1702.910 ;
        RECT 1944.485 1702.895 1944.815 1702.900 ;
      LAYER via3 ;
        RECT 1944.260 3501.500 1944.580 3501.820 ;
        RECT 1944.260 1702.900 1944.580 1703.220 ;
      LAYER met4 ;
        RECT 1944.255 3501.495 1944.585 3501.825 ;
        RECT 1944.270 1703.225 1944.570 3501.495 ;
        RECT 1944.255 1702.895 1944.585 1703.225 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2879.300 3501.650 2879.440 3517.600 ;
        RECT 1917.840 3501.330 1918.100 3501.650 ;
        RECT 2879.240 3501.330 2879.500 3501.650 ;
        RECT 1917.900 2500.090 1918.040 3501.330 ;
        RECT 1914.150 2499.410 1914.430 2500.000 ;
        RECT 1916.060 2499.950 1918.040 2500.090 ;
        RECT 1916.060 2499.410 1916.200 2499.950 ;
        RECT 1914.150 2499.270 1916.200 2499.410 ;
        RECT 1914.150 2496.000 1914.430 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2553.605 3429.665 2553.775 3477.435 ;
        RECT 2553.145 3332.765 2553.315 3380.875 ;
        RECT 2553.605 2815.285 2553.775 2849.455 ;
        RECT 1945.945 1685.465 1946.115 1690.395 ;
        RECT 1993.785 1685.465 1993.955 1690.055 ;
        RECT 2231.145 1689.885 2232.695 1690.055 ;
      LAYER mcon ;
        RECT 2553.605 3477.265 2553.775 3477.435 ;
        RECT 2553.145 3380.705 2553.315 3380.875 ;
        RECT 2553.605 2849.285 2553.775 2849.455 ;
        RECT 1945.945 1690.225 1946.115 1690.395 ;
        RECT 1993.785 1689.885 1993.955 1690.055 ;
        RECT 2232.525 1689.885 2232.695 1690.055 ;
      LAYER met1 ;
        RECT 2553.530 3477.420 2553.850 3477.480 ;
        RECT 2553.335 3477.280 2553.850 3477.420 ;
        RECT 2553.530 3477.220 2553.850 3477.280 ;
        RECT 2553.545 3429.820 2553.835 3429.865 ;
        RECT 2553.990 3429.820 2554.310 3429.880 ;
        RECT 2553.545 3429.680 2554.310 3429.820 ;
        RECT 2553.545 3429.635 2553.835 3429.680 ;
        RECT 2553.990 3429.620 2554.310 3429.680 ;
        RECT 2553.070 3380.860 2553.390 3380.920 ;
        RECT 2552.875 3380.720 2553.390 3380.860 ;
        RECT 2553.070 3380.660 2553.390 3380.720 ;
        RECT 2553.085 3332.920 2553.375 3332.965 ;
        RECT 2553.530 3332.920 2553.850 3332.980 ;
        RECT 2553.085 3332.780 2553.850 3332.920 ;
        RECT 2553.085 3332.735 2553.375 3332.780 ;
        RECT 2553.530 3332.720 2553.850 3332.780 ;
        RECT 2553.070 3270.700 2553.390 3270.760 ;
        RECT 2553.990 3270.700 2554.310 3270.760 ;
        RECT 2553.070 3270.560 2554.310 3270.700 ;
        RECT 2553.070 3270.500 2553.390 3270.560 ;
        RECT 2553.990 3270.500 2554.310 3270.560 ;
        RECT 2553.070 3174.140 2553.390 3174.200 ;
        RECT 2553.990 3174.140 2554.310 3174.200 ;
        RECT 2553.070 3174.000 2554.310 3174.140 ;
        RECT 2553.070 3173.940 2553.390 3174.000 ;
        RECT 2553.990 3173.940 2554.310 3174.000 ;
        RECT 2553.070 2981.020 2553.390 2981.080 ;
        RECT 2553.990 2981.020 2554.310 2981.080 ;
        RECT 2553.070 2980.880 2554.310 2981.020 ;
        RECT 2553.070 2980.820 2553.390 2980.880 ;
        RECT 2553.990 2980.820 2554.310 2980.880 ;
        RECT 2552.150 2946.340 2552.470 2946.400 ;
        RECT 2553.530 2946.340 2553.850 2946.400 ;
        RECT 2552.150 2946.200 2553.850 2946.340 ;
        RECT 2552.150 2946.140 2552.470 2946.200 ;
        RECT 2553.530 2946.140 2553.850 2946.200 ;
        RECT 2553.530 2849.440 2553.850 2849.500 ;
        RECT 2553.335 2849.300 2553.850 2849.440 ;
        RECT 2553.530 2849.240 2553.850 2849.300 ;
        RECT 2553.545 2815.440 2553.835 2815.485 ;
        RECT 2554.450 2815.440 2554.770 2815.500 ;
        RECT 2553.545 2815.300 2554.770 2815.440 ;
        RECT 2553.545 2815.255 2553.835 2815.300 ;
        RECT 2554.450 2815.240 2554.770 2815.300 ;
        RECT 2553.530 2753.220 2553.850 2753.280 ;
        RECT 2554.910 2753.220 2555.230 2753.280 ;
        RECT 2553.530 2753.080 2555.230 2753.220 ;
        RECT 2553.530 2753.020 2553.850 2753.080 ;
        RECT 2554.910 2753.020 2555.230 2753.080 ;
        RECT 2554.910 2719.220 2555.230 2719.280 ;
        RECT 2554.540 2719.080 2555.230 2719.220 ;
        RECT 2554.540 2718.600 2554.680 2719.080 ;
        RECT 2554.910 2719.020 2555.230 2719.080 ;
        RECT 2554.450 2718.340 2554.770 2718.600 ;
        RECT 2554.450 2670.400 2554.770 2670.660 ;
        RECT 2554.540 2669.920 2554.680 2670.400 ;
        RECT 2554.910 2669.920 2555.230 2669.980 ;
        RECT 2554.540 2669.780 2555.230 2669.920 ;
        RECT 2554.910 2669.720 2555.230 2669.780 ;
        RECT 2554.910 2649.520 2555.230 2649.580 ;
        RECT 2555.830 2649.520 2556.150 2649.580 ;
        RECT 2554.910 2649.380 2556.150 2649.520 ;
        RECT 2554.910 2649.320 2555.230 2649.380 ;
        RECT 2555.830 2649.320 2556.150 2649.380 ;
        RECT 2554.910 2573.360 2555.230 2573.420 ;
        RECT 2555.830 2573.360 2556.150 2573.420 ;
        RECT 2554.910 2573.220 2556.150 2573.360 ;
        RECT 2554.910 2573.160 2555.230 2573.220 ;
        RECT 2555.830 2573.160 2556.150 2573.220 ;
        RECT 2553.990 2511.820 2554.310 2511.880 ;
        RECT 2554.910 2511.820 2555.230 2511.880 ;
        RECT 2553.990 2511.680 2555.230 2511.820 ;
        RECT 2553.990 2511.620 2554.310 2511.680 ;
        RECT 2554.910 2511.620 2555.230 2511.680 ;
        RECT 2553.070 2401.320 2553.390 2401.380 ;
        RECT 2553.990 2401.320 2554.310 2401.380 ;
        RECT 2553.070 2401.180 2554.310 2401.320 ;
        RECT 2553.070 2401.120 2553.390 2401.180 ;
        RECT 2553.990 2401.120 2554.310 2401.180 ;
        RECT 2553.070 2304.760 2553.390 2304.820 ;
        RECT 2553.990 2304.760 2554.310 2304.820 ;
        RECT 2553.070 2304.620 2554.310 2304.760 ;
        RECT 2553.070 2304.560 2553.390 2304.620 ;
        RECT 2553.990 2304.560 2554.310 2304.620 ;
        RECT 2553.070 2208.200 2553.390 2208.260 ;
        RECT 2553.990 2208.200 2554.310 2208.260 ;
        RECT 2553.070 2208.060 2554.310 2208.200 ;
        RECT 2553.070 2208.000 2553.390 2208.060 ;
        RECT 2553.990 2208.000 2554.310 2208.060 ;
        RECT 2553.070 2111.640 2553.390 2111.700 ;
        RECT 2553.990 2111.640 2554.310 2111.700 ;
        RECT 2553.070 2111.500 2554.310 2111.640 ;
        RECT 2553.070 2111.440 2553.390 2111.500 ;
        RECT 2553.990 2111.440 2554.310 2111.500 ;
        RECT 2553.070 2015.080 2553.390 2015.140 ;
        RECT 2553.990 2015.080 2554.310 2015.140 ;
        RECT 2553.070 2014.940 2554.310 2015.080 ;
        RECT 2553.070 2014.880 2553.390 2014.940 ;
        RECT 2553.990 2014.880 2554.310 2014.940 ;
        RECT 2553.070 1918.520 2553.390 1918.580 ;
        RECT 2553.990 1918.520 2554.310 1918.580 ;
        RECT 2553.070 1918.380 2554.310 1918.520 ;
        RECT 2553.070 1918.320 2553.390 1918.380 ;
        RECT 2553.990 1918.320 2554.310 1918.380 ;
        RECT 2553.070 1821.960 2553.390 1822.020 ;
        RECT 2553.990 1821.960 2554.310 1822.020 ;
        RECT 2553.070 1821.820 2554.310 1821.960 ;
        RECT 2553.070 1821.760 2553.390 1821.820 ;
        RECT 2553.990 1821.760 2554.310 1821.820 ;
        RECT 2553.070 1725.400 2553.390 1725.460 ;
        RECT 2553.990 1725.400 2554.310 1725.460 ;
        RECT 2553.070 1725.260 2554.310 1725.400 ;
        RECT 2553.070 1725.200 2553.390 1725.260 ;
        RECT 2553.990 1725.200 2554.310 1725.260 ;
        RECT 1943.570 1690.380 1943.890 1690.440 ;
        RECT 1945.885 1690.380 1946.175 1690.425 ;
        RECT 1943.570 1690.240 1946.175 1690.380 ;
        RECT 1943.570 1690.180 1943.890 1690.240 ;
        RECT 1945.885 1690.195 1946.175 1690.240 ;
        RECT 1993.725 1690.040 1994.015 1690.085 ;
        RECT 2231.085 1690.040 2231.375 1690.085 ;
        RECT 1993.725 1689.900 2231.375 1690.040 ;
        RECT 1993.725 1689.855 1994.015 1689.900 ;
        RECT 2231.085 1689.855 2231.375 1689.900 ;
        RECT 2232.465 1690.040 2232.755 1690.085 ;
        RECT 2553.070 1690.040 2553.390 1690.100 ;
        RECT 2232.465 1689.900 2553.390 1690.040 ;
        RECT 2232.465 1689.855 2232.755 1689.900 ;
        RECT 2553.070 1689.840 2553.390 1689.900 ;
        RECT 1945.885 1685.620 1946.175 1685.665 ;
        RECT 1993.725 1685.620 1994.015 1685.665 ;
        RECT 1945.885 1685.480 1994.015 1685.620 ;
        RECT 1945.885 1685.435 1946.175 1685.480 ;
        RECT 1993.725 1685.435 1994.015 1685.480 ;
      LAYER via ;
        RECT 2553.560 3477.220 2553.820 3477.480 ;
        RECT 2554.020 3429.620 2554.280 3429.880 ;
        RECT 2553.100 3380.660 2553.360 3380.920 ;
        RECT 2553.560 3332.720 2553.820 3332.980 ;
        RECT 2553.100 3270.500 2553.360 3270.760 ;
        RECT 2554.020 3270.500 2554.280 3270.760 ;
        RECT 2553.100 3173.940 2553.360 3174.200 ;
        RECT 2554.020 3173.940 2554.280 3174.200 ;
        RECT 2553.100 2980.820 2553.360 2981.080 ;
        RECT 2554.020 2980.820 2554.280 2981.080 ;
        RECT 2552.180 2946.140 2552.440 2946.400 ;
        RECT 2553.560 2946.140 2553.820 2946.400 ;
        RECT 2553.560 2849.240 2553.820 2849.500 ;
        RECT 2554.480 2815.240 2554.740 2815.500 ;
        RECT 2553.560 2753.020 2553.820 2753.280 ;
        RECT 2554.940 2753.020 2555.200 2753.280 ;
        RECT 2554.940 2719.020 2555.200 2719.280 ;
        RECT 2554.480 2718.340 2554.740 2718.600 ;
        RECT 2554.480 2670.400 2554.740 2670.660 ;
        RECT 2554.940 2669.720 2555.200 2669.980 ;
        RECT 2554.940 2649.320 2555.200 2649.580 ;
        RECT 2555.860 2649.320 2556.120 2649.580 ;
        RECT 2554.940 2573.160 2555.200 2573.420 ;
        RECT 2555.860 2573.160 2556.120 2573.420 ;
        RECT 2554.020 2511.620 2554.280 2511.880 ;
        RECT 2554.940 2511.620 2555.200 2511.880 ;
        RECT 2553.100 2401.120 2553.360 2401.380 ;
        RECT 2554.020 2401.120 2554.280 2401.380 ;
        RECT 2553.100 2304.560 2553.360 2304.820 ;
        RECT 2554.020 2304.560 2554.280 2304.820 ;
        RECT 2553.100 2208.000 2553.360 2208.260 ;
        RECT 2554.020 2208.000 2554.280 2208.260 ;
        RECT 2553.100 2111.440 2553.360 2111.700 ;
        RECT 2554.020 2111.440 2554.280 2111.700 ;
        RECT 2553.100 2014.880 2553.360 2015.140 ;
        RECT 2554.020 2014.880 2554.280 2015.140 ;
        RECT 2553.100 1918.320 2553.360 1918.580 ;
        RECT 2554.020 1918.320 2554.280 1918.580 ;
        RECT 2553.100 1821.760 2553.360 1822.020 ;
        RECT 2554.020 1821.760 2554.280 1822.020 ;
        RECT 2553.100 1725.200 2553.360 1725.460 ;
        RECT 2554.020 1725.200 2554.280 1725.460 ;
        RECT 1943.600 1690.180 1943.860 1690.440 ;
        RECT 2553.100 1689.840 2553.360 1690.100 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2554.790 3519.700 2555.350 3524.800 ;
=======
        RECT 2554.790 3517.600 2555.350 3524.800 ;
<<<<<<< HEAD
        RECT 2555.000 3501.650 2555.140 3517.600 ;
        RECT 1938.540 3501.330 1938.800 3501.650 ;
        RECT 2554.940 3501.330 2555.200 3501.650 ;
        RECT 1938.600 2516.330 1938.740 3501.330 ;
        RECT 1933.020 2516.010 1933.280 2516.330 ;
        RECT 1938.540 2516.010 1938.800 2516.330 ;
        RECT 1933.080 2500.000 1933.220 2516.010 ;
        RECT 1933.010 2496.000 1933.290 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2555.000 3511.930 2555.140 3517.600 ;
        RECT 2553.620 3511.790 2555.140 3511.930 ;
        RECT 2553.620 3477.510 2553.760 3511.790 ;
        RECT 2553.560 3477.190 2553.820 3477.510 ;
        RECT 2554.020 3429.590 2554.280 3429.910 ;
        RECT 2554.080 3394.970 2554.220 3429.590 ;
        RECT 2553.160 3394.830 2554.220 3394.970 ;
        RECT 2553.160 3380.950 2553.300 3394.830 ;
        RECT 2553.100 3380.630 2553.360 3380.950 ;
        RECT 2553.560 3332.690 2553.820 3333.010 ;
        RECT 2553.620 3298.410 2553.760 3332.690 ;
        RECT 2553.620 3298.270 2554.220 3298.410 ;
        RECT 2554.080 3270.790 2554.220 3298.270 ;
        RECT 2553.100 3270.470 2553.360 3270.790 ;
        RECT 2554.020 3270.470 2554.280 3270.790 ;
        RECT 2553.160 3222.250 2553.300 3270.470 ;
        RECT 2553.160 3222.110 2554.220 3222.250 ;
        RECT 2554.080 3174.230 2554.220 3222.110 ;
        RECT 2553.100 3173.910 2553.360 3174.230 ;
        RECT 2554.020 3173.910 2554.280 3174.230 ;
        RECT 2553.160 3125.690 2553.300 3173.910 ;
        RECT 2553.160 3125.550 2554.220 3125.690 ;
        RECT 2554.080 2981.110 2554.220 3125.550 ;
        RECT 2553.100 2980.850 2553.360 2981.110 ;
        RECT 2553.100 2980.790 2553.760 2980.850 ;
        RECT 2554.020 2980.790 2554.280 2981.110 ;
        RECT 2553.160 2980.710 2553.760 2980.790 ;
        RECT 2553.620 2980.170 2553.760 2980.710 ;
        RECT 2553.620 2980.030 2554.220 2980.170 ;
        RECT 2554.080 2959.770 2554.220 2980.030 ;
        RECT 2553.620 2959.630 2554.220 2959.770 ;
        RECT 2553.620 2946.430 2553.760 2959.630 ;
        RECT 2552.180 2946.110 2552.440 2946.430 ;
        RECT 2553.560 2946.110 2553.820 2946.430 ;
        RECT 2552.240 2898.685 2552.380 2946.110 ;
        RECT 2552.170 2898.315 2552.450 2898.685 ;
        RECT 2553.090 2898.315 2553.370 2898.685 ;
        RECT 2553.160 2863.210 2553.300 2898.315 ;
        RECT 2553.160 2863.070 2553.760 2863.210 ;
        RECT 2553.620 2849.530 2553.760 2863.070 ;
        RECT 2553.560 2849.210 2553.820 2849.530 ;
        RECT 2554.480 2815.210 2554.740 2815.530 ;
        RECT 2554.540 2801.445 2554.680 2815.210 ;
        RECT 2553.550 2801.075 2553.830 2801.445 ;
        RECT 2554.470 2801.075 2554.750 2801.445 ;
        RECT 2553.620 2753.310 2553.760 2801.075 ;
        RECT 2553.560 2752.990 2553.820 2753.310 ;
        RECT 2554.940 2752.990 2555.200 2753.310 ;
        RECT 2555.000 2719.310 2555.140 2752.990 ;
        RECT 2554.940 2718.990 2555.200 2719.310 ;
        RECT 2554.480 2718.310 2554.740 2718.630 ;
        RECT 2554.540 2670.690 2554.680 2718.310 ;
        RECT 2554.480 2670.370 2554.740 2670.690 ;
        RECT 2554.940 2669.690 2555.200 2670.010 ;
        RECT 2555.000 2649.610 2555.140 2669.690 ;
        RECT 2554.940 2649.290 2555.200 2649.610 ;
        RECT 2555.860 2649.290 2556.120 2649.610 ;
        RECT 2555.920 2573.450 2556.060 2649.290 ;
        RECT 2554.940 2573.130 2555.200 2573.450 ;
        RECT 2555.860 2573.130 2556.120 2573.450 ;
        RECT 2555.000 2511.910 2555.140 2573.130 ;
        RECT 2554.020 2511.765 2554.280 2511.910 ;
        RECT 2552.630 2511.395 2552.910 2511.765 ;
        RECT 2554.010 2511.395 2554.290 2511.765 ;
        RECT 2554.940 2511.590 2555.200 2511.910 ;
        RECT 2552.700 2463.485 2552.840 2511.395 ;
        RECT 2552.630 2463.115 2552.910 2463.485 ;
        RECT 2553.550 2463.115 2553.830 2463.485 ;
        RECT 2553.620 2449.770 2553.760 2463.115 ;
        RECT 2553.620 2449.630 2554.220 2449.770 ;
        RECT 2554.080 2401.410 2554.220 2449.630 ;
        RECT 2553.100 2401.090 2553.360 2401.410 ;
        RECT 2554.020 2401.090 2554.280 2401.410 ;
        RECT 2553.160 2400.810 2553.300 2401.090 ;
        RECT 2553.160 2400.670 2553.760 2400.810 ;
        RECT 2553.620 2353.210 2553.760 2400.670 ;
        RECT 2553.620 2353.070 2554.220 2353.210 ;
        RECT 2554.080 2304.850 2554.220 2353.070 ;
        RECT 2553.100 2304.530 2553.360 2304.850 ;
        RECT 2554.020 2304.530 2554.280 2304.850 ;
        RECT 2553.160 2304.250 2553.300 2304.530 ;
        RECT 2553.160 2304.110 2553.760 2304.250 ;
        RECT 2553.620 2256.650 2553.760 2304.110 ;
        RECT 2553.620 2256.510 2554.220 2256.650 ;
        RECT 2554.080 2208.290 2554.220 2256.510 ;
        RECT 2553.100 2207.970 2553.360 2208.290 ;
        RECT 2554.020 2207.970 2554.280 2208.290 ;
        RECT 2553.160 2207.690 2553.300 2207.970 ;
        RECT 2553.160 2207.550 2553.760 2207.690 ;
        RECT 2553.620 2160.090 2553.760 2207.550 ;
        RECT 2553.620 2159.950 2554.220 2160.090 ;
        RECT 2554.080 2111.730 2554.220 2159.950 ;
        RECT 2553.100 2111.410 2553.360 2111.730 ;
        RECT 2554.020 2111.410 2554.280 2111.730 ;
        RECT 2553.160 2111.130 2553.300 2111.410 ;
        RECT 2553.160 2110.990 2553.760 2111.130 ;
        RECT 2553.620 2063.530 2553.760 2110.990 ;
        RECT 2553.620 2063.390 2554.220 2063.530 ;
        RECT 2554.080 2015.170 2554.220 2063.390 ;
        RECT 2553.100 2014.850 2553.360 2015.170 ;
        RECT 2554.020 2014.850 2554.280 2015.170 ;
        RECT 2553.160 2014.570 2553.300 2014.850 ;
        RECT 2553.160 2014.430 2553.760 2014.570 ;
        RECT 2553.620 1966.970 2553.760 2014.430 ;
        RECT 2553.620 1966.830 2554.220 1966.970 ;
        RECT 2554.080 1918.610 2554.220 1966.830 ;
        RECT 2553.100 1918.290 2553.360 1918.610 ;
        RECT 2554.020 1918.290 2554.280 1918.610 ;
        RECT 2553.160 1918.010 2553.300 1918.290 ;
        RECT 2553.160 1917.870 2553.760 1918.010 ;
        RECT 2553.620 1870.410 2553.760 1917.870 ;
        RECT 2553.620 1870.270 2554.220 1870.410 ;
        RECT 2554.080 1822.050 2554.220 1870.270 ;
        RECT 2553.100 1821.730 2553.360 1822.050 ;
        RECT 2554.020 1821.730 2554.280 1822.050 ;
        RECT 2553.160 1773.170 2553.300 1821.730 ;
        RECT 2553.160 1773.030 2554.220 1773.170 ;
        RECT 2554.080 1725.490 2554.220 1773.030 ;
        RECT 2553.100 1725.170 2553.360 1725.490 ;
        RECT 2554.020 1725.170 2554.280 1725.490 ;
        RECT 1943.590 1700.000 1943.870 1704.000 ;
        RECT 1943.660 1690.470 1943.800 1700.000 ;
        RECT 1943.600 1690.150 1943.860 1690.470 ;
        RECT 2553.160 1690.130 2553.300 1725.170 ;
        RECT 2553.100 1689.810 2553.360 1690.130 ;
      LAYER via2 ;
        RECT 2552.170 2898.360 2552.450 2898.640 ;
        RECT 2553.090 2898.360 2553.370 2898.640 ;
        RECT 2553.550 2801.120 2553.830 2801.400 ;
        RECT 2554.470 2801.120 2554.750 2801.400 ;
        RECT 2552.630 2511.440 2552.910 2511.720 ;
        RECT 2554.010 2511.440 2554.290 2511.720 ;
        RECT 2552.630 2463.160 2552.910 2463.440 ;
        RECT 2553.550 2463.160 2553.830 2463.440 ;
      LAYER met3 ;
        RECT 2552.145 2898.650 2552.475 2898.665 ;
        RECT 2553.065 2898.650 2553.395 2898.665 ;
        RECT 2552.145 2898.350 2553.395 2898.650 ;
        RECT 2552.145 2898.335 2552.475 2898.350 ;
        RECT 2553.065 2898.335 2553.395 2898.350 ;
        RECT 2553.525 2801.410 2553.855 2801.425 ;
        RECT 2554.445 2801.410 2554.775 2801.425 ;
        RECT 2553.525 2801.110 2554.775 2801.410 ;
        RECT 2553.525 2801.095 2553.855 2801.110 ;
        RECT 2554.445 2801.095 2554.775 2801.110 ;
        RECT 2552.605 2511.730 2552.935 2511.745 ;
        RECT 2553.985 2511.730 2554.315 2511.745 ;
        RECT 2552.605 2511.430 2554.315 2511.730 ;
        RECT 2552.605 2511.415 2552.935 2511.430 ;
        RECT 2553.985 2511.415 2554.315 2511.430 ;
        RECT 2552.605 2463.450 2552.935 2463.465 ;
        RECT 2553.525 2463.450 2553.855 2463.465 ;
        RECT 2552.605 2463.150 2553.855 2463.450 ;
        RECT 2552.605 2463.135 2552.935 2463.150 ;
        RECT 2553.525 2463.135 2553.855 2463.150 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2227.925 3422.185 2228.095 3463.835 ;
        RECT 2230.685 3332.765 2230.855 3415.555 ;
        RECT 2229.765 3104.965 2229.935 3139.475 ;
        RECT 2229.305 2753.065 2229.475 2801.175 ;
        RECT 2229.765 2428.705 2229.935 2463.215 ;
        RECT 2229.765 2331.805 2229.935 2366.655 ;
        RECT 2229.305 1973.445 2229.475 2021.555 ;
        RECT 2230.685 1787.125 2230.855 1835.235 ;
        RECT 2230.225 1690.565 2230.395 1738.675 ;
      LAYER mcon ;
        RECT 2227.925 3463.665 2228.095 3463.835 ;
        RECT 2230.685 3415.385 2230.855 3415.555 ;
        RECT 2229.765 3139.305 2229.935 3139.475 ;
        RECT 2229.305 2801.005 2229.475 2801.175 ;
        RECT 2229.765 2463.045 2229.935 2463.215 ;
        RECT 2229.765 2366.485 2229.935 2366.655 ;
        RECT 2229.305 2021.385 2229.475 2021.555 ;
        RECT 2230.685 1835.065 2230.855 1835.235 ;
        RECT 2230.225 1738.505 2230.395 1738.675 ;
      LAYER met1 ;
        RECT 2227.850 3470.620 2228.170 3470.680 ;
        RECT 2229.690 3470.620 2230.010 3470.680 ;
        RECT 2227.850 3470.480 2230.010 3470.620 ;
        RECT 2227.850 3470.420 2228.170 3470.480 ;
        RECT 2229.690 3470.420 2230.010 3470.480 ;
        RECT 2227.850 3463.820 2228.170 3463.880 ;
        RECT 2227.655 3463.680 2228.170 3463.820 ;
        RECT 2227.850 3463.620 2228.170 3463.680 ;
        RECT 2227.865 3422.340 2228.155 3422.385 ;
        RECT 2228.770 3422.340 2229.090 3422.400 ;
        RECT 2227.865 3422.200 2229.090 3422.340 ;
        RECT 2227.865 3422.155 2228.155 3422.200 ;
        RECT 2228.770 3422.140 2229.090 3422.200 ;
        RECT 2228.770 3415.540 2229.090 3415.600 ;
        RECT 2230.625 3415.540 2230.915 3415.585 ;
        RECT 2228.770 3415.400 2230.915 3415.540 ;
        RECT 2228.770 3415.340 2229.090 3415.400 ;
        RECT 2230.625 3415.355 2230.915 3415.400 ;
        RECT 2230.625 3332.920 2230.915 3332.965 ;
        RECT 2231.070 3332.920 2231.390 3332.980 ;
        RECT 2230.625 3332.780 2231.390 3332.920 ;
        RECT 2230.625 3332.735 2230.915 3332.780 ;
        RECT 2231.070 3332.720 2231.390 3332.780 ;
        RECT 2229.690 3236.360 2230.010 3236.420 ;
        RECT 2230.150 3236.360 2230.470 3236.420 ;
        RECT 2229.690 3236.220 2230.470 3236.360 ;
        RECT 2229.690 3236.160 2230.010 3236.220 ;
        RECT 2230.150 3236.160 2230.470 3236.220 ;
        RECT 2229.690 3202.020 2230.010 3202.080 ;
        RECT 2230.150 3202.020 2230.470 3202.080 ;
        RECT 2229.690 3201.880 2230.470 3202.020 ;
        RECT 2229.690 3201.820 2230.010 3201.880 ;
        RECT 2230.150 3201.820 2230.470 3201.880 ;
        RECT 2229.230 3153.400 2229.550 3153.460 ;
        RECT 2230.150 3153.400 2230.470 3153.460 ;
        RECT 2229.230 3153.260 2230.470 3153.400 ;
        RECT 2229.230 3153.200 2229.550 3153.260 ;
        RECT 2230.150 3153.200 2230.470 3153.260 ;
        RECT 2229.690 3139.460 2230.010 3139.520 ;
        RECT 2229.495 3139.320 2230.010 3139.460 ;
        RECT 2229.690 3139.260 2230.010 3139.320 ;
        RECT 2229.705 3105.120 2229.995 3105.165 ;
        RECT 2230.610 3105.120 2230.930 3105.180 ;
        RECT 2229.705 3104.980 2230.930 3105.120 ;
        RECT 2229.705 3104.935 2229.995 3104.980 ;
        RECT 2230.610 3104.920 2230.930 3104.980 ;
        RECT 2230.610 3056.640 2230.930 3056.900 ;
        RECT 2230.700 3056.160 2230.840 3056.640 ;
        RECT 2231.070 3056.160 2231.390 3056.220 ;
        RECT 2230.700 3056.020 2231.390 3056.160 ;
        RECT 2231.070 3055.960 2231.390 3056.020 ;
        RECT 2231.070 2912.340 2231.390 2912.400 ;
        RECT 2230.700 2912.200 2231.390 2912.340 ;
        RECT 2230.700 2911.720 2230.840 2912.200 ;
        RECT 2231.070 2912.140 2231.390 2912.200 ;
        RECT 2230.610 2911.460 2230.930 2911.720 ;
        RECT 2229.230 2815.580 2229.550 2815.840 ;
        RECT 2229.320 2815.160 2229.460 2815.580 ;
        RECT 2229.230 2814.900 2229.550 2815.160 ;
        RECT 2229.230 2801.160 2229.550 2801.220 ;
        RECT 2229.035 2801.020 2229.550 2801.160 ;
        RECT 2229.230 2800.960 2229.550 2801.020 ;
        RECT 2229.245 2753.220 2229.535 2753.265 ;
        RECT 2230.150 2753.220 2230.470 2753.280 ;
        RECT 2229.245 2753.080 2230.470 2753.220 ;
        RECT 2229.245 2753.035 2229.535 2753.080 ;
        RECT 2230.150 2753.020 2230.470 2753.080 ;
        RECT 2229.230 2718.200 2229.550 2718.260 ;
        RECT 2230.150 2718.200 2230.470 2718.260 ;
        RECT 2229.230 2718.060 2230.470 2718.200 ;
        RECT 2229.230 2718.000 2229.550 2718.060 ;
        RECT 2230.150 2718.000 2230.470 2718.060 ;
        RECT 2229.230 2670.260 2229.550 2670.320 ;
        RECT 2230.150 2670.260 2230.470 2670.320 ;
        RECT 2229.230 2670.120 2230.470 2670.260 ;
        RECT 2229.230 2670.060 2229.550 2670.120 ;
        RECT 2230.150 2670.060 2230.470 2670.120 ;
        RECT 2230.150 2622.120 2230.470 2622.380 ;
        RECT 2230.240 2621.980 2230.380 2622.120 ;
        RECT 2230.610 2621.980 2230.930 2622.040 ;
        RECT 2230.240 2621.840 2230.930 2621.980 ;
        RECT 2230.610 2621.780 2230.930 2621.840 ;
        RECT 2229.690 2560.100 2230.010 2560.160 ;
        RECT 2231.070 2560.100 2231.390 2560.160 ;
        RECT 2229.690 2559.960 2231.390 2560.100 ;
        RECT 2229.690 2559.900 2230.010 2559.960 ;
        RECT 2231.070 2559.900 2231.390 2559.960 ;
        RECT 2230.150 2511.820 2230.470 2511.880 ;
        RECT 2231.070 2511.820 2231.390 2511.880 ;
        RECT 2230.150 2511.680 2231.390 2511.820 ;
        RECT 2230.150 2511.620 2230.470 2511.680 ;
        RECT 2231.070 2511.620 2231.390 2511.680 ;
        RECT 2229.690 2463.200 2230.010 2463.260 ;
        RECT 2229.495 2463.060 2230.010 2463.200 ;
        RECT 2229.690 2463.000 2230.010 2463.060 ;
        RECT 2229.690 2428.860 2230.010 2428.920 ;
        RECT 2229.495 2428.720 2230.010 2428.860 ;
        RECT 2229.690 2428.660 2230.010 2428.720 ;
        RECT 2229.230 2380.580 2229.550 2380.640 ;
        RECT 2230.150 2380.580 2230.470 2380.640 ;
        RECT 2229.230 2380.440 2230.470 2380.580 ;
        RECT 2229.230 2380.380 2229.550 2380.440 ;
        RECT 2230.150 2380.380 2230.470 2380.440 ;
        RECT 2229.690 2366.640 2230.010 2366.700 ;
        RECT 2229.495 2366.500 2230.010 2366.640 ;
        RECT 2229.690 2366.440 2230.010 2366.500 ;
        RECT 2229.690 2331.960 2230.010 2332.020 ;
        RECT 2229.495 2331.820 2230.010 2331.960 ;
        RECT 2229.690 2331.760 2230.010 2331.820 ;
        RECT 2228.770 2235.540 2229.090 2235.800 ;
        RECT 2228.860 2235.400 2229.000 2235.540 ;
        RECT 2229.230 2235.400 2229.550 2235.460 ;
        RECT 2228.860 2235.260 2229.550 2235.400 ;
        RECT 2229.230 2235.200 2229.550 2235.260 ;
        RECT 2227.850 2221.800 2228.170 2221.860 ;
        RECT 2229.230 2221.800 2229.550 2221.860 ;
        RECT 2227.850 2221.660 2229.550 2221.800 ;
        RECT 2227.850 2221.600 2228.170 2221.660 ;
        RECT 2229.230 2221.600 2229.550 2221.660 ;
        RECT 2227.850 2125.240 2228.170 2125.300 ;
        RECT 2229.230 2125.240 2229.550 2125.300 ;
        RECT 2227.850 2125.100 2229.550 2125.240 ;
        RECT 2227.850 2125.040 2228.170 2125.100 ;
        RECT 2229.230 2125.040 2229.550 2125.100 ;
        RECT 2228.770 2042.420 2229.090 2042.680 ;
        RECT 2228.860 2041.940 2229.000 2042.420 ;
        RECT 2229.230 2041.940 2229.550 2042.000 ;
        RECT 2228.860 2041.800 2229.550 2041.940 ;
        RECT 2229.230 2041.740 2229.550 2041.800 ;
        RECT 2229.230 2021.540 2229.550 2021.600 ;
        RECT 2229.035 2021.400 2229.550 2021.540 ;
        RECT 2229.230 2021.340 2229.550 2021.400 ;
        RECT 2229.245 1973.600 2229.535 1973.645 ;
        RECT 2229.690 1973.600 2230.010 1973.660 ;
        RECT 2229.245 1973.460 2230.010 1973.600 ;
        RECT 2229.245 1973.415 2229.535 1973.460 ;
        RECT 2229.690 1973.400 2230.010 1973.460 ;
        RECT 2229.690 1931.920 2230.010 1932.180 ;
        RECT 2229.780 1931.500 2229.920 1931.920 ;
        RECT 2229.690 1931.240 2230.010 1931.500 ;
        RECT 2229.690 1897.580 2230.010 1897.840 ;
        RECT 2229.780 1897.160 2229.920 1897.580 ;
        RECT 2229.690 1896.900 2230.010 1897.160 ;
        RECT 2230.610 1835.220 2230.930 1835.280 ;
        RECT 2230.415 1835.080 2230.930 1835.220 ;
        RECT 2230.610 1835.020 2230.930 1835.080 ;
        RECT 2230.625 1787.280 2230.915 1787.325 ;
        RECT 2231.070 1787.280 2231.390 1787.340 ;
        RECT 2230.625 1787.140 2231.390 1787.280 ;
        RECT 2230.625 1787.095 2230.915 1787.140 ;
        RECT 2231.070 1787.080 2231.390 1787.140 ;
        RECT 2230.150 1738.660 2230.470 1738.720 ;
        RECT 2229.955 1738.520 2230.470 1738.660 ;
        RECT 2230.150 1738.460 2230.470 1738.520 ;
        RECT 2230.165 1690.720 2230.455 1690.765 ;
        RECT 2231.070 1690.720 2231.390 1690.780 ;
        RECT 2230.165 1690.580 2231.390 1690.720 ;
        RECT 2230.165 1690.535 2230.455 1690.580 ;
        RECT 2231.070 1690.520 2231.390 1690.580 ;
        RECT 1945.410 1685.280 1945.730 1685.340 ;
        RECT 2231.070 1685.280 2231.390 1685.340 ;
        RECT 1945.410 1685.140 2231.390 1685.280 ;
        RECT 1945.410 1685.080 1945.730 1685.140 ;
        RECT 2231.070 1685.080 2231.390 1685.140 ;
      LAYER via ;
        RECT 2227.880 3470.420 2228.140 3470.680 ;
        RECT 2229.720 3470.420 2229.980 3470.680 ;
        RECT 2227.880 3463.620 2228.140 3463.880 ;
        RECT 2228.800 3422.140 2229.060 3422.400 ;
        RECT 2228.800 3415.340 2229.060 3415.600 ;
        RECT 2231.100 3332.720 2231.360 3332.980 ;
        RECT 2229.720 3236.160 2229.980 3236.420 ;
        RECT 2230.180 3236.160 2230.440 3236.420 ;
        RECT 2229.720 3201.820 2229.980 3202.080 ;
        RECT 2230.180 3201.820 2230.440 3202.080 ;
        RECT 2229.260 3153.200 2229.520 3153.460 ;
        RECT 2230.180 3153.200 2230.440 3153.460 ;
        RECT 2229.720 3139.260 2229.980 3139.520 ;
        RECT 2230.640 3104.920 2230.900 3105.180 ;
        RECT 2230.640 3056.640 2230.900 3056.900 ;
        RECT 2231.100 3055.960 2231.360 3056.220 ;
        RECT 2231.100 2912.140 2231.360 2912.400 ;
        RECT 2230.640 2911.460 2230.900 2911.720 ;
        RECT 2229.260 2815.580 2229.520 2815.840 ;
        RECT 2229.260 2814.900 2229.520 2815.160 ;
        RECT 2229.260 2800.960 2229.520 2801.220 ;
        RECT 2230.180 2753.020 2230.440 2753.280 ;
        RECT 2229.260 2718.000 2229.520 2718.260 ;
        RECT 2230.180 2718.000 2230.440 2718.260 ;
        RECT 2229.260 2670.060 2229.520 2670.320 ;
        RECT 2230.180 2670.060 2230.440 2670.320 ;
        RECT 2230.180 2622.120 2230.440 2622.380 ;
        RECT 2230.640 2621.780 2230.900 2622.040 ;
        RECT 2229.720 2559.900 2229.980 2560.160 ;
        RECT 2231.100 2559.900 2231.360 2560.160 ;
        RECT 2230.180 2511.620 2230.440 2511.880 ;
        RECT 2231.100 2511.620 2231.360 2511.880 ;
        RECT 2229.720 2463.000 2229.980 2463.260 ;
        RECT 2229.720 2428.660 2229.980 2428.920 ;
        RECT 2229.260 2380.380 2229.520 2380.640 ;
        RECT 2230.180 2380.380 2230.440 2380.640 ;
        RECT 2229.720 2366.440 2229.980 2366.700 ;
        RECT 2229.720 2331.760 2229.980 2332.020 ;
        RECT 2228.800 2235.540 2229.060 2235.800 ;
        RECT 2229.260 2235.200 2229.520 2235.460 ;
        RECT 2227.880 2221.600 2228.140 2221.860 ;
        RECT 2229.260 2221.600 2229.520 2221.860 ;
        RECT 2227.880 2125.040 2228.140 2125.300 ;
        RECT 2229.260 2125.040 2229.520 2125.300 ;
        RECT 2228.800 2042.420 2229.060 2042.680 ;
        RECT 2229.260 2041.740 2229.520 2042.000 ;
        RECT 2229.260 2021.340 2229.520 2021.600 ;
        RECT 2229.720 1973.400 2229.980 1973.660 ;
        RECT 2229.720 1931.920 2229.980 1932.180 ;
        RECT 2229.720 1931.240 2229.980 1931.500 ;
        RECT 2229.720 1897.580 2229.980 1897.840 ;
        RECT 2229.720 1896.900 2229.980 1897.160 ;
        RECT 2230.640 1835.020 2230.900 1835.280 ;
        RECT 2231.100 1787.080 2231.360 1787.340 ;
        RECT 2230.180 1738.460 2230.440 1738.720 ;
        RECT 2231.100 1690.520 2231.360 1690.780 ;
        RECT 1945.440 1685.080 1945.700 1685.340 ;
        RECT 2231.100 1685.080 2231.360 1685.340 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2230.490 3519.700 2231.050 3524.800 ;
=======
        RECT 2230.490 3517.600 2231.050 3524.800 ;
        RECT 2230.700 3517.370 2230.840 3517.600 ;
        RECT 2229.780 3517.230 2230.840 3517.370 ;
        RECT 2229.780 3470.710 2229.920 3517.230 ;
        RECT 2227.880 3470.390 2228.140 3470.710 ;
        RECT 2229.720 3470.390 2229.980 3470.710 ;
        RECT 2227.940 3463.910 2228.080 3470.390 ;
        RECT 2227.880 3463.590 2228.140 3463.910 ;
        RECT 2228.800 3422.110 2229.060 3422.430 ;
        RECT 2228.860 3415.630 2229.000 3422.110 ;
        RECT 2228.800 3415.310 2229.060 3415.630 ;
        RECT 2231.100 3332.690 2231.360 3333.010 ;
        RECT 2231.160 3298.410 2231.300 3332.690 ;
        RECT 2230.240 3298.270 2231.300 3298.410 ;
        RECT 2230.240 3236.450 2230.380 3298.270 ;
        RECT 2229.720 3236.130 2229.980 3236.450 ;
        RECT 2230.180 3236.130 2230.440 3236.450 ;
        RECT 2229.780 3202.110 2229.920 3236.130 ;
        RECT 2229.720 3201.790 2229.980 3202.110 ;
        RECT 2230.180 3201.790 2230.440 3202.110 ;
        RECT 2230.240 3153.490 2230.380 3201.790 ;
        RECT 2229.260 3153.170 2229.520 3153.490 ;
        RECT 2230.180 3153.170 2230.440 3153.490 ;
        RECT 2229.320 3152.890 2229.460 3153.170 ;
        RECT 2229.320 3152.750 2229.920 3152.890 ;
        RECT 2229.780 3139.550 2229.920 3152.750 ;
        RECT 2229.720 3139.230 2229.980 3139.550 ;
        RECT 2230.640 3104.890 2230.900 3105.210 ;
        RECT 2230.700 3056.930 2230.840 3104.890 ;
        RECT 2230.640 3056.610 2230.900 3056.930 ;
        RECT 2231.100 3055.930 2231.360 3056.250 ;
        RECT 2231.160 3036.045 2231.300 3055.930 ;
        RECT 2231.090 3035.675 2231.370 3036.045 ;
        RECT 2231.090 2959.515 2231.370 2959.885 ;
        RECT 2231.160 2912.430 2231.300 2959.515 ;
        RECT 2231.100 2912.110 2231.360 2912.430 ;
        RECT 2230.640 2911.430 2230.900 2911.750 ;
        RECT 2230.700 2863.210 2230.840 2911.430 ;
        RECT 2229.780 2863.070 2230.840 2863.210 ;
        RECT 2229.780 2849.610 2229.920 2863.070 ;
        RECT 2229.320 2849.470 2229.920 2849.610 ;
        RECT 2229.320 2815.870 2229.460 2849.470 ;
        RECT 2229.260 2815.550 2229.520 2815.870 ;
        RECT 2229.260 2814.870 2229.520 2815.190 ;
        RECT 2229.320 2801.250 2229.460 2814.870 ;
        RECT 2229.260 2800.930 2229.520 2801.250 ;
        RECT 2230.180 2752.990 2230.440 2753.310 ;
        RECT 2230.240 2718.290 2230.380 2752.990 ;
        RECT 2229.260 2717.970 2229.520 2718.290 ;
        RECT 2230.180 2717.970 2230.440 2718.290 ;
        RECT 2229.320 2670.350 2229.460 2717.970 ;
        RECT 2229.260 2670.030 2229.520 2670.350 ;
        RECT 2230.180 2670.030 2230.440 2670.350 ;
        RECT 2230.240 2622.410 2230.380 2670.030 ;
        RECT 2230.180 2622.090 2230.440 2622.410 ;
        RECT 2230.640 2621.750 2230.900 2622.070 ;
        RECT 2230.700 2608.325 2230.840 2621.750 ;
        RECT 2229.710 2607.955 2229.990 2608.325 ;
        RECT 2230.630 2607.955 2230.910 2608.325 ;
        RECT 2229.780 2560.190 2229.920 2607.955 ;
        RECT 2229.720 2559.870 2229.980 2560.190 ;
        RECT 2231.100 2559.870 2231.360 2560.190 ;
        RECT 2231.160 2511.910 2231.300 2559.870 ;
        RECT 2230.180 2511.765 2230.440 2511.910 ;
        RECT 2228.790 2511.395 2229.070 2511.765 ;
        RECT 2230.170 2511.395 2230.450 2511.765 ;
        RECT 2231.100 2511.590 2231.360 2511.910 ;
        RECT 2228.860 2463.485 2229.000 2511.395 ;
        RECT 2228.790 2463.115 2229.070 2463.485 ;
        RECT 2229.710 2463.115 2229.990 2463.485 ;
        RECT 2229.720 2462.970 2229.980 2463.115 ;
        RECT 2229.720 2428.630 2229.980 2428.950 ;
        RECT 2229.780 2415.090 2229.920 2428.630 ;
        RECT 2229.780 2414.950 2230.380 2415.090 ;
        RECT 2230.240 2380.670 2230.380 2414.950 ;
        RECT 2229.260 2380.410 2229.520 2380.670 ;
        RECT 2229.260 2380.350 2229.920 2380.410 ;
        RECT 2230.180 2380.350 2230.440 2380.670 ;
        RECT 2229.320 2380.270 2229.920 2380.350 ;
        RECT 2229.780 2366.730 2229.920 2380.270 ;
        RECT 2229.720 2366.410 2229.980 2366.730 ;
        RECT 2229.720 2331.730 2229.980 2332.050 ;
        RECT 2229.780 2318.530 2229.920 2331.730 ;
        RECT 2229.780 2318.390 2230.380 2318.530 ;
        RECT 2230.240 2270.365 2230.380 2318.390 ;
        RECT 2228.790 2269.995 2229.070 2270.365 ;
        RECT 2230.170 2269.995 2230.450 2270.365 ;
        RECT 2228.860 2235.830 2229.000 2269.995 ;
        RECT 2228.800 2235.510 2229.060 2235.830 ;
        RECT 2229.260 2235.170 2229.520 2235.490 ;
        RECT 2229.320 2221.890 2229.460 2235.170 ;
        RECT 2227.880 2221.570 2228.140 2221.890 ;
        RECT 2229.260 2221.570 2229.520 2221.890 ;
        RECT 2227.940 2173.805 2228.080 2221.570 ;
        RECT 2227.870 2173.435 2228.150 2173.805 ;
        RECT 2228.790 2173.435 2229.070 2173.805 ;
        RECT 2228.860 2138.330 2229.000 2173.435 ;
        RECT 2228.860 2138.190 2229.460 2138.330 ;
        RECT 2229.320 2125.330 2229.460 2138.190 ;
        RECT 2227.880 2125.010 2228.140 2125.330 ;
        RECT 2229.260 2125.010 2229.520 2125.330 ;
        RECT 2227.940 2077.245 2228.080 2125.010 ;
        RECT 2227.870 2076.875 2228.150 2077.245 ;
        RECT 2228.790 2076.875 2229.070 2077.245 ;
        RECT 2228.860 2042.710 2229.000 2076.875 ;
        RECT 2228.800 2042.390 2229.060 2042.710 ;
        RECT 2229.260 2041.710 2229.520 2042.030 ;
        RECT 2229.320 2021.630 2229.460 2041.710 ;
        RECT 2229.260 2021.310 2229.520 2021.630 ;
        RECT 2229.720 1973.370 2229.980 1973.690 ;
        RECT 2229.780 1932.210 2229.920 1973.370 ;
        RECT 2229.720 1931.890 2229.980 1932.210 ;
        RECT 2229.720 1931.210 2229.980 1931.530 ;
        RECT 2229.780 1897.870 2229.920 1931.210 ;
        RECT 2229.720 1897.550 2229.980 1897.870 ;
        RECT 2229.720 1896.870 2229.980 1897.190 ;
        RECT 2229.780 1849.330 2229.920 1896.870 ;
        RECT 2229.780 1849.190 2230.840 1849.330 ;
        RECT 2230.700 1835.310 2230.840 1849.190 ;
        RECT 2230.640 1834.990 2230.900 1835.310 ;
        RECT 2231.100 1787.050 2231.360 1787.370 ;
        RECT 2231.160 1752.770 2231.300 1787.050 ;
        RECT 2230.240 1752.630 2231.300 1752.770 ;
        RECT 2230.240 1738.750 2230.380 1752.630 ;
        RECT 2230.180 1738.430 2230.440 1738.750 ;
        RECT 1945.430 1700.000 1945.710 1704.000 ;
        RECT 1945.500 1685.370 1945.640 1700.000 ;
        RECT 2231.100 1690.490 2231.360 1690.810 ;
        RECT 2231.160 1685.370 2231.300 1690.490 ;
        RECT 1945.440 1685.050 1945.700 1685.370 ;
        RECT 2231.100 1685.050 2231.360 1685.370 ;
      LAYER via2 ;
        RECT 2231.090 3035.720 2231.370 3036.000 ;
        RECT 2231.090 2959.560 2231.370 2959.840 ;
        RECT 2229.710 2608.000 2229.990 2608.280 ;
        RECT 2230.630 2608.000 2230.910 2608.280 ;
        RECT 2228.790 2511.440 2229.070 2511.720 ;
        RECT 2230.170 2511.440 2230.450 2511.720 ;
        RECT 2228.790 2463.160 2229.070 2463.440 ;
        RECT 2229.710 2463.160 2229.990 2463.440 ;
        RECT 2228.790 2270.040 2229.070 2270.320 ;
        RECT 2230.170 2270.040 2230.450 2270.320 ;
        RECT 2227.870 2173.480 2228.150 2173.760 ;
        RECT 2228.790 2173.480 2229.070 2173.760 ;
        RECT 2227.870 2076.920 2228.150 2077.200 ;
        RECT 2228.790 2076.920 2229.070 2077.200 ;
      LAYER met3 ;
        RECT 2230.350 3036.010 2230.730 3036.020 ;
        RECT 2231.065 3036.010 2231.395 3036.025 ;
        RECT 2230.350 3035.710 2231.395 3036.010 ;
        RECT 2230.350 3035.700 2230.730 3035.710 ;
        RECT 2231.065 3035.695 2231.395 3035.710 ;
        RECT 2230.350 2959.850 2230.730 2959.860 ;
        RECT 2231.065 2959.850 2231.395 2959.865 ;
        RECT 2230.350 2959.550 2231.395 2959.850 ;
        RECT 2230.350 2959.540 2230.730 2959.550 ;
        RECT 2231.065 2959.535 2231.395 2959.550 ;
        RECT 2229.685 2608.290 2230.015 2608.305 ;
        RECT 2230.605 2608.290 2230.935 2608.305 ;
        RECT 2229.685 2607.990 2230.935 2608.290 ;
        RECT 2229.685 2607.975 2230.015 2607.990 ;
        RECT 2230.605 2607.975 2230.935 2607.990 ;
        RECT 2228.765 2511.730 2229.095 2511.745 ;
        RECT 2230.145 2511.730 2230.475 2511.745 ;
        RECT 2228.765 2511.430 2230.475 2511.730 ;
        RECT 2228.765 2511.415 2229.095 2511.430 ;
        RECT 2230.145 2511.415 2230.475 2511.430 ;
        RECT 2228.765 2463.450 2229.095 2463.465 ;
        RECT 2229.685 2463.450 2230.015 2463.465 ;
        RECT 2228.765 2463.150 2230.015 2463.450 ;
        RECT 2228.765 2463.135 2229.095 2463.150 ;
        RECT 2229.685 2463.135 2230.015 2463.150 ;
        RECT 2228.765 2270.330 2229.095 2270.345 ;
        RECT 2230.145 2270.330 2230.475 2270.345 ;
        RECT 2228.765 2270.030 2230.475 2270.330 ;
        RECT 2228.765 2270.015 2229.095 2270.030 ;
        RECT 2230.145 2270.015 2230.475 2270.030 ;
        RECT 2227.845 2173.770 2228.175 2173.785 ;
        RECT 2228.765 2173.770 2229.095 2173.785 ;
        RECT 2227.845 2173.470 2229.095 2173.770 ;
        RECT 2227.845 2173.455 2228.175 2173.470 ;
        RECT 2228.765 2173.455 2229.095 2173.470 ;
        RECT 2227.845 2077.210 2228.175 2077.225 ;
        RECT 2228.765 2077.210 2229.095 2077.225 ;
        RECT 2227.845 2076.910 2229.095 2077.210 ;
        RECT 2227.845 2076.895 2228.175 2076.910 ;
        RECT 2228.765 2076.895 2229.095 2076.910 ;
      LAYER via3 ;
        RECT 2230.380 3035.700 2230.700 3036.020 ;
        RECT 2230.380 2959.540 2230.700 2959.860 ;
      LAYER met4 ;
<<<<<<< HEAD
        RECT 1945.175 3502.175 1945.505 3502.505 ;
        RECT 1945.190 1702.545 1945.490 3502.175 ;
        RECT 1945.175 1702.215 1945.505 1702.545 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2230.375 3035.695 2230.705 3036.025 ;
        RECT 2230.390 2959.865 2230.690 3035.695 ;
        RECT 2230.375 2959.535 2230.705 2959.865 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1905.850 3501.900 1906.170 3501.960 ;
        RECT 1946.790 3501.900 1947.110 3501.960 ;
        RECT 1905.850 3501.760 1947.110 3501.900 ;
        RECT 1905.850 3501.700 1906.170 3501.760 ;
        RECT 1946.790 3501.700 1947.110 3501.760 ;
      LAYER via ;
        RECT 1905.880 3501.700 1906.140 3501.960 ;
        RECT 1946.820 3501.700 1947.080 3501.960 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1905.730 3519.700 1906.290 3524.800 ;
=======
        RECT 1905.730 3517.600 1906.290 3524.800 ;
<<<<<<< HEAD
        RECT 1905.940 3502.330 1906.080 3517.600 ;
        RECT 1905.880 3502.010 1906.140 3502.330 ;
        RECT 1946.820 3502.010 1947.080 3502.330 ;
        RECT 1946.880 1703.810 1947.020 3502.010 ;
        RECT 1947.270 1703.810 1947.550 1704.000 ;
        RECT 1946.880 1703.670 1947.550 1703.810 ;
        RECT 1947.270 1700.000 1947.550 1703.670 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1905.940 3501.990 1906.080 3517.600 ;
        RECT 1905.880 3501.670 1906.140 3501.990 ;
        RECT 1946.820 3501.670 1947.080 3501.990 ;
        RECT 1946.880 1704.000 1947.020 3501.670 ;
        RECT 1946.810 1700.000 1947.090 1704.000 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1581.550 3483.880 1581.870 3483.940 ;
        RECT 1586.610 3483.880 1586.930 3483.940 ;
        RECT 1581.550 3483.740 1586.930 3483.880 ;
        RECT 1581.550 3483.680 1581.870 3483.740 ;
        RECT 1586.610 3483.680 1586.930 3483.740 ;
        RECT 1586.610 3073.840 1586.930 3073.900 ;
        RECT 1952.770 3073.840 1953.090 3073.900 ;
        RECT 1586.610 3073.700 1953.090 3073.840 ;
        RECT 1586.610 3073.640 1586.930 3073.700 ;
        RECT 1952.770 3073.640 1953.090 3073.700 ;
      LAYER via ;
        RECT 1581.580 3483.680 1581.840 3483.940 ;
        RECT 1586.640 3483.680 1586.900 3483.940 ;
        RECT 1586.640 3073.640 1586.900 3073.900 ;
        RECT 1952.800 3073.640 1953.060 3073.900 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1581.430 3519.700 1581.990 3524.800 ;
=======
        RECT 1581.430 3517.600 1581.990 3524.800 ;
        RECT 1581.640 3483.970 1581.780 3517.600 ;
        RECT 1581.580 3483.650 1581.840 3483.970 ;
        RECT 1586.640 3483.650 1586.900 3483.970 ;
        RECT 1586.700 3073.930 1586.840 3483.650 ;
        RECT 1586.640 3073.610 1586.900 3073.930 ;
        RECT 1952.800 3073.610 1953.060 3073.930 ;
        RECT 1952.860 2300.285 1953.000 3073.610 ;
        RECT 1952.790 2299.915 1953.070 2300.285 ;
      LAYER via2 ;
        RECT 1952.790 2299.960 1953.070 2300.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1138.105 2059.530 1138.435 2059.545 ;
        RECT 1150.000 2059.530 1154.000 2059.680 ;
        RECT 1138.105 2059.230 1154.000 2059.530 ;
        RECT 1138.105 2059.215 1138.435 2059.230 ;
        RECT 1150.000 2059.080 1154.000 2059.230 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1946.000 2300.250 1950.000 2300.400 ;
        RECT 1952.765 2300.250 1953.095 2300.265 ;
        RECT 1946.000 2299.950 1953.095 2300.250 ;
        RECT 1946.000 2299.800 1950.000 2299.950 ;
        RECT 1952.765 2299.935 1953.095 2299.950 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1137.650 268.840 1137.970 268.900 ;
        RECT 2900.830 268.840 2901.150 268.900 ;
        RECT 1137.650 268.700 2901.150 268.840 ;
        RECT 1137.650 268.640 1137.970 268.700 ;
        RECT 2900.830 268.640 2901.150 268.700 ;
      LAYER via ;
        RECT 1137.680 268.640 1137.940 268.900 ;
        RECT 2900.860 268.640 2901.120 268.900 ;
      LAYER met2 ;
        RECT 1137.670 1832.755 1137.950 1833.125 ;
        RECT 1137.740 268.930 1137.880 1832.755 ;
        RECT 1137.680 268.610 1137.940 268.930 ;
        RECT 2900.860 268.610 2901.120 268.930 ;
        RECT 2900.920 264.365 2901.060 268.610 ;
        RECT 2900.850 263.995 2901.130 264.365 ;
      LAYER via2 ;
        RECT 1137.670 1832.800 1137.950 1833.080 ;
        RECT 2900.850 264.040 2901.130 264.320 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 263.580 2924.800 264.780 ;
=======
        RECT 1138.105 1739.930 1138.435 1739.945 ;
        RECT 1150.000 1739.930 1154.000 1740.080 ;
        RECT 1138.105 1739.630 1154.000 1739.930 ;
        RECT 1138.105 1739.615 1138.435 1739.630 ;
        RECT 1150.000 1739.480 1154.000 1739.630 ;
=======
        RECT 1137.645 1833.090 1137.975 1833.105 ;
        RECT 1150.000 1833.090 1154.000 1833.240 ;
        RECT 1137.645 1832.790 1154.000 1833.090 ;
        RECT 1137.645 1832.775 1137.975 1832.790 ;
        RECT 1150.000 1832.640 1154.000 1832.790 ;
>>>>>>> re-updated local openlane
        RECT 2900.825 264.330 2901.155 264.345 ;
        RECT 2917.600 264.330 2924.800 264.780 ;
        RECT 2900.825 264.030 2924.800 264.330 ;
        RECT 2900.825 264.015 2901.155 264.030 ;
        RECT 2917.600 263.580 2924.800 264.030 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1257.250 3498.500 1257.570 3498.560 ;
        RECT 1262.310 3498.500 1262.630 3498.560 ;
        RECT 1257.250 3498.360 1262.630 3498.500 ;
        RECT 1257.250 3498.300 1257.570 3498.360 ;
        RECT 1262.310 3498.300 1262.630 3498.360 ;
        RECT 1262.310 2516.920 1262.630 2516.980 ;
        RECT 1920.570 2516.920 1920.890 2516.980 ;
        RECT 1262.310 2516.780 1920.890 2516.920 ;
        RECT 1262.310 2516.720 1262.630 2516.780 ;
        RECT 1920.570 2516.720 1920.890 2516.780 ;
      LAYER via ;
        RECT 1257.280 3498.300 1257.540 3498.560 ;
        RECT 1262.340 3498.300 1262.600 3498.560 ;
        RECT 1262.340 2516.720 1262.600 2516.980 ;
        RECT 1920.600 2516.720 1920.860 2516.980 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1257.130 3519.700 1257.690 3524.800 ;
=======
        RECT 1257.130 3517.600 1257.690 3524.800 ;
        RECT 1257.340 3498.590 1257.480 3517.600 ;
        RECT 1257.280 3498.270 1257.540 3498.590 ;
        RECT 1262.340 3498.270 1262.600 3498.590 ;
<<<<<<< HEAD
        RECT 1262.400 2509.190 1262.540 3498.270 ;
        RECT 1262.340 2508.870 1262.600 2509.190 ;
        RECT 1959.700 2496.290 1959.960 2496.610 ;
        RECT 1959.760 2167.005 1959.900 2496.290 ;
        RECT 1959.690 2166.635 1959.970 2167.005 ;
      LAYER via2 ;
        RECT 1959.690 2166.680 1959.970 2166.960 ;
      LAYER met3 ;
        RECT 1946.000 2166.970 1950.000 2167.120 ;
        RECT 1959.665 2166.970 1959.995 2166.985 ;
        RECT 1946.000 2166.670 1959.995 2166.970 ;
        RECT 1946.000 2166.520 1950.000 2166.670 ;
        RECT 1959.665 2166.655 1959.995 2166.670 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1262.400 2517.010 1262.540 3498.270 ;
        RECT 1262.340 2516.690 1262.600 2517.010 ;
        RECT 1920.600 2516.690 1920.860 2517.010 ;
        RECT 1920.660 2500.000 1920.800 2516.690 ;
        RECT 1920.590 2496.000 1920.870 2500.000 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.490 3498.500 932.810 3498.560 ;
        RECT 938.010 3498.500 938.330 3498.560 ;
        RECT 932.490 3498.360 938.330 3498.500 ;
        RECT 932.490 3498.300 932.810 3498.360 ;
        RECT 938.010 3498.300 938.330 3498.360 ;
        RECT 938.010 2194.260 938.330 2194.320 ;
        RECT 1131.670 2194.260 1131.990 2194.320 ;
        RECT 938.010 2194.120 1131.990 2194.260 ;
        RECT 938.010 2194.060 938.330 2194.120 ;
        RECT 1131.670 2194.060 1131.990 2194.120 ;
      LAYER via ;
        RECT 932.520 3498.300 932.780 3498.560 ;
        RECT 938.040 3498.300 938.300 3498.560 ;
        RECT 938.040 2194.060 938.300 2194.320 ;
        RECT 1131.700 2194.060 1131.960 2194.320 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 932.370 3519.700 932.930 3524.800 ;
=======
        RECT 932.370 3517.600 932.930 3524.800 ;
        RECT 932.580 3498.590 932.720 3517.600 ;
        RECT 932.520 3498.270 932.780 3498.590 ;
        RECT 938.040 3498.270 938.300 3498.590 ;
<<<<<<< HEAD
        RECT 938.100 1696.930 938.240 3498.270 ;
        RECT 1948.650 1700.000 1948.930 1704.000 ;
        RECT 1948.720 1696.930 1948.860 1700.000 ;
        RECT 938.040 1696.610 938.300 1696.930 ;
        RECT 1948.660 1696.610 1948.920 1696.930 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 938.100 2194.350 938.240 3498.270 ;
        RECT 938.040 2194.030 938.300 2194.350 ;
        RECT 1131.700 2194.030 1131.960 2194.350 ;
        RECT 1131.760 2188.765 1131.900 2194.030 ;
        RECT 1131.690 2188.395 1131.970 2188.765 ;
      LAYER via2 ;
        RECT 1131.690 2188.440 1131.970 2188.720 ;
      LAYER met3 ;
        RECT 1131.665 2188.730 1131.995 2188.745 ;
        RECT 1150.000 2188.730 1154.000 2188.880 ;
        RECT 1131.665 2188.430 1154.000 2188.730 ;
        RECT 1131.665 2188.415 1131.995 2188.430 ;
        RECT 1150.000 2188.280 1154.000 2188.430 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 608.190 3498.500 608.510 3498.560 ;
        RECT 613.710 3498.500 614.030 3498.560 ;
        RECT 608.190 3498.360 614.030 3498.500 ;
        RECT 608.190 3498.300 608.510 3498.360 ;
        RECT 613.710 3498.300 614.030 3498.360 ;
        RECT 613.710 2283.680 614.030 2283.740 ;
        RECT 1131.670 2283.680 1131.990 2283.740 ;
        RECT 613.710 2283.540 1131.990 2283.680 ;
        RECT 613.710 2283.480 614.030 2283.540 ;
        RECT 1131.670 2283.480 1131.990 2283.540 ;
      LAYER via ;
        RECT 608.220 3498.300 608.480 3498.560 ;
        RECT 613.740 3498.300 614.000 3498.560 ;
        RECT 613.740 2283.480 614.000 2283.740 ;
        RECT 1131.700 2283.480 1131.960 2283.740 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 608.070 3519.700 608.630 3524.800 ;
=======
        RECT 608.070 3517.600 608.630 3524.800 ;
        RECT 608.280 3498.590 608.420 3517.600 ;
        RECT 608.220 3498.270 608.480 3498.590 ;
        RECT 613.740 3498.270 614.000 3498.590 ;
<<<<<<< HEAD
        RECT 613.800 2522.110 613.940 3498.270 ;
        RECT 613.740 2521.790 614.000 2522.110 ;
        RECT 1939.920 2521.790 1940.180 2522.110 ;
        RECT 1939.980 2500.000 1940.120 2521.790 ;
        RECT 1939.910 2496.000 1940.190 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 613.800 2283.770 613.940 3498.270 ;
        RECT 613.740 2283.450 614.000 2283.770 ;
        RECT 1131.700 2283.450 1131.960 2283.770 ;
        RECT 1131.760 2277.845 1131.900 2283.450 ;
        RECT 1131.690 2277.475 1131.970 2277.845 ;
      LAYER via2 ;
        RECT 1131.690 2277.520 1131.970 2277.800 ;
      LAYER met3 ;
        RECT 1131.665 2277.810 1131.995 2277.825 ;
        RECT 1150.000 2277.810 1154.000 2277.960 ;
        RECT 1131.665 2277.510 1154.000 2277.810 ;
        RECT 1131.665 2277.495 1131.995 2277.510 ;
        RECT 1150.000 2277.360 1154.000 2277.510 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 283.890 3500.880 284.210 3500.940 ;
        RECT 289.410 3500.880 289.730 3500.940 ;
        RECT 283.890 3500.740 289.730 3500.880 ;
        RECT 283.890 3500.680 284.210 3500.740 ;
        RECT 289.410 3500.680 289.730 3500.740 ;
        RECT 289.410 2501.280 289.730 2501.340 ;
        RECT 1959.670 2501.280 1959.990 2501.340 ;
        RECT 289.410 2501.140 1959.990 2501.280 ;
        RECT 289.410 2501.080 289.730 2501.140 ;
        RECT 1959.670 2501.080 1959.990 2501.140 ;
      LAYER via ;
        RECT 283.920 3500.680 284.180 3500.940 ;
        RECT 289.440 3500.680 289.700 3500.940 ;
        RECT 289.440 2501.080 289.700 2501.340 ;
        RECT 1959.700 2501.080 1959.960 2501.340 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 283.770 3519.700 284.330 3524.800 ;
=======
        RECT 283.770 3517.600 284.330 3524.800 ;
        RECT 283.980 3500.970 284.120 3517.600 ;
        RECT 283.920 3500.650 284.180 3500.970 ;
        RECT 289.440 3500.650 289.700 3500.970 ;
        RECT 289.500 2501.370 289.640 3500.650 ;
        RECT 289.440 2501.050 289.700 2501.370 ;
        RECT 1959.700 2501.050 1959.960 2501.370 ;
        RECT 1959.760 2433.565 1959.900 2501.050 ;
        RECT 1959.690 2433.195 1959.970 2433.565 ;
      LAYER via2 ;
        RECT 1959.690 2433.240 1959.970 2433.520 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1131.665 2139.770 1131.995 2139.785 ;
        RECT 1150.000 2139.770 1154.000 2139.920 ;
        RECT 1131.665 2139.470 1154.000 2139.770 ;
        RECT 1131.665 2139.455 1131.995 2139.470 ;
        RECT 1150.000 2139.320 1154.000 2139.470 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1946.000 2433.530 1950.000 2433.680 ;
        RECT 1959.665 2433.530 1959.995 2433.545 ;
        RECT 1946.000 2433.230 1959.995 2433.530 ;
        RECT 1946.000 2433.080 1950.000 2433.230 ;
        RECT 1959.665 2433.215 1959.995 2433.230 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3477.760 17.410 3477.820 ;
        RECT 51.590 3477.760 51.910 3477.820 ;
        RECT 17.090 3477.620 51.910 3477.760 ;
        RECT 17.090 3477.560 17.410 3477.620 ;
        RECT 51.590 3477.560 51.910 3477.620 ;
        RECT 51.590 2366.640 51.910 2366.700 ;
        RECT 1131.670 2366.640 1131.990 2366.700 ;
        RECT 51.590 2366.500 1131.990 2366.640 ;
        RECT 51.590 2366.440 51.910 2366.500 ;
        RECT 1131.670 2366.440 1131.990 2366.500 ;
      LAYER via ;
        RECT 17.120 3477.560 17.380 3477.820 ;
        RECT 51.620 3477.560 51.880 3477.820 ;
        RECT 51.620 2366.440 51.880 2366.700 ;
        RECT 1131.700 2366.440 1131.960 2366.700 ;
      LAYER met2 ;
        RECT 17.110 3483.115 17.390 3483.485 ;
        RECT 17.180 3477.850 17.320 3483.115 ;
        RECT 17.120 3477.530 17.380 3477.850 ;
        RECT 51.620 3477.530 51.880 3477.850 ;
        RECT 51.680 2366.730 51.820 3477.530 ;
        RECT 51.620 2366.410 51.880 2366.730 ;
        RECT 1131.700 2366.410 1131.960 2366.730 ;
        RECT 1131.760 2366.245 1131.900 2366.410 ;
        RECT 1131.690 2365.875 1131.970 2366.245 ;
      LAYER via2 ;
        RECT 17.110 3483.160 17.390 3483.440 ;
        RECT 1131.690 2365.920 1131.970 2366.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3482.700 0.300 3483.900 ;
=======
        RECT -4.800 3483.450 2.400 3483.900 ;
        RECT 17.085 3483.450 17.415 3483.465 ;
        RECT -4.800 3483.150 17.415 3483.450 ;
        RECT -4.800 3482.700 2.400 3483.150 ;
        RECT 17.085 3483.135 17.415 3483.150 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1131.665 2366.210 1131.995 2366.225 ;
        RECT 1150.000 2366.210 1154.000 2366.360 ;
        RECT 1131.665 2365.910 1154.000 2366.210 ;
        RECT 1131.665 2365.895 1131.995 2365.910 ;
        RECT 1150.000 2365.760 1154.000 2365.910 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2515.560 17.410 2515.620 ;
        RECT 1927.010 2515.560 1927.330 2515.620 ;
        RECT 17.090 2515.420 1927.330 2515.560 ;
        RECT 17.090 2515.360 17.410 2515.420 ;
        RECT 1927.010 2515.360 1927.330 2515.420 ;
      LAYER via ;
        RECT 17.120 2515.360 17.380 2515.620 ;
        RECT 1927.040 2515.360 1927.300 2515.620 ;
      LAYER met2 ;
        RECT 17.110 3195.475 17.390 3195.845 ;
        RECT 17.180 2515.650 17.320 3195.475 ;
        RECT 17.120 2515.330 17.380 2515.650 ;
        RECT 1927.040 2515.330 1927.300 2515.650 ;
        RECT 1927.100 2500.000 1927.240 2515.330 ;
        RECT 1927.030 2496.000 1927.310 2500.000 ;
      LAYER via2 ;
        RECT 17.110 3195.520 17.390 3195.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3195.060 0.300 3196.260 ;
=======
        RECT -4.800 3195.810 2.400 3196.260 ;
        RECT 17.085 3195.810 17.415 3195.825 ;
        RECT -4.800 3195.510 17.415 3195.810 ;
        RECT -4.800 3195.060 2.400 3195.510 ;
        RECT 17.085 3195.495 17.415 3195.510 ;
<<<<<<< HEAD
        RECT 1947.245 2302.290 1947.575 2302.305 ;
        RECT 1947.030 2301.975 1947.575 2302.290 ;
        RECT 1947.030 2300.400 1947.330 2301.975 ;
        RECT 1946.000 2299.800 1950.000 2300.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2515.220 17.870 2515.280 ;
        RECT 1933.450 2515.220 1933.770 2515.280 ;
        RECT 17.550 2515.080 1933.770 2515.220 ;
        RECT 17.550 2515.020 17.870 2515.080 ;
        RECT 1933.450 2515.020 1933.770 2515.080 ;
      LAYER via ;
        RECT 17.580 2515.020 17.840 2515.280 ;
        RECT 1933.480 2515.020 1933.740 2515.280 ;
      LAYER met2 ;
        RECT 17.570 2908.515 17.850 2908.885 ;
        RECT 17.640 2515.310 17.780 2908.515 ;
        RECT 17.580 2514.990 17.840 2515.310 ;
        RECT 1933.480 2514.990 1933.740 2515.310 ;
        RECT 1933.540 2500.000 1933.680 2514.990 ;
        RECT 1933.470 2496.000 1933.750 2500.000 ;
      LAYER via2 ;
        RECT 17.570 2908.560 17.850 2908.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2908.100 0.300 2909.300 ;
=======
        RECT -4.800 2908.850 2.400 2909.300 ;
        RECT 17.545 2908.850 17.875 2908.865 ;
        RECT -4.800 2908.550 17.875 2908.850 ;
        RECT -4.800 2908.100 2.400 2908.550 ;
<<<<<<< HEAD
        RECT 17.085 2908.535 17.415 2908.550 ;
        RECT 1131.665 2219.330 1131.995 2219.345 ;
        RECT 1150.000 2219.330 1154.000 2219.480 ;
        RECT 1131.665 2219.030 1154.000 2219.330 ;
        RECT 1131.665 2219.015 1131.995 2219.030 ;
        RECT 1150.000 2218.880 1154.000 2219.030 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 17.545 2908.535 17.875 2908.550 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 2514.880 18.330 2514.940 ;
        RECT 1939.890 2514.880 1940.210 2514.940 ;
        RECT 18.010 2514.740 1940.210 2514.880 ;
        RECT 18.010 2514.680 18.330 2514.740 ;
        RECT 1939.890 2514.680 1940.210 2514.740 ;
      LAYER via ;
        RECT 18.040 2514.680 18.300 2514.940 ;
        RECT 1939.920 2514.680 1940.180 2514.940 ;
      LAYER met2 ;
        RECT 18.030 2620.875 18.310 2621.245 ;
        RECT 18.100 2514.970 18.240 2620.875 ;
        RECT 18.040 2514.650 18.300 2514.970 ;
        RECT 1939.920 2514.650 1940.180 2514.970 ;
        RECT 1939.980 2500.000 1940.120 2514.650 ;
        RECT 1939.910 2496.000 1940.190 2500.000 ;
      LAYER via2 ;
        RECT 18.030 2620.920 18.310 2621.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2620.460 0.300 2621.660 ;
=======
        RECT -4.800 2621.210 2.400 2621.660 ;
        RECT 18.005 2621.210 18.335 2621.225 ;
        RECT -4.800 2620.910 18.335 2621.210 ;
        RECT -4.800 2620.460 2.400 2620.910 ;
<<<<<<< HEAD
        RECT 16.165 2620.895 16.495 2620.910 ;
        RECT 1131.665 2299.570 1131.995 2299.585 ;
        RECT 1150.000 2299.570 1154.000 2299.720 ;
        RECT 1131.665 2299.270 1154.000 2299.570 ;
        RECT 1131.665 2299.255 1131.995 2299.270 ;
        RECT 1150.000 2299.120 1154.000 2299.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 18.005 2620.895 18.335 2620.910 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 65.850 2449.600 66.170 2449.660 ;
        RECT 1131.670 2449.600 1131.990 2449.660 ;
        RECT 65.850 2449.460 1131.990 2449.600 ;
        RECT 65.850 2449.400 66.170 2449.460 ;
        RECT 1131.670 2449.400 1131.990 2449.460 ;
        RECT 16.630 2339.100 16.950 2339.160 ;
        RECT 65.850 2339.100 66.170 2339.160 ;
        RECT 16.630 2338.960 66.170 2339.100 ;
        RECT 16.630 2338.900 16.950 2338.960 ;
        RECT 65.850 2338.900 66.170 2338.960 ;
      LAYER via ;
        RECT 65.880 2449.400 66.140 2449.660 ;
        RECT 1131.700 2449.400 1131.960 2449.660 ;
        RECT 16.660 2338.900 16.920 2339.160 ;
        RECT 65.880 2338.900 66.140 2339.160 ;
      LAYER met2 ;
        RECT 1131.690 2454.955 1131.970 2455.325 ;
        RECT 1131.760 2449.690 1131.900 2454.955 ;
        RECT 65.880 2449.370 66.140 2449.690 ;
        RECT 1131.700 2449.370 1131.960 2449.690 ;
        RECT 65.940 2339.190 66.080 2449.370 ;
        RECT 16.660 2338.870 16.920 2339.190 ;
        RECT 65.880 2338.870 66.140 2339.190 ;
        RECT 16.720 2334.285 16.860 2338.870 ;
        RECT 16.650 2333.915 16.930 2334.285 ;
      LAYER via2 ;
        RECT 1131.690 2455.000 1131.970 2455.280 ;
        RECT 16.650 2333.960 16.930 2334.240 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT -4.800 2333.500 0.300 2334.700 ;
=======
        RECT 1946.000 2433.530 1950.000 2433.680 ;
        RECT 1959.870 2433.530 1960.250 2433.540 ;
        RECT 1946.000 2433.230 1960.250 2433.530 ;
        RECT 1946.000 2433.080 1950.000 2433.230 ;
        RECT 1959.870 2433.220 1960.250 2433.230 ;
        RECT 290.070 2341.050 290.450 2341.060 ;
        RECT 336.990 2341.050 337.370 2341.060 ;
        RECT 290.070 2340.750 337.370 2341.050 ;
        RECT 290.070 2340.740 290.450 2340.750 ;
        RECT 336.990 2340.740 337.370 2340.750 ;
        RECT 386.670 2341.050 387.050 2341.060 ;
        RECT 433.590 2341.050 433.970 2341.060 ;
        RECT 386.670 2340.750 433.970 2341.050 ;
        RECT 386.670 2340.740 387.050 2340.750 ;
        RECT 433.590 2340.740 433.970 2340.750 ;
        RECT 483.270 2341.050 483.650 2341.060 ;
        RECT 530.190 2341.050 530.570 2341.060 ;
        RECT 483.270 2340.750 530.570 2341.050 ;
        RECT 483.270 2340.740 483.650 2340.750 ;
        RECT 530.190 2340.740 530.570 2340.750 ;
        RECT 773.070 2341.050 773.450 2341.060 ;
        RECT 819.990 2341.050 820.370 2341.060 ;
        RECT 773.070 2340.750 820.370 2341.050 ;
        RECT 773.070 2340.740 773.450 2340.750 ;
        RECT 819.990 2340.740 820.370 2340.750 ;
        RECT 966.270 2341.050 966.650 2341.060 ;
        RECT 980.990 2341.050 981.370 2341.060 ;
        RECT 966.270 2340.750 981.370 2341.050 ;
        RECT 966.270 2340.740 966.650 2340.750 ;
        RECT 980.990 2340.740 981.370 2340.750 ;
        RECT 1062.870 2341.050 1063.250 2341.060 ;
        RECT 1109.790 2341.050 1110.170 2341.060 ;
        RECT 1062.870 2340.750 1110.170 2341.050 ;
        RECT 1062.870 2340.740 1063.250 2340.750 ;
        RECT 1109.790 2340.740 1110.170 2340.750 ;
=======
        RECT 1131.665 2455.290 1131.995 2455.305 ;
        RECT 1150.000 2455.290 1154.000 2455.440 ;
        RECT 1131.665 2454.990 1154.000 2455.290 ;
        RECT 1131.665 2454.975 1131.995 2454.990 ;
        RECT 1150.000 2454.840 1154.000 2454.990 ;
>>>>>>> re-updated local openlane
        RECT -4.800 2334.250 2.400 2334.700 ;
        RECT 16.625 2334.250 16.955 2334.265 ;
        RECT -4.800 2333.950 16.955 2334.250 ;
        RECT -4.800 2333.500 2.400 2333.950 ;
<<<<<<< HEAD
        RECT 26.030 2333.940 26.410 2333.950 ;
      LAYER via3 ;
        RECT 1959.900 2433.220 1960.220 2433.540 ;
        RECT 290.100 2340.740 290.420 2341.060 ;
        RECT 337.020 2340.740 337.340 2341.060 ;
        RECT 386.700 2340.740 387.020 2341.060 ;
        RECT 433.620 2340.740 433.940 2341.060 ;
        RECT 483.300 2340.740 483.620 2341.060 ;
        RECT 530.220 2340.740 530.540 2341.060 ;
        RECT 773.100 2340.740 773.420 2341.060 ;
        RECT 820.020 2340.740 820.340 2341.060 ;
        RECT 966.300 2340.740 966.620 2341.060 ;
        RECT 981.020 2340.740 981.340 2341.060 ;
        RECT 1062.900 2340.740 1063.220 2341.060 ;
        RECT 1109.820 2340.740 1110.140 2341.060 ;
        RECT 26.060 2333.940 26.380 2334.260 ;
      LAYER met4 ;
        RECT 1959.895 2433.215 1960.225 2433.545 ;
        RECT 289.670 2340.310 290.850 2341.490 ;
        RECT 336.590 2340.310 337.770 2341.490 ;
        RECT 386.270 2340.310 387.450 2341.490 ;
        RECT 433.190 2340.310 434.370 2341.490 ;
        RECT 482.870 2340.310 484.050 2341.490 ;
        RECT 529.790 2340.310 530.970 2341.490 ;
        RECT 772.670 2340.310 773.850 2341.490 ;
        RECT 820.015 2340.735 820.345 2341.065 ;
        RECT 820.030 2334.690 820.330 2340.735 ;
        RECT 965.870 2340.310 967.050 2341.490 ;
        RECT 980.590 2340.310 981.770 2341.490 ;
        RECT 1062.470 2340.310 1063.650 2341.490 ;
        RECT 1109.815 2340.735 1110.145 2341.065 ;
        RECT 1109.830 2334.690 1110.130 2340.735 ;
        RECT 1159.990 2340.310 1161.170 2341.490 ;
        RECT 1182.990 2340.310 1184.170 2341.490 ;
        RECT 25.630 2333.510 26.810 2334.690 ;
        RECT 819.590 2333.510 820.770 2334.690 ;
        RECT 1109.390 2333.510 1110.570 2334.690 ;
        RECT 1160.430 2327.890 1160.730 2340.310 ;
        RECT 1183.430 2327.890 1183.730 2340.310 ;
        RECT 1959.910 2334.690 1960.210 2433.215 ;
        RECT 1959.470 2333.510 1960.650 2334.690 ;
        RECT 1159.990 2326.710 1161.170 2327.890 ;
        RECT 1182.990 2326.710 1184.170 2327.890 ;
      LAYER met5 ;
        RECT 59.460 2340.100 97.860 2341.700 ;
        RECT 59.460 2334.900 61.060 2340.100 ;
        RECT 25.420 2333.300 61.060 2334.900 ;
        RECT 96.260 2334.900 97.860 2340.100 ;
        RECT 143.180 2340.100 194.460 2341.700 ;
        RECT 143.180 2334.900 144.780 2340.100 ;
        RECT 96.260 2333.300 144.780 2334.900 ;
        RECT 192.860 2334.900 194.460 2340.100 ;
        RECT 239.780 2340.100 291.060 2341.700 ;
        RECT 336.380 2340.100 387.660 2341.700 ;
        RECT 432.980 2340.100 484.260 2341.700 ;
        RECT 529.580 2340.100 580.860 2341.700 ;
        RECT 239.780 2334.900 241.380 2340.100 ;
        RECT 192.860 2333.300 241.380 2334.900 ;
        RECT 579.260 2334.900 580.860 2340.100 ;
        RECT 626.180 2340.100 677.460 2341.700 ;
        RECT 626.180 2334.900 627.780 2340.100 ;
        RECT 579.260 2333.300 627.780 2334.900 ;
        RECT 675.860 2334.900 677.460 2340.100 ;
        RECT 722.780 2340.100 774.060 2341.700 ;
        RECT 833.180 2340.100 871.580 2341.700 ;
        RECT 722.780 2334.900 724.380 2340.100 ;
        RECT 833.180 2334.900 834.780 2340.100 ;
        RECT 675.860 2333.300 724.380 2334.900 ;
        RECT 819.380 2333.300 834.780 2334.900 ;
        RECT 869.980 2328.100 871.580 2340.100 ;
        RECT 929.780 2340.100 967.260 2341.700 ;
        RECT 980.380 2340.100 1014.180 2341.700 ;
        RECT 929.780 2334.900 931.380 2340.100 ;
        RECT 915.980 2333.300 931.380 2334.900 ;
        RECT 1012.580 2334.900 1014.180 2340.100 ;
        RECT 1026.380 2340.100 1063.860 2341.700 ;
        RECT 1122.980 2340.100 1161.380 2341.700 ;
        RECT 1182.780 2340.100 1207.380 2341.700 ;
        RECT 1026.380 2334.900 1027.980 2340.100 ;
        RECT 1122.980 2334.900 1124.580 2340.100 ;
        RECT 1205.780 2338.300 1207.380 2340.100 ;
        RECT 1217.740 2340.100 1257.060 2341.700 ;
        RECT 1217.740 2338.300 1219.340 2340.100 ;
        RECT 1205.780 2336.700 1219.340 2338.300 ;
        RECT 1255.460 2338.300 1257.060 2340.100 ;
        RECT 1316.180 2340.100 1354.580 2341.700 ;
        RECT 1255.460 2336.700 1303.980 2338.300 ;
        RECT 1012.580 2333.300 1027.980 2334.900 ;
        RECT 1109.180 2333.300 1124.580 2334.900 ;
        RECT 1302.380 2334.900 1303.980 2336.700 ;
        RECT 1316.180 2334.900 1317.780 2340.100 ;
        RECT 1302.380 2333.300 1317.780 2334.900 ;
        RECT 915.980 2328.100 917.580 2333.300 ;
        RECT 1352.980 2328.100 1354.580 2340.100 ;
        RECT 1412.780 2340.100 1451.180 2341.700 ;
        RECT 1412.780 2334.900 1414.380 2340.100 ;
        RECT 1398.980 2333.300 1414.380 2334.900 ;
        RECT 1398.980 2328.100 1400.580 2333.300 ;
        RECT 869.980 2326.500 917.580 2328.100 ;
        RECT 1159.780 2326.500 1184.380 2328.100 ;
        RECT 1352.980 2326.500 1400.580 2328.100 ;
        RECT 1449.580 2328.100 1451.180 2340.100 ;
        RECT 1509.380 2340.100 1547.780 2341.700 ;
        RECT 1509.380 2334.900 1510.980 2340.100 ;
        RECT 1495.580 2333.300 1510.980 2334.900 ;
        RECT 1495.580 2328.100 1497.180 2333.300 ;
        RECT 1449.580 2326.500 1497.180 2328.100 ;
        RECT 1546.180 2328.100 1547.780 2340.100 ;
        RECT 1605.980 2340.100 1644.380 2341.700 ;
        RECT 1605.980 2334.900 1607.580 2340.100 ;
        RECT 1592.180 2333.300 1607.580 2334.900 ;
        RECT 1592.180 2328.100 1593.780 2333.300 ;
        RECT 1546.180 2326.500 1593.780 2328.100 ;
        RECT 1642.780 2328.100 1644.380 2340.100 ;
        RECT 1702.580 2340.100 1740.980 2341.700 ;
        RECT 1702.580 2334.900 1704.180 2340.100 ;
        RECT 1688.780 2333.300 1704.180 2334.900 ;
        RECT 1688.780 2328.100 1690.380 2333.300 ;
        RECT 1642.780 2326.500 1690.380 2328.100 ;
        RECT 1739.380 2328.100 1740.980 2340.100 ;
        RECT 1799.180 2340.100 1837.580 2341.700 ;
        RECT 1799.180 2334.900 1800.780 2340.100 ;
        RECT 1785.380 2333.300 1800.780 2334.900 ;
        RECT 1785.380 2328.100 1786.980 2333.300 ;
        RECT 1739.380 2326.500 1786.980 2328.100 ;
        RECT 1835.980 2328.100 1837.580 2340.100 ;
        RECT 1895.780 2340.100 1933.260 2341.700 ;
        RECT 1895.780 2334.900 1897.380 2340.100 ;
        RECT 1881.980 2333.300 1897.380 2334.900 ;
        RECT 1931.660 2334.900 1933.260 2340.100 ;
        RECT 1931.660 2333.300 1960.860 2334.900 ;
        RECT 1881.980 2328.100 1883.580 2333.300 ;
        RECT 1835.980 2326.500 1883.580 2328.100 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 2333.935 16.955 2333.950 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 48.445 1684.445 48.615 1685.295 ;
        RECT 96.285 1684.445 96.455 1685.635 ;
        RECT 110.545 1685.465 111.175 1685.635 ;
        RECT 158.845 1684.105 159.015 1684.955 ;
        RECT 193.345 1683.425 193.515 1684.275 ;
        RECT 241.185 1683.425 241.355 1684.615 ;
        RECT 255.445 1684.105 255.615 1684.955 ;
        RECT 289.945 1683.425 290.115 1684.275 ;
        RECT 337.785 1683.425 337.955 1684.615 ;
        RECT 352.045 1684.105 352.215 1684.955 ;
        RECT 386.545 1683.425 386.715 1684.275 ;
        RECT 434.385 1683.425 434.555 1684.615 ;
        RECT 448.645 1684.105 448.815 1684.955 ;
        RECT 483.145 1683.425 483.315 1684.275 ;
        RECT 530.985 1683.425 531.155 1684.615 ;
        RECT 545.245 1684.105 545.415 1684.955 ;
        RECT 593.085 1684.105 593.715 1684.275 ;
        RECT 641.845 1684.105 642.015 1684.955 ;
        RECT 689.685 1684.105 690.315 1684.275 ;
        RECT 738.445 1684.105 738.615 1684.955 ;
        RECT 786.285 1684.105 786.915 1684.275 ;
        RECT 835.045 1684.105 835.215 1684.955 ;
        RECT 882.885 1684.105 883.515 1684.275 ;
        RECT 931.645 1684.105 931.815 1684.955 ;
        RECT 979.485 1684.105 980.115 1684.275 ;
        RECT 1028.245 1684.105 1028.415 1684.955 ;
        RECT 1159.345 1684.785 1159.515 1685.635 ;
        RECT 1231.565 1684.445 1231.735 1685.635 ;
        RECT 1249.505 1684.615 1249.675 1685.295 ;
        RECT 1249.045 1684.445 1249.675 1684.615 ;
        RECT 1296.885 1684.445 1297.055 1685.295 ;
        RECT 1594.965 1684.445 1595.135 1685.635 ;
        RECT 1606.925 1684.445 1607.095 1685.975 ;
        RECT 1690.185 1684.785 1690.355 1686.315 ;
        RECT 1690.645 1685.125 1690.815 1686.655 ;
        RECT 1076.085 1684.105 1076.715 1684.275 ;
        RECT 1883.845 1684.105 1884.015 1685.295 ;
        RECT 1937.665 1684.105 1937.835 1685.635 ;
      LAYER mcon ;
        RECT 1690.645 1686.485 1690.815 1686.655 ;
        RECT 1690.185 1686.145 1690.355 1686.315 ;
        RECT 1606.925 1685.805 1607.095 1685.975 ;
        RECT 96.285 1685.465 96.455 1685.635 ;
        RECT 111.005 1685.465 111.175 1685.635 ;
        RECT 1159.345 1685.465 1159.515 1685.635 ;
        RECT 48.445 1685.125 48.615 1685.295 ;
        RECT 158.845 1684.785 159.015 1684.955 ;
        RECT 255.445 1684.785 255.615 1684.955 ;
        RECT 241.185 1684.445 241.355 1684.615 ;
        RECT 193.345 1684.105 193.515 1684.275 ;
        RECT 352.045 1684.785 352.215 1684.955 ;
        RECT 337.785 1684.445 337.955 1684.615 ;
        RECT 289.945 1684.105 290.115 1684.275 ;
        RECT 448.645 1684.785 448.815 1684.955 ;
        RECT 434.385 1684.445 434.555 1684.615 ;
        RECT 386.545 1684.105 386.715 1684.275 ;
        RECT 545.245 1684.785 545.415 1684.955 ;
        RECT 530.985 1684.445 531.155 1684.615 ;
        RECT 483.145 1684.105 483.315 1684.275 ;
        RECT 641.845 1684.785 642.015 1684.955 ;
        RECT 738.445 1684.785 738.615 1684.955 ;
        RECT 835.045 1684.785 835.215 1684.955 ;
        RECT 931.645 1684.785 931.815 1684.955 ;
        RECT 1028.245 1684.785 1028.415 1684.955 ;
        RECT 1231.565 1685.465 1231.735 1685.635 ;
        RECT 1594.965 1685.465 1595.135 1685.635 ;
        RECT 1249.505 1685.125 1249.675 1685.295 ;
        RECT 1296.885 1685.125 1297.055 1685.295 ;
        RECT 1937.665 1685.465 1937.835 1685.635 ;
        RECT 1883.845 1685.125 1884.015 1685.295 ;
        RECT 593.545 1684.105 593.715 1684.275 ;
        RECT 690.145 1684.105 690.315 1684.275 ;
        RECT 786.745 1684.105 786.915 1684.275 ;
        RECT 883.345 1684.105 883.515 1684.275 ;
        RECT 979.945 1684.105 980.115 1684.275 ;
        RECT 1076.545 1684.105 1076.715 1684.275 ;
      LAYER met1 ;
        RECT 1793.150 1686.980 1793.470 1687.040 ;
        RECT 1706.300 1686.840 1793.470 1686.980 ;
        RECT 1690.585 1686.640 1690.875 1686.685 ;
        RECT 1706.300 1686.640 1706.440 1686.840 ;
        RECT 1793.150 1686.780 1793.470 1686.840 ;
        RECT 1690.585 1686.500 1706.440 1686.640 ;
        RECT 1690.585 1686.455 1690.875 1686.500 ;
        RECT 1690.125 1686.300 1690.415 1686.345 ;
        RECT 1666.280 1686.160 1690.415 1686.300 ;
        RECT 1606.865 1685.960 1607.155 1686.005 ;
        RECT 1666.280 1685.960 1666.420 1686.160 ;
        RECT 1690.125 1686.115 1690.415 1686.160 ;
        RECT 1558.640 1685.820 1569.820 1685.960 ;
        RECT 96.225 1685.620 96.515 1685.665 ;
        RECT 110.485 1685.620 110.775 1685.665 ;
        RECT 96.225 1685.480 110.775 1685.620 ;
        RECT 96.225 1685.435 96.515 1685.480 ;
        RECT 110.485 1685.435 110.775 1685.480 ;
        RECT 110.945 1685.620 111.235 1685.665 ;
        RECT 1159.285 1685.620 1159.575 1685.665 ;
        RECT 1231.505 1685.620 1231.795 1685.665 ;
        RECT 110.945 1685.480 144.740 1685.620 ;
        RECT 110.945 1685.435 111.235 1685.480 ;
        RECT 18.470 1685.280 18.790 1685.340 ;
        RECT 48.385 1685.280 48.675 1685.325 ;
        RECT 18.470 1685.140 48.675 1685.280 ;
        RECT 144.600 1685.280 144.740 1685.480 ;
        RECT 1159.285 1685.480 1231.795 1685.620 ;
        RECT 1159.285 1685.435 1159.575 1685.480 ;
        RECT 1231.505 1685.435 1231.795 1685.480 ;
        RECT 1249.445 1685.280 1249.735 1685.325 ;
        RECT 1296.825 1685.280 1297.115 1685.325 ;
        RECT 1558.640 1685.280 1558.780 1685.820 ;
        RECT 1569.680 1685.620 1569.820 1685.820 ;
        RECT 1606.865 1685.820 1666.420 1685.960 ;
        RECT 1606.865 1685.775 1607.155 1685.820 ;
        RECT 1594.905 1685.620 1595.195 1685.665 ;
        RECT 1937.605 1685.620 1937.895 1685.665 ;
        RECT 1569.680 1685.480 1595.195 1685.620 ;
        RECT 1594.905 1685.435 1595.195 1685.480 ;
        RECT 1920.200 1685.480 1937.895 1685.620 ;
        RECT 1690.585 1685.280 1690.875 1685.325 ;
        RECT 144.600 1685.140 158.540 1685.280 ;
        RECT 18.470 1685.080 18.790 1685.140 ;
        RECT 48.385 1685.095 48.675 1685.140 ;
        RECT 158.400 1684.940 158.540 1685.140 ;
        RECT 1249.445 1685.140 1297.115 1685.280 ;
        RECT 1249.445 1685.095 1249.735 1685.140 ;
        RECT 1296.825 1685.095 1297.115 1685.140 ;
        RECT 1514.020 1685.140 1558.780 1685.280 ;
        RECT 1690.200 1685.140 1690.875 1685.280 ;
        RECT 158.785 1684.940 159.075 1684.985 ;
        RECT 255.385 1684.940 255.675 1684.985 ;
        RECT 351.985 1684.940 352.275 1684.985 ;
        RECT 448.585 1684.940 448.875 1684.985 ;
        RECT 545.185 1684.940 545.475 1684.985 ;
        RECT 641.785 1684.940 642.075 1684.985 ;
        RECT 738.385 1684.940 738.675 1684.985 ;
        RECT 834.985 1684.940 835.275 1684.985 ;
        RECT 931.585 1684.940 931.875 1684.985 ;
        RECT 1028.185 1684.940 1028.475 1684.985 ;
        RECT 1159.285 1684.940 1159.575 1684.985 ;
        RECT 1514.020 1684.940 1514.160 1685.140 ;
        RECT 1690.200 1684.985 1690.340 1685.140 ;
        RECT 1690.585 1685.095 1690.875 1685.140 ;
        RECT 1801.890 1685.280 1802.210 1685.340 ;
        RECT 1883.785 1685.280 1884.075 1685.325 ;
        RECT 1920.200 1685.280 1920.340 1685.480 ;
        RECT 1937.605 1685.435 1937.895 1685.480 ;
        RECT 1801.890 1685.140 1884.075 1685.280 ;
        RECT 1801.890 1685.080 1802.210 1685.140 ;
        RECT 1883.785 1685.095 1884.075 1685.140 ;
        RECT 1897.660 1685.140 1920.340 1685.280 ;
        RECT 158.400 1684.800 159.075 1684.940 ;
        RECT 158.785 1684.755 159.075 1684.800 ;
        RECT 255.000 1684.800 255.675 1684.940 ;
        RECT 48.385 1684.600 48.675 1684.645 ;
        RECT 96.225 1684.600 96.515 1684.645 ;
        RECT 48.385 1684.460 96.515 1684.600 ;
        RECT 48.385 1684.415 48.675 1684.460 ;
        RECT 96.225 1684.415 96.515 1684.460 ;
        RECT 241.125 1684.600 241.415 1684.645 ;
        RECT 255.000 1684.600 255.140 1684.800 ;
        RECT 255.385 1684.755 255.675 1684.800 ;
        RECT 351.600 1684.800 352.275 1684.940 ;
        RECT 241.125 1684.460 255.140 1684.600 ;
        RECT 337.725 1684.600 338.015 1684.645 ;
        RECT 351.600 1684.600 351.740 1684.800 ;
        RECT 351.985 1684.755 352.275 1684.800 ;
        RECT 448.200 1684.800 448.875 1684.940 ;
        RECT 337.725 1684.460 351.740 1684.600 ;
        RECT 434.325 1684.600 434.615 1684.645 ;
        RECT 448.200 1684.600 448.340 1684.800 ;
        RECT 448.585 1684.755 448.875 1684.800 ;
        RECT 544.800 1684.800 545.475 1684.940 ;
        RECT 434.325 1684.460 448.340 1684.600 ;
        RECT 530.925 1684.600 531.215 1684.645 ;
        RECT 544.800 1684.600 544.940 1684.800 ;
        RECT 545.185 1684.755 545.475 1684.800 ;
        RECT 641.400 1684.800 642.075 1684.940 ;
        RECT 641.400 1684.600 641.540 1684.800 ;
        RECT 641.785 1684.755 642.075 1684.800 ;
        RECT 738.000 1684.800 738.675 1684.940 ;
        RECT 738.000 1684.600 738.140 1684.800 ;
        RECT 738.385 1684.755 738.675 1684.800 ;
        RECT 834.600 1684.800 835.275 1684.940 ;
        RECT 834.600 1684.600 834.740 1684.800 ;
        RECT 834.985 1684.755 835.275 1684.800 ;
        RECT 931.200 1684.800 931.875 1684.940 ;
        RECT 931.200 1684.600 931.340 1684.800 ;
        RECT 931.585 1684.755 931.875 1684.800 ;
        RECT 1027.800 1684.800 1028.475 1684.940 ;
        RECT 1027.800 1684.600 1027.940 1684.800 ;
        RECT 1028.185 1684.755 1028.475 1684.800 ;
        RECT 1124.400 1684.800 1159.575 1684.940 ;
        RECT 1124.400 1684.600 1124.540 1684.800 ;
        RECT 1159.285 1684.755 1159.575 1684.800 ;
        RECT 1304.260 1684.800 1514.160 1684.940 ;
        RECT 530.925 1684.460 544.940 1684.600 ;
        RECT 599.540 1684.460 641.540 1684.600 ;
        RECT 696.140 1684.460 738.140 1684.600 ;
        RECT 792.740 1684.460 834.740 1684.600 ;
        RECT 889.340 1684.460 931.340 1684.600 ;
        RECT 985.940 1684.460 1027.940 1684.600 ;
        RECT 1082.540 1684.460 1124.540 1684.600 ;
        RECT 1231.505 1684.600 1231.795 1684.645 ;
        RECT 1248.985 1684.600 1249.275 1684.645 ;
        RECT 1231.505 1684.460 1249.275 1684.600 ;
        RECT 241.125 1684.415 241.415 1684.460 ;
        RECT 337.725 1684.415 338.015 1684.460 ;
        RECT 434.325 1684.415 434.615 1684.460 ;
        RECT 530.925 1684.415 531.215 1684.460 ;
        RECT 158.785 1684.260 159.075 1684.305 ;
        RECT 193.285 1684.260 193.575 1684.305 ;
        RECT 158.785 1684.120 193.575 1684.260 ;
        RECT 158.785 1684.075 159.075 1684.120 ;
        RECT 193.285 1684.075 193.575 1684.120 ;
        RECT 255.385 1684.260 255.675 1684.305 ;
        RECT 289.885 1684.260 290.175 1684.305 ;
        RECT 255.385 1684.120 290.175 1684.260 ;
        RECT 255.385 1684.075 255.675 1684.120 ;
        RECT 289.885 1684.075 290.175 1684.120 ;
        RECT 351.985 1684.260 352.275 1684.305 ;
        RECT 386.485 1684.260 386.775 1684.305 ;
        RECT 351.985 1684.120 386.775 1684.260 ;
        RECT 351.985 1684.075 352.275 1684.120 ;
        RECT 386.485 1684.075 386.775 1684.120 ;
        RECT 448.585 1684.260 448.875 1684.305 ;
        RECT 483.085 1684.260 483.375 1684.305 ;
        RECT 448.585 1684.120 483.375 1684.260 ;
        RECT 448.585 1684.075 448.875 1684.120 ;
        RECT 483.085 1684.075 483.375 1684.120 ;
        RECT 545.185 1684.260 545.475 1684.305 ;
        RECT 593.025 1684.260 593.315 1684.305 ;
        RECT 545.185 1684.120 593.315 1684.260 ;
        RECT 545.185 1684.075 545.475 1684.120 ;
        RECT 593.025 1684.075 593.315 1684.120 ;
        RECT 593.485 1684.260 593.775 1684.305 ;
        RECT 599.540 1684.260 599.680 1684.460 ;
        RECT 593.485 1684.120 599.680 1684.260 ;
        RECT 641.785 1684.260 642.075 1684.305 ;
        RECT 689.625 1684.260 689.915 1684.305 ;
        RECT 641.785 1684.120 689.915 1684.260 ;
        RECT 593.485 1684.075 593.775 1684.120 ;
        RECT 641.785 1684.075 642.075 1684.120 ;
        RECT 689.625 1684.075 689.915 1684.120 ;
        RECT 690.085 1684.260 690.375 1684.305 ;
        RECT 696.140 1684.260 696.280 1684.460 ;
        RECT 690.085 1684.120 696.280 1684.260 ;
        RECT 738.385 1684.260 738.675 1684.305 ;
        RECT 786.225 1684.260 786.515 1684.305 ;
        RECT 738.385 1684.120 786.515 1684.260 ;
        RECT 690.085 1684.075 690.375 1684.120 ;
        RECT 738.385 1684.075 738.675 1684.120 ;
        RECT 786.225 1684.075 786.515 1684.120 ;
        RECT 786.685 1684.260 786.975 1684.305 ;
        RECT 792.740 1684.260 792.880 1684.460 ;
        RECT 786.685 1684.120 792.880 1684.260 ;
        RECT 834.985 1684.260 835.275 1684.305 ;
        RECT 882.825 1684.260 883.115 1684.305 ;
        RECT 834.985 1684.120 883.115 1684.260 ;
        RECT 786.685 1684.075 786.975 1684.120 ;
        RECT 834.985 1684.075 835.275 1684.120 ;
        RECT 882.825 1684.075 883.115 1684.120 ;
        RECT 883.285 1684.260 883.575 1684.305 ;
        RECT 889.340 1684.260 889.480 1684.460 ;
        RECT 883.285 1684.120 889.480 1684.260 ;
        RECT 931.585 1684.260 931.875 1684.305 ;
        RECT 979.425 1684.260 979.715 1684.305 ;
        RECT 931.585 1684.120 979.715 1684.260 ;
        RECT 883.285 1684.075 883.575 1684.120 ;
        RECT 931.585 1684.075 931.875 1684.120 ;
        RECT 979.425 1684.075 979.715 1684.120 ;
        RECT 979.885 1684.260 980.175 1684.305 ;
        RECT 985.940 1684.260 986.080 1684.460 ;
        RECT 979.885 1684.120 986.080 1684.260 ;
        RECT 1028.185 1684.260 1028.475 1684.305 ;
        RECT 1076.025 1684.260 1076.315 1684.305 ;
        RECT 1028.185 1684.120 1076.315 1684.260 ;
        RECT 979.885 1684.075 980.175 1684.120 ;
        RECT 1028.185 1684.075 1028.475 1684.120 ;
        RECT 1076.025 1684.075 1076.315 1684.120 ;
        RECT 1076.485 1684.260 1076.775 1684.305 ;
        RECT 1082.540 1684.260 1082.680 1684.460 ;
        RECT 1231.505 1684.415 1231.795 1684.460 ;
        RECT 1248.985 1684.415 1249.275 1684.460 ;
        RECT 1296.825 1684.600 1297.115 1684.645 ;
        RECT 1304.260 1684.600 1304.400 1684.800 ;
        RECT 1690.125 1684.755 1690.415 1684.985 ;
        RECT 1897.660 1684.940 1897.800 1685.140 ;
        RECT 1890.760 1684.800 1897.800 1684.940 ;
        RECT 1296.825 1684.460 1304.400 1684.600 ;
        RECT 1594.905 1684.600 1595.195 1684.645 ;
        RECT 1606.865 1684.600 1607.155 1684.645 ;
        RECT 1594.905 1684.460 1607.155 1684.600 ;
        RECT 1296.825 1684.415 1297.115 1684.460 ;
        RECT 1594.905 1684.415 1595.195 1684.460 ;
        RECT 1606.865 1684.415 1607.155 1684.460 ;
        RECT 1076.485 1684.120 1082.680 1684.260 ;
        RECT 1883.785 1684.260 1884.075 1684.305 ;
        RECT 1890.760 1684.260 1890.900 1684.800 ;
        RECT 1883.785 1684.120 1890.900 1684.260 ;
        RECT 1937.605 1684.260 1937.895 1684.305 ;
        RECT 1948.630 1684.260 1948.950 1684.320 ;
        RECT 1937.605 1684.120 1948.950 1684.260 ;
        RECT 1076.485 1684.075 1076.775 1684.120 ;
        RECT 1883.785 1684.075 1884.075 1684.120 ;
        RECT 1937.605 1684.075 1937.895 1684.120 ;
        RECT 1948.630 1684.060 1948.950 1684.120 ;
        RECT 193.285 1683.580 193.575 1683.625 ;
        RECT 241.125 1683.580 241.415 1683.625 ;
        RECT 193.285 1683.440 241.415 1683.580 ;
        RECT 193.285 1683.395 193.575 1683.440 ;
        RECT 241.125 1683.395 241.415 1683.440 ;
        RECT 289.885 1683.580 290.175 1683.625 ;
        RECT 337.725 1683.580 338.015 1683.625 ;
        RECT 289.885 1683.440 338.015 1683.580 ;
        RECT 289.885 1683.395 290.175 1683.440 ;
        RECT 337.725 1683.395 338.015 1683.440 ;
        RECT 386.485 1683.580 386.775 1683.625 ;
        RECT 434.325 1683.580 434.615 1683.625 ;
        RECT 386.485 1683.440 434.615 1683.580 ;
        RECT 386.485 1683.395 386.775 1683.440 ;
        RECT 434.325 1683.395 434.615 1683.440 ;
        RECT 483.085 1683.580 483.375 1683.625 ;
        RECT 530.925 1683.580 531.215 1683.625 ;
        RECT 483.085 1683.440 531.215 1683.580 ;
        RECT 483.085 1683.395 483.375 1683.440 ;
        RECT 530.925 1683.395 531.215 1683.440 ;
      LAYER via ;
        RECT 1793.180 1686.780 1793.440 1687.040 ;
        RECT 18.500 1685.080 18.760 1685.340 ;
        RECT 1801.920 1685.080 1802.180 1685.340 ;
        RECT 1948.660 1684.060 1948.920 1684.320 ;
      LAYER met2 ;
        RECT 18.490 2046.275 18.770 2046.645 ;
        RECT 18.560 1685.370 18.700 2046.275 ;
        RECT 1948.650 1700.000 1948.930 1704.000 ;
        RECT 1793.180 1686.925 1793.440 1687.070 ;
        RECT 1793.170 1686.555 1793.450 1686.925 ;
        RECT 1801.910 1686.555 1802.190 1686.925 ;
        RECT 1801.980 1685.370 1802.120 1686.555 ;
        RECT 18.500 1685.050 18.760 1685.370 ;
        RECT 1801.920 1685.050 1802.180 1685.370 ;
        RECT 1948.720 1684.350 1948.860 1700.000 ;
        RECT 1948.660 1684.030 1948.920 1684.350 ;
      LAYER via2 ;
        RECT 18.490 2046.320 18.770 2046.600 ;
        RECT 1793.170 1686.600 1793.450 1686.880 ;
        RECT 1801.910 1686.600 1802.190 1686.880 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT -4.800 2045.860 0.300 2047.060 ;
=======
        RECT 1137.645 2379.130 1137.975 2379.145 ;
        RECT 1150.000 2379.130 1154.000 2379.280 ;
        RECT 1137.645 2378.830 1154.000 2379.130 ;
        RECT 1137.645 2378.815 1137.975 2378.830 ;
        RECT 1150.000 2378.680 1154.000 2378.830 ;
=======
>>>>>>> re-updated local openlane
        RECT -4.800 2046.610 2.400 2047.060 ;
        RECT 18.465 2046.610 18.795 2046.625 ;
        RECT -4.800 2046.310 18.795 2046.610 ;
        RECT -4.800 2045.860 2.400 2046.310 ;
<<<<<<< HEAD
        RECT 14.325 2046.295 14.655 2046.310 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 18.465 2046.295 18.795 2046.310 ;
        RECT 1793.145 1686.890 1793.475 1686.905 ;
        RECT 1801.885 1686.890 1802.215 1686.905 ;
        RECT 1793.145 1686.590 1802.215 1686.890 ;
        RECT 1793.145 1686.575 1793.475 1686.590 ;
        RECT 1801.885 1686.575 1802.215 1686.590 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1137.190 503.440 1137.510 503.500 ;
        RECT 2900.830 503.440 2901.150 503.500 ;
        RECT 1137.190 503.300 2901.150 503.440 ;
        RECT 1137.190 503.240 1137.510 503.300 ;
        RECT 2900.830 503.240 2901.150 503.300 ;
      LAYER via ;
        RECT 1137.220 503.240 1137.480 503.500 ;
        RECT 2900.860 503.240 2901.120 503.500 ;
      LAYER met2 ;
        RECT 1137.210 1921.835 1137.490 1922.205 ;
        RECT 1137.280 503.530 1137.420 1921.835 ;
        RECT 1137.220 503.210 1137.480 503.530 ;
        RECT 2900.860 503.210 2901.120 503.530 ;
        RECT 2900.920 498.965 2901.060 503.210 ;
        RECT 2900.850 498.595 2901.130 498.965 ;
      LAYER via2 ;
        RECT 1137.210 1921.880 1137.490 1922.160 ;
        RECT 2900.850 498.640 2901.130 498.920 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 498.180 2924.800 499.380 ;
=======
        RECT 1946.000 1767.130 1950.000 1767.280 ;
        RECT 1962.885 1767.130 1963.215 1767.145 ;
        RECT 1946.000 1766.830 1963.215 1767.130 ;
        RECT 1946.000 1766.680 1950.000 1766.830 ;
        RECT 1962.885 1766.815 1963.215 1766.830 ;
=======
        RECT 1137.185 1922.170 1137.515 1922.185 ;
        RECT 1150.000 1922.170 1154.000 1922.320 ;
        RECT 1137.185 1921.870 1154.000 1922.170 ;
        RECT 1137.185 1921.855 1137.515 1921.870 ;
        RECT 1150.000 1921.720 1154.000 1921.870 ;
>>>>>>> re-updated local openlane
        RECT 2900.825 498.930 2901.155 498.945 ;
        RECT 2917.600 498.930 2924.800 499.380 ;
        RECT 2900.825 498.630 2924.800 498.930 ;
        RECT 2900.825 498.615 2901.155 498.630 ;
        RECT 2917.600 498.180 2924.800 498.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 99.890 2505.020 100.210 2505.080 ;
        RECT 1946.330 2505.020 1946.650 2505.080 ;
        RECT 99.890 2504.880 1946.650 2505.020 ;
        RECT 99.890 2504.820 100.210 2504.880 ;
        RECT 1946.330 2504.820 1946.650 2504.880 ;
        RECT 15.250 1766.200 15.570 1766.260 ;
        RECT 99.890 1766.200 100.210 1766.260 ;
        RECT 15.250 1766.060 100.210 1766.200 ;
        RECT 15.250 1766.000 15.570 1766.060 ;
        RECT 99.890 1766.000 100.210 1766.060 ;
      LAYER via ;
        RECT 99.920 2504.820 100.180 2505.080 ;
        RECT 1946.360 2504.820 1946.620 2505.080 ;
        RECT 15.280 1766.000 15.540 1766.260 ;
        RECT 99.920 1766.000 100.180 1766.260 ;
      LAYER met2 ;
        RECT 99.920 2504.790 100.180 2505.110 ;
        RECT 1946.360 2504.790 1946.620 2505.110 ;
        RECT 99.980 1766.290 100.120 2504.790 ;
        RECT 1946.420 2500.000 1946.560 2504.790 ;
        RECT 1946.350 2496.000 1946.630 2500.000 ;
        RECT 15.280 1765.970 15.540 1766.290 ;
        RECT 99.920 1765.970 100.180 1766.290 ;
        RECT 15.340 1759.685 15.480 1765.970 ;
        RECT 15.270 1759.315 15.550 1759.685 ;
      LAYER via2 ;
        RECT 15.270 1759.360 15.550 1759.640 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT -4.800 1758.900 0.300 1760.100 ;
=======
        RECT 1131.665 2459.370 1131.995 2459.385 ;
        RECT 1150.000 2459.370 1154.000 2459.520 ;
        RECT 1131.665 2459.070 1154.000 2459.370 ;
        RECT 1131.665 2459.055 1131.995 2459.070 ;
        RECT 1150.000 2458.920 1154.000 2459.070 ;
=======
>>>>>>> re-updated local openlane
        RECT -4.800 1759.650 2.400 1760.100 ;
        RECT 15.245 1759.650 15.575 1759.665 ;
        RECT -4.800 1759.350 15.575 1759.650 ;
        RECT -4.800 1758.900 2.400 1759.350 ;
<<<<<<< HEAD
        RECT 15.705 1759.335 16.035 1759.350 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 15.245 1759.335 15.575 1759.350 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1136.730 738.040 1137.050 738.100 ;
        RECT 2900.830 738.040 2901.150 738.100 ;
        RECT 1136.730 737.900 2901.150 738.040 ;
        RECT 1136.730 737.840 1137.050 737.900 ;
        RECT 2900.830 737.840 2901.150 737.900 ;
      LAYER via ;
        RECT 1136.760 737.840 1137.020 738.100 ;
        RECT 2900.860 737.840 2901.120 738.100 ;
      LAYER met2 ;
        RECT 1136.750 2010.915 1137.030 2011.285 ;
        RECT 1136.820 738.130 1136.960 2010.915 ;
        RECT 1136.760 737.810 1137.020 738.130 ;
        RECT 2900.860 737.810 2901.120 738.130 ;
        RECT 2900.920 733.565 2901.060 737.810 ;
        RECT 2900.850 733.195 2901.130 733.565 ;
      LAYER via2 ;
        RECT 1136.750 2010.960 1137.030 2011.240 ;
        RECT 2900.850 733.240 2901.130 733.520 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 732.780 2924.800 733.980 ;
=======
=======
        RECT 1136.725 2011.250 1137.055 2011.265 ;
        RECT 1150.000 2011.250 1154.000 2011.400 ;
        RECT 1136.725 2010.950 1154.000 2011.250 ;
        RECT 1136.725 2010.935 1137.055 2010.950 ;
        RECT 1150.000 2010.800 1154.000 2010.950 ;
>>>>>>> re-updated local openlane
        RECT 2900.825 733.530 2901.155 733.545 ;
        RECT 2917.600 733.530 2924.800 733.980 ;
        RECT 2900.825 733.230 2924.800 733.530 ;
        RECT 2900.825 733.215 2901.155 733.230 ;
        RECT 2917.600 732.780 2924.800 733.230 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1962.890 972.640 1963.210 972.700 ;
        RECT 2900.830 972.640 2901.150 972.700 ;
        RECT 1962.890 972.500 2901.150 972.640 ;
        RECT 1962.890 972.440 1963.210 972.500 ;
        RECT 2900.830 972.440 2901.150 972.500 ;
      LAYER via ;
        RECT 1962.920 972.440 1963.180 972.700 ;
        RECT 2900.860 972.440 2901.120 972.700 ;
      LAYER met2 ;
        RECT 1962.910 1766.795 1963.190 1767.165 ;
        RECT 1962.980 972.730 1963.120 1766.795 ;
        RECT 1962.920 972.410 1963.180 972.730 ;
        RECT 2900.860 972.410 2901.120 972.730 ;
        RECT 2900.920 968.165 2901.060 972.410 ;
        RECT 2900.850 967.795 2901.130 968.165 ;
      LAYER via2 ;
        RECT 1962.910 1766.840 1963.190 1767.120 ;
        RECT 2900.850 967.840 2901.130 968.120 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 967.380 2924.800 968.580 ;
=======
        RECT 1137.645 1819.490 1137.975 1819.505 ;
        RECT 1150.000 1819.490 1154.000 1819.640 ;
        RECT 1137.645 1819.190 1154.000 1819.490 ;
        RECT 1137.645 1819.175 1137.975 1819.190 ;
        RECT 1150.000 1819.040 1154.000 1819.190 ;
=======
        RECT 1946.000 1767.130 1950.000 1767.280 ;
        RECT 1962.885 1767.130 1963.215 1767.145 ;
        RECT 1946.000 1766.830 1963.215 1767.130 ;
        RECT 1946.000 1766.680 1950.000 1766.830 ;
        RECT 1962.885 1766.815 1963.215 1766.830 ;
>>>>>>> re-updated local openlane
        RECT 2900.825 968.130 2901.155 968.145 ;
        RECT 2917.600 968.130 2924.800 968.580 ;
        RECT 2900.825 967.830 2924.800 968.130 ;
        RECT 2900.825 967.815 2901.155 967.830 ;
        RECT 2917.600 967.380 2924.800 967.830 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1963.350 1207.240 1963.670 1207.300 ;
        RECT 2900.830 1207.240 2901.150 1207.300 ;
        RECT 1963.350 1207.100 2901.150 1207.240 ;
        RECT 1963.350 1207.040 1963.670 1207.100 ;
        RECT 2900.830 1207.040 2901.150 1207.100 ;
      LAYER via ;
        RECT 1963.380 1207.040 1963.640 1207.300 ;
        RECT 2900.860 1207.040 2901.120 1207.300 ;
      LAYER met2 ;
        RECT 1963.370 1900.075 1963.650 1900.445 ;
        RECT 1963.440 1207.330 1963.580 1900.075 ;
        RECT 1963.380 1207.010 1963.640 1207.330 ;
        RECT 2900.860 1207.010 2901.120 1207.330 ;
        RECT 2900.920 1202.765 2901.060 1207.010 ;
        RECT 2900.850 1202.395 2901.130 1202.765 ;
      LAYER via2 ;
        RECT 1963.370 1900.120 1963.650 1900.400 ;
        RECT 2900.850 1202.440 2901.130 1202.720 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1201.980 2924.800 1203.180 ;
=======
=======
        RECT 1946.000 1900.410 1950.000 1900.560 ;
        RECT 1963.345 1900.410 1963.675 1900.425 ;
        RECT 1946.000 1900.110 1963.675 1900.410 ;
        RECT 1946.000 1899.960 1950.000 1900.110 ;
        RECT 1963.345 1900.095 1963.675 1900.110 ;
>>>>>>> re-updated local openlane
        RECT 2900.825 1202.730 2901.155 1202.745 ;
        RECT 2917.600 1202.730 2924.800 1203.180 ;
        RECT 2900.825 1202.430 2924.800 1202.730 ;
        RECT 2900.825 1202.415 2901.155 1202.430 ;
        RECT 2917.600 1201.980 2924.800 1202.430 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1888.370 2512.160 1888.690 2512.220 ;
        RECT 1977.150 2512.160 1977.470 2512.220 ;
        RECT 1888.370 2512.020 1977.470 2512.160 ;
        RECT 1888.370 2511.960 1888.690 2512.020 ;
        RECT 1977.150 2511.960 1977.470 2512.020 ;
        RECT 1977.150 1441.840 1977.470 1441.900 ;
        RECT 2900.830 1441.840 2901.150 1441.900 ;
        RECT 1977.150 1441.700 2901.150 1441.840 ;
        RECT 1977.150 1441.640 1977.470 1441.700 ;
        RECT 2900.830 1441.640 2901.150 1441.700 ;
      LAYER via ;
        RECT 1888.400 2511.960 1888.660 2512.220 ;
        RECT 1977.180 2511.960 1977.440 2512.220 ;
        RECT 1977.180 1441.640 1977.440 1441.900 ;
        RECT 2900.860 1441.640 2901.120 1441.900 ;
      LAYER met2 ;
        RECT 1888.400 2511.930 1888.660 2512.250 ;
        RECT 1977.180 2511.930 1977.440 2512.250 ;
        RECT 1888.460 2500.000 1888.600 2511.930 ;
        RECT 1888.390 2496.000 1888.670 2500.000 ;
        RECT 1977.240 1441.930 1977.380 2511.930 ;
        RECT 1977.180 1441.610 1977.440 1441.930 ;
        RECT 2900.860 1441.610 2901.120 1441.930 ;
        RECT 2900.920 1437.365 2901.060 1441.610 ;
        RECT 2900.850 1436.995 2901.130 1437.365 ;
      LAYER via2 ;
        RECT 2900.850 1437.040 2901.130 1437.320 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1436.580 2924.800 1437.780 ;
=======
        RECT 1137.185 1899.730 1137.515 1899.745 ;
        RECT 1150.000 1899.730 1154.000 1899.880 ;
        RECT 1137.185 1899.430 1154.000 1899.730 ;
        RECT 1137.185 1899.415 1137.515 1899.430 ;
        RECT 1150.000 1899.280 1154.000 1899.430 ;
=======
>>>>>>> re-updated local openlane
        RECT 2900.825 1437.330 2901.155 1437.345 ;
        RECT 2917.600 1437.330 2924.800 1437.780 ;
        RECT 2900.825 1437.030 2924.800 1437.330 ;
        RECT 2900.825 1437.015 2901.155 1437.030 ;
        RECT 2917.600 1436.580 2924.800 1437.030 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1894.810 2511.820 1895.130 2511.880 ;
        RECT 1990.950 2511.820 1991.270 2511.880 ;
        RECT 1894.810 2511.680 1991.270 2511.820 ;
        RECT 1894.810 2511.620 1895.130 2511.680 ;
        RECT 1990.950 2511.620 1991.270 2511.680 ;
        RECT 1990.950 1676.440 1991.270 1676.500 ;
        RECT 2900.830 1676.440 2901.150 1676.500 ;
        RECT 1990.950 1676.300 2901.150 1676.440 ;
        RECT 1990.950 1676.240 1991.270 1676.300 ;
        RECT 2900.830 1676.240 2901.150 1676.300 ;
      LAYER via ;
        RECT 1894.840 2511.620 1895.100 2511.880 ;
        RECT 1990.980 2511.620 1991.240 2511.880 ;
        RECT 1990.980 1676.240 1991.240 1676.500 ;
        RECT 2900.860 1676.240 2901.120 1676.500 ;
      LAYER met2 ;
        RECT 1894.840 2511.590 1895.100 2511.910 ;
        RECT 1990.980 2511.590 1991.240 2511.910 ;
        RECT 1894.900 2500.000 1895.040 2511.590 ;
        RECT 1894.830 2496.000 1895.110 2500.000 ;
        RECT 1991.040 1676.530 1991.180 2511.590 ;
        RECT 1990.980 1676.210 1991.240 1676.530 ;
        RECT 2900.860 1676.210 2901.120 1676.530 ;
        RECT 2900.920 1671.965 2901.060 1676.210 ;
        RECT 2900.850 1671.595 2901.130 1671.965 ;
      LAYER via2 ;
        RECT 2900.850 1671.640 2901.130 1671.920 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1671.180 2924.800 1672.380 ;
=======
        RECT 2900.825 1671.930 2901.155 1671.945 ;
        RECT 2917.600 1671.930 2924.800 1672.380 ;
        RECT 2900.825 1671.630 2924.800 1671.930 ;
        RECT 2900.825 1671.615 2901.155 1671.630 ;
        RECT 2917.600 1671.180 2924.800 1671.630 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1905.780 2924.800 1906.980 ;
=======
        RECT 1136.470 1979.290 1136.850 1979.300 ;
        RECT 1150.000 1979.290 1154.000 1979.440 ;
        RECT 1136.470 1978.990 1154.000 1979.290 ;
        RECT 1136.470 1978.980 1136.850 1978.990 ;
        RECT 1150.000 1978.840 1154.000 1978.990 ;
=======
        RECT 1136.470 2099.650 1136.850 2099.660 ;
        RECT 1150.000 2099.650 1154.000 2099.800 ;
        RECT 1136.470 2099.350 1154.000 2099.650 ;
        RECT 1136.470 2099.340 1136.850 2099.350 ;
        RECT 1150.000 2099.200 1154.000 2099.350 ;
>>>>>>> re-updated local openlane
        RECT 2898.270 1906.530 2898.650 1906.540 ;
        RECT 2917.600 1906.530 2924.800 1906.980 ;
        RECT 2898.270 1906.230 2924.800 1906.530 ;
        RECT 2898.270 1906.220 2898.650 1906.230 ;
        RECT 2917.600 1905.780 2924.800 1906.230 ;
      LAYER via3 ;
        RECT 1136.500 2099.340 1136.820 2099.660 ;
        RECT 2898.300 1906.220 2898.620 1906.540 ;
      LAYER met4 ;
        RECT 1136.495 2099.335 1136.825 2099.665 ;
        RECT 1136.510 1906.290 1136.810 2099.335 ;
        RECT 2897.870 1908.510 2899.050 1909.690 ;
        RECT 2898.310 1906.545 2898.610 1908.510 ;
        RECT 1136.070 1905.110 1137.250 1906.290 ;
        RECT 2898.295 1906.215 2898.625 1906.545 ;
      LAYER met5 ;
        RECT 1170.820 1911.700 1222.100 1913.300 ;
        RECT 1170.820 1906.500 1172.420 1911.700 ;
        RECT 1135.860 1904.900 1172.420 1906.500 ;
        RECT 1220.500 1906.500 1222.100 1911.700 ;
        RECT 1267.420 1911.700 1318.700 1913.300 ;
        RECT 1267.420 1906.500 1269.020 1911.700 ;
        RECT 1220.500 1904.900 1269.020 1906.500 ;
        RECT 1317.100 1906.500 1318.700 1911.700 ;
        RECT 1364.020 1911.700 1415.300 1913.300 ;
        RECT 1364.020 1906.500 1365.620 1911.700 ;
        RECT 1317.100 1904.900 1365.620 1906.500 ;
        RECT 1413.700 1906.500 1415.300 1911.700 ;
        RECT 1460.620 1911.700 1511.900 1913.300 ;
        RECT 1460.620 1906.500 1462.220 1911.700 ;
        RECT 1413.700 1904.900 1462.220 1906.500 ;
        RECT 1510.300 1906.500 1511.900 1911.700 ;
        RECT 1557.220 1911.700 1608.500 1913.300 ;
        RECT 1557.220 1906.500 1558.820 1911.700 ;
        RECT 1510.300 1904.900 1558.820 1906.500 ;
        RECT 1606.900 1906.500 1608.500 1911.700 ;
        RECT 1653.820 1911.700 1705.100 1913.300 ;
        RECT 1653.820 1906.500 1655.420 1911.700 ;
        RECT 1606.900 1904.900 1655.420 1906.500 ;
        RECT 1703.500 1906.500 1705.100 1911.700 ;
        RECT 1750.420 1911.700 1801.700 1913.300 ;
        RECT 1750.420 1906.500 1752.020 1911.700 ;
        RECT 1703.500 1904.900 1752.020 1906.500 ;
        RECT 1800.100 1906.500 1801.700 1911.700 ;
        RECT 1847.020 1911.700 1898.300 1913.300 ;
        RECT 1847.020 1906.500 1848.620 1911.700 ;
        RECT 1800.100 1904.900 1848.620 1906.500 ;
        RECT 1896.700 1906.500 1898.300 1911.700 ;
        RECT 1943.620 1911.700 1994.900 1913.300 ;
        RECT 1943.620 1906.500 1945.220 1911.700 ;
        RECT 1896.700 1904.900 1945.220 1906.500 ;
        RECT 1993.300 1906.500 1994.900 1911.700 ;
        RECT 2040.220 1911.700 2091.500 1913.300 ;
        RECT 2040.220 1906.500 2041.820 1911.700 ;
        RECT 1993.300 1904.900 2041.820 1906.500 ;
        RECT 2089.900 1906.500 2091.500 1911.700 ;
        RECT 2136.820 1911.700 2188.100 1913.300 ;
        RECT 2136.820 1906.500 2138.420 1911.700 ;
        RECT 2089.900 1904.900 2138.420 1906.500 ;
        RECT 2186.500 1906.500 2188.100 1911.700 ;
        RECT 2233.420 1911.700 2284.700 1913.300 ;
        RECT 2233.420 1906.500 2235.020 1911.700 ;
        RECT 2186.500 1904.900 2235.020 1906.500 ;
        RECT 2283.100 1906.500 2284.700 1911.700 ;
        RECT 2330.020 1911.700 2381.300 1913.300 ;
        RECT 2330.020 1906.500 2331.620 1911.700 ;
        RECT 2283.100 1904.900 2331.620 1906.500 ;
        RECT 2379.700 1906.500 2381.300 1911.700 ;
        RECT 2426.620 1911.700 2477.900 1913.300 ;
        RECT 2426.620 1906.500 2428.220 1911.700 ;
        RECT 2379.700 1904.900 2428.220 1906.500 ;
        RECT 2476.300 1906.500 2477.900 1911.700 ;
        RECT 2523.220 1911.700 2574.500 1913.300 ;
        RECT 2523.220 1906.500 2524.820 1911.700 ;
        RECT 2476.300 1904.900 2524.820 1906.500 ;
        RECT 2572.900 1906.500 2574.500 1911.700 ;
        RECT 2620.740 1911.700 2740.100 1913.300 ;
        RECT 2620.740 1906.500 2622.340 1911.700 ;
        RECT 2572.900 1904.900 2622.340 1906.500 ;
        RECT 2738.500 1906.500 2740.100 1911.700 ;
        RECT 2766.100 1911.700 2837.620 1913.300 ;
        RECT 2766.100 1906.500 2767.700 1911.700 ;
        RECT 2738.500 1904.900 2767.700 1906.500 ;
        RECT 2836.020 1906.500 2837.620 1911.700 ;
        RECT 2882.940 1911.700 2899.260 1913.300 ;
        RECT 2882.940 1906.500 2884.540 1911.700 ;
        RECT 2897.660 1908.300 2899.260 1911.700 ;
        RECT 2836.020 1904.900 2884.540 1906.500 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1944.950 2139.180 1945.270 2139.240 ;
        RECT 2899.450 2139.180 2899.770 2139.240 ;
        RECT 1944.950 2139.040 2899.770 2139.180 ;
        RECT 1944.950 2138.980 1945.270 2139.040 ;
        RECT 2899.450 2138.980 2899.770 2139.040 ;
      LAYER via ;
        RECT 1944.980 2138.980 1945.240 2139.240 ;
        RECT 2899.480 2138.980 2899.740 2139.240 ;
      LAYER met2 ;
        RECT 2899.470 2140.795 2899.750 2141.165 ;
        RECT 2899.540 2139.270 2899.680 2140.795 ;
        RECT 1944.980 2138.950 1945.240 2139.270 ;
        RECT 2899.480 2138.950 2899.740 2139.270 ;
        RECT 1945.040 2101.045 1945.180 2138.950 ;
        RECT 1941.290 2100.675 1941.570 2101.045 ;
        RECT 1944.970 2100.675 1945.250 2101.045 ;
        RECT 1941.360 2069.765 1941.500 2100.675 ;
        RECT 1941.290 2069.395 1941.570 2069.765 ;
        RECT 1942.670 2068.715 1942.950 2069.085 ;
        RECT 1942.740 1980.685 1942.880 2068.715 ;
        RECT 1941.750 1980.570 1942.030 1980.685 ;
        RECT 1940.900 1980.430 1942.030 1980.570 ;
        RECT 1940.900 1979.890 1941.040 1980.430 ;
        RECT 1941.750 1980.315 1942.030 1980.430 ;
        RECT 1942.670 1980.315 1942.950 1980.685 ;
        RECT 1940.900 1979.750 1941.960 1979.890 ;
        RECT 1941.820 1932.290 1941.960 1979.750 ;
        RECT 1941.360 1932.150 1941.960 1932.290 ;
        RECT 1941.360 1931.725 1941.500 1932.150 ;
        RECT 1941.290 1931.355 1941.570 1931.725 ;
        RECT 1943.130 1931.355 1943.410 1931.725 ;
        RECT 1943.200 1884.125 1943.340 1931.355 ;
        RECT 1941.750 1884.010 1942.030 1884.125 ;
        RECT 1940.900 1883.870 1942.030 1884.010 ;
        RECT 1940.900 1883.330 1941.040 1883.870 ;
        RECT 1941.750 1883.755 1942.030 1883.870 ;
        RECT 1943.130 1883.755 1943.410 1884.125 ;
        RECT 1940.900 1883.190 1941.960 1883.330 ;
        RECT 1941.820 1835.730 1941.960 1883.190 ;
        RECT 1941.360 1835.590 1941.960 1835.730 ;
        RECT 1941.360 1835.165 1941.500 1835.590 ;
        RECT 1941.290 1834.795 1941.570 1835.165 ;
        RECT 1941.290 1787.450 1941.570 1787.565 ;
        RECT 1940.900 1787.310 1941.570 1787.450 ;
        RECT 1940.900 1739.850 1941.040 1787.310 ;
        RECT 1941.290 1787.195 1941.570 1787.310 ;
        RECT 1941.290 1739.850 1941.570 1739.965 ;
        RECT 1940.900 1739.710 1941.570 1739.850 ;
        RECT 1941.290 1739.595 1941.570 1739.710 ;
        RECT 1942.210 1738.915 1942.490 1739.285 ;
        RECT 1942.280 1704.490 1942.420 1738.915 ;
        RECT 1941.360 1704.350 1942.420 1704.490 ;
        RECT 1940.370 1703.810 1940.650 1704.000 ;
        RECT 1941.360 1703.810 1941.500 1704.350 ;
        RECT 1940.370 1703.670 1941.500 1703.810 ;
        RECT 1940.370 1700.000 1940.650 1703.670 ;
      LAYER via2 ;
        RECT 2899.470 2140.840 2899.750 2141.120 ;
        RECT 1941.290 2100.720 1941.570 2101.000 ;
        RECT 1944.970 2100.720 1945.250 2101.000 ;
        RECT 1941.290 2069.440 1941.570 2069.720 ;
        RECT 1942.670 2068.760 1942.950 2069.040 ;
        RECT 1941.750 1980.360 1942.030 1980.640 ;
        RECT 1942.670 1980.360 1942.950 1980.640 ;
        RECT 1941.290 1931.400 1941.570 1931.680 ;
        RECT 1943.130 1931.400 1943.410 1931.680 ;
        RECT 1941.750 1883.800 1942.030 1884.080 ;
        RECT 1943.130 1883.800 1943.410 1884.080 ;
        RECT 1941.290 1834.840 1941.570 1835.120 ;
        RECT 1941.290 1787.240 1941.570 1787.520 ;
        RECT 1941.290 1739.640 1941.570 1739.920 ;
        RECT 1942.210 1738.960 1942.490 1739.240 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 2140.380 2924.800 2141.580 ;
=======
        RECT 2900.825 2141.130 2901.155 2141.145 ;
=======
        RECT 2899.445 2141.130 2899.775 2141.145 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 2141.130 2924.800 2141.580 ;
        RECT 2899.445 2140.830 2924.800 2141.130 ;
        RECT 2899.445 2140.815 2899.775 2140.830 ;
        RECT 2917.600 2140.380 2924.800 2140.830 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1941.265 2101.010 1941.595 2101.025 ;
        RECT 1944.945 2101.010 1945.275 2101.025 ;
        RECT 1941.265 2100.710 1945.275 2101.010 ;
        RECT 1941.265 2100.695 1941.595 2100.710 ;
        RECT 1944.945 2100.695 1945.275 2100.710 ;
        RECT 1941.265 2069.415 1941.595 2069.745 ;
        RECT 1941.280 2069.050 1941.580 2069.415 ;
        RECT 1942.645 2069.050 1942.975 2069.065 ;
        RECT 1941.280 2068.750 1942.975 2069.050 ;
        RECT 1942.645 2068.735 1942.975 2068.750 ;
        RECT 1941.725 1980.650 1942.055 1980.665 ;
        RECT 1942.645 1980.650 1942.975 1980.665 ;
        RECT 1941.725 1980.350 1942.975 1980.650 ;
        RECT 1941.725 1980.335 1942.055 1980.350 ;
        RECT 1942.645 1980.335 1942.975 1980.350 ;
        RECT 1941.265 1931.690 1941.595 1931.705 ;
        RECT 1943.105 1931.690 1943.435 1931.705 ;
        RECT 1941.265 1931.390 1943.435 1931.690 ;
        RECT 1941.265 1931.375 1941.595 1931.390 ;
        RECT 1943.105 1931.375 1943.435 1931.390 ;
        RECT 1941.725 1884.090 1942.055 1884.105 ;
        RECT 1943.105 1884.090 1943.435 1884.105 ;
        RECT 1941.725 1883.790 1943.435 1884.090 ;
        RECT 1941.725 1883.775 1942.055 1883.790 ;
        RECT 1943.105 1883.775 1943.435 1883.790 ;
        RECT 1941.265 1835.130 1941.595 1835.145 ;
        RECT 1941.265 1834.815 1941.810 1835.130 ;
        RECT 1941.510 1834.460 1941.810 1834.815 ;
        RECT 1941.470 1834.140 1941.850 1834.460 ;
        RECT 1941.470 1787.900 1941.850 1788.220 ;
        RECT 1941.510 1787.545 1941.810 1787.900 ;
        RECT 1941.265 1787.230 1941.810 1787.545 ;
        RECT 1941.265 1787.215 1941.595 1787.230 ;
        RECT 1941.265 1739.930 1941.595 1739.945 ;
        RECT 1941.265 1739.630 1942.730 1739.930 ;
        RECT 1941.265 1739.615 1941.595 1739.630 ;
        RECT 1942.430 1739.265 1942.730 1739.630 ;
        RECT 1942.185 1738.950 1942.730 1739.265 ;
        RECT 1942.185 1738.935 1942.515 1738.950 ;
      LAYER via3 ;
        RECT 1941.500 1834.140 1941.820 1834.460 ;
        RECT 1941.500 1787.900 1941.820 1788.220 ;
      LAYER met4 ;
        RECT 1941.495 1834.135 1941.825 1834.465 ;
        RECT 1941.510 1788.225 1941.810 1834.135 ;
        RECT 1941.495 1787.895 1941.825 1788.225 ;
>>>>>>> re-updated local openlane
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1606.390 84.560 1606.710 84.620 ;
        RECT 1618.350 84.560 1618.670 84.620 ;
        RECT 1606.390 84.420 1618.670 84.560 ;
        RECT 1606.390 84.360 1606.710 84.420 ;
        RECT 1618.350 84.360 1618.670 84.420 ;
        RECT 1799.130 84.220 1799.450 84.280 ;
        RECT 1806.490 84.220 1806.810 84.280 ;
        RECT 1799.130 84.080 1806.810 84.220 ;
        RECT 1799.130 84.020 1799.450 84.080 ;
        RECT 1806.490 84.020 1806.810 84.080 ;
        RECT 1932.070 84.220 1932.390 84.280 ;
        RECT 1946.330 84.220 1946.650 84.280 ;
        RECT 1932.070 84.080 1946.650 84.220 ;
        RECT 1932.070 84.020 1932.390 84.080 ;
        RECT 1946.330 84.020 1946.650 84.080 ;
        RECT 2608.730 84.220 2609.050 84.280 ;
        RECT 2632.650 84.220 2632.970 84.280 ;
        RECT 2608.730 84.080 2632.970 84.220 ;
        RECT 2608.730 84.020 2609.050 84.080 ;
        RECT 2632.650 84.020 2632.970 84.080 ;
        RECT 1435.730 83.880 1436.050 83.940 ;
        RECT 1490.010 83.880 1490.330 83.940 ;
        RECT 1435.730 83.740 1490.330 83.880 ;
        RECT 1435.730 83.680 1436.050 83.740 ;
        RECT 1490.010 83.680 1490.330 83.740 ;
        RECT 1642.270 83.540 1642.590 83.600 ;
        RECT 1690.110 83.540 1690.430 83.600 ;
        RECT 1642.270 83.400 1690.430 83.540 ;
        RECT 1642.270 83.340 1642.590 83.400 ;
        RECT 1690.110 83.340 1690.430 83.400 ;
      LAYER via ;
        RECT 1606.420 84.360 1606.680 84.620 ;
        RECT 1618.380 84.360 1618.640 84.620 ;
        RECT 1799.160 84.020 1799.420 84.280 ;
        RECT 1806.520 84.020 1806.780 84.280 ;
        RECT 1932.100 84.020 1932.360 84.280 ;
        RECT 1946.360 84.020 1946.620 84.280 ;
        RECT 2608.760 84.020 2609.020 84.280 ;
        RECT 2632.680 84.020 2632.940 84.280 ;
        RECT 1435.760 83.680 1436.020 83.940 ;
        RECT 1490.040 83.680 1490.300 83.940 ;
        RECT 1642.300 83.340 1642.560 83.600 ;
        RECT 1690.140 83.340 1690.400 83.600 ;
      LAYER met2 ;
        RECT 1153.310 2498.050 1153.590 2500.000 ;
        RECT 1155.150 2498.050 1155.430 2498.165 ;
        RECT 1153.310 2497.910 1155.430 2498.050 ;
        RECT 1153.310 2496.000 1153.590 2497.910 ;
        RECT 1155.150 2497.795 1155.430 2497.910 ;
        RECT 1946.350 85.155 1946.630 85.525 ;
        RECT 1993.730 85.155 1994.010 85.525 ;
        RECT 2268.810 85.155 2269.090 85.525 ;
        RECT 1606.410 84.475 1606.690 84.845 ;
        RECT 1606.420 84.330 1606.680 84.475 ;
        RECT 1618.380 84.330 1618.640 84.650 ;
        RECT 1690.130 84.475 1690.410 84.845 ;
        RECT 1435.750 83.795 1436.030 84.165 ;
        RECT 1511.650 84.050 1511.930 84.165 ;
        RECT 1435.760 83.650 1436.020 83.795 ;
        RECT 1490.040 83.650 1490.300 83.970 ;
        RECT 1510.800 83.910 1511.930 84.050 ;
        RECT 1490.100 83.485 1490.240 83.650 ;
        RECT 1510.800 83.485 1510.940 83.910 ;
        RECT 1511.650 83.795 1511.930 83.910 ;
        RECT 1618.440 83.485 1618.580 84.330 ;
        RECT 1690.200 83.630 1690.340 84.475 ;
        RECT 1946.420 84.310 1946.560 85.155 ;
        RECT 1993.800 84.730 1993.940 85.155 ;
        RECT 1994.650 84.730 1994.930 84.845 ;
        RECT 1993.800 84.590 1994.930 84.730 ;
        RECT 1994.650 84.475 1994.930 84.590 ;
        RECT 2069.630 84.475 2069.910 84.845 ;
        RECT 2076.530 84.475 2076.810 84.845 ;
        RECT 1799.160 84.165 1799.420 84.310 ;
        RECT 1806.520 84.165 1806.780 84.310 ;
        RECT 1932.100 84.165 1932.360 84.310 ;
        RECT 1799.150 83.795 1799.430 84.165 ;
        RECT 1806.510 83.795 1806.790 84.165 ;
        RECT 1932.090 83.795 1932.370 84.165 ;
        RECT 1946.360 83.990 1946.620 84.310 ;
        RECT 1642.300 83.485 1642.560 83.630 ;
        RECT 1490.030 83.115 1490.310 83.485 ;
        RECT 1510.730 83.115 1511.010 83.485 ;
        RECT 1618.370 83.115 1618.650 83.485 ;
        RECT 1642.290 83.115 1642.570 83.485 ;
        RECT 1690.140 83.310 1690.400 83.630 ;
        RECT 2069.700 83.485 2069.840 84.475 ;
        RECT 2076.600 83.485 2076.740 84.475 ;
        RECT 2268.880 84.050 2269.020 85.155 ;
        RECT 2304.230 84.475 2304.510 84.845 ;
        RECT 2269.270 84.050 2269.550 84.165 ;
        RECT 2268.880 83.910 2269.550 84.050 ;
        RECT 2269.270 83.795 2269.550 83.910 ;
        RECT 2069.630 83.115 2069.910 83.485 ;
        RECT 2076.530 83.115 2076.810 83.485 ;
        RECT 2304.300 82.805 2304.440 84.475 ;
        RECT 2608.760 84.165 2609.020 84.310 ;
        RECT 2632.680 84.165 2632.940 84.310 ;
        RECT 2608.750 83.795 2609.030 84.165 ;
        RECT 2632.670 83.795 2632.950 84.165 ;
        RECT 2304.230 82.435 2304.510 82.805 ;
      LAYER via2 ;
        RECT 1155.150 2497.840 1155.430 2498.120 ;
        RECT 1946.350 85.200 1946.630 85.480 ;
        RECT 1993.730 85.200 1994.010 85.480 ;
        RECT 2268.810 85.200 2269.090 85.480 ;
        RECT 1606.410 84.520 1606.690 84.800 ;
        RECT 1690.130 84.520 1690.410 84.800 ;
        RECT 1435.750 83.840 1436.030 84.120 ;
        RECT 1511.650 83.840 1511.930 84.120 ;
        RECT 1994.650 84.520 1994.930 84.800 ;
        RECT 2069.630 84.520 2069.910 84.800 ;
        RECT 2076.530 84.520 2076.810 84.800 ;
        RECT 1799.150 83.840 1799.430 84.120 ;
        RECT 1806.510 83.840 1806.790 84.120 ;
        RECT 1932.090 83.840 1932.370 84.120 ;
        RECT 1490.030 83.160 1490.310 83.440 ;
        RECT 1510.730 83.160 1511.010 83.440 ;
        RECT 1618.370 83.160 1618.650 83.440 ;
        RECT 1642.290 83.160 1642.570 83.440 ;
        RECT 2304.230 84.520 2304.510 84.800 ;
        RECT 2269.270 83.840 2269.550 84.120 ;
        RECT 2069.630 83.160 2069.910 83.440 ;
        RECT 2076.530 83.160 2076.810 83.440 ;
        RECT 2608.750 83.840 2609.030 84.120 ;
        RECT 2632.670 83.840 2632.950 84.120 ;
        RECT 2304.230 82.480 2304.510 82.760 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 87.460 2924.800 88.660 ;
=======
        RECT 1155.125 2498.130 1155.455 2498.145 ;
        RECT 1158.550 2498.130 1158.930 2498.140 ;
        RECT 1155.125 2497.830 1158.930 2498.130 ;
        RECT 1155.125 2497.815 1155.455 2497.830 ;
        RECT 1158.550 2497.820 1158.930 2497.830 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2916.710 87.910 2924.800 88.210 ;
        RECT 1946.325 85.490 1946.655 85.505 ;
        RECT 1993.705 85.490 1994.035 85.505 ;
        RECT 2268.785 85.490 2269.115 85.505 ;
        RECT 1337.990 85.190 1339.210 85.490 ;
        RECT 1337.990 84.810 1338.290 85.190 ;
        RECT 1338.910 84.820 1339.210 85.190 ;
        RECT 1946.325 85.190 1994.035 85.490 ;
        RECT 1946.325 85.175 1946.655 85.190 ;
        RECT 1993.705 85.175 1994.035 85.190 ;
        RECT 2234.990 85.190 2269.115 85.490 ;
        RECT 1290.150 84.510 1338.290 84.810 ;
        RECT 1290.150 84.130 1290.450 84.510 ;
        RECT 1338.870 84.500 1339.250 84.820 ;
        RECT 1606.385 84.810 1606.715 84.825 ;
        RECT 1410.670 84.510 1435.810 84.810 ;
        RECT 1269.910 83.830 1290.450 84.130 ;
        RECT 1158.550 83.450 1158.930 83.460 ;
        RECT 1269.910 83.450 1270.210 83.830 ;
        RECT 1158.550 83.150 1270.210 83.450 ;
        RECT 1338.870 83.450 1339.250 83.460 ;
        RECT 1410.670 83.450 1410.970 84.510 ;
        RECT 1435.510 84.145 1435.810 84.510 ;
        RECT 1545.910 84.510 1606.715 84.810 ;
        RECT 1435.510 83.830 1436.055 84.145 ;
        RECT 1435.725 83.815 1436.055 83.830 ;
        RECT 1511.625 84.130 1511.955 84.145 ;
        RECT 1545.910 84.130 1546.210 84.510 ;
        RECT 1606.385 84.495 1606.715 84.510 ;
        RECT 1690.105 84.810 1690.435 84.825 ;
        RECT 1883.510 84.810 1883.890 84.820 ;
        RECT 1690.105 84.510 1704.450 84.810 ;
        RECT 1690.105 84.495 1690.435 84.510 ;
        RECT 1511.625 83.830 1546.210 84.130 ;
        RECT 1511.625 83.815 1511.955 83.830 ;
        RECT 1338.870 83.150 1410.970 83.450 ;
        RECT 1490.005 83.450 1490.335 83.465 ;
        RECT 1510.705 83.450 1511.035 83.465 ;
        RECT 1490.005 83.150 1511.035 83.450 ;
        RECT 1158.550 83.140 1158.930 83.150 ;
        RECT 1338.870 83.140 1339.250 83.150 ;
        RECT 1490.005 83.135 1490.335 83.150 ;
        RECT 1510.705 83.135 1511.035 83.150 ;
        RECT 1618.345 83.450 1618.675 83.465 ;
        RECT 1642.265 83.450 1642.595 83.465 ;
        RECT 1618.345 83.150 1642.595 83.450 ;
        RECT 1704.150 83.450 1704.450 84.510 ;
        RECT 1849.510 84.510 1883.890 84.810 ;
        RECT 1799.125 84.130 1799.455 84.145 ;
        RECT 1752.910 83.830 1799.455 84.130 ;
        RECT 1752.910 83.450 1753.210 83.830 ;
        RECT 1799.125 83.815 1799.455 83.830 ;
        RECT 1806.485 84.130 1806.815 84.145 ;
        RECT 1806.485 83.830 1835.090 84.130 ;
        RECT 1806.485 83.815 1806.815 83.830 ;
        RECT 1704.150 83.150 1753.210 83.450 ;
        RECT 1834.790 83.450 1835.090 83.830 ;
        RECT 1849.510 83.450 1849.810 84.510 ;
        RECT 1883.510 84.500 1883.890 84.510 ;
        RECT 1994.625 84.810 1994.955 84.825 ;
        RECT 2069.605 84.810 2069.935 84.825 ;
        RECT 2076.505 84.810 2076.835 84.825 ;
        RECT 2234.990 84.810 2235.290 85.190 ;
        RECT 2268.785 85.175 2269.115 85.190 ;
        RECT 1994.625 84.510 2021.850 84.810 ;
        RECT 1994.625 84.495 1994.955 84.510 ;
        RECT 1932.065 84.130 1932.395 84.145 ;
        RECT 1834.790 83.150 1849.810 83.450 ;
        RECT 1931.390 83.830 1932.395 84.130 ;
        RECT 1618.345 83.135 1618.675 83.150 ;
        RECT 1642.265 83.135 1642.595 83.150 ;
        RECT 1883.510 82.770 1883.890 82.780 ;
        RECT 1931.390 82.770 1931.690 83.830 ;
        RECT 1932.065 83.815 1932.395 83.830 ;
        RECT 2021.550 83.450 2021.850 84.510 ;
        RECT 2069.605 84.510 2076.835 84.810 ;
        RECT 2069.605 84.495 2069.935 84.510 ;
        RECT 2076.505 84.495 2076.835 84.510 ;
        RECT 2089.630 84.510 2235.290 84.810 ;
        RECT 2304.205 84.810 2304.535 84.825 ;
        RECT 2304.205 84.510 2353.050 84.810 ;
        RECT 2069.605 83.450 2069.935 83.465 ;
        RECT 2021.550 83.150 2069.935 83.450 ;
        RECT 2069.605 83.135 2069.935 83.150 ;
        RECT 2076.505 83.450 2076.835 83.465 ;
        RECT 2089.630 83.450 2089.930 84.510 ;
        RECT 2304.205 84.495 2304.535 84.510 ;
        RECT 2269.245 84.130 2269.575 84.145 ;
        RECT 2269.910 84.130 2270.290 84.140 ;
        RECT 2269.245 83.830 2270.290 84.130 ;
        RECT 2352.750 84.130 2353.050 84.510 ;
        RECT 2669.230 84.510 2739.450 84.810 ;
        RECT 2572.630 84.130 2574.770 84.300 ;
        RECT 2608.725 84.130 2609.055 84.145 ;
        RECT 2352.750 83.830 2400.890 84.130 ;
        RECT 2269.245 83.815 2269.575 83.830 ;
        RECT 2269.910 83.820 2270.290 83.830 ;
        RECT 2076.505 83.150 2089.930 83.450 ;
        RECT 2400.590 83.450 2400.890 83.830 ;
        RECT 2429.110 83.830 2511.290 84.130 ;
        RECT 2429.110 83.450 2429.410 83.830 ;
        RECT 2400.590 83.150 2429.410 83.450 ;
        RECT 2510.990 83.450 2511.290 83.830 ;
        RECT 2559.750 84.000 2609.055 84.130 ;
        RECT 2559.750 83.830 2572.930 84.000 ;
        RECT 2574.470 83.830 2609.055 84.000 ;
        RECT 2559.750 83.450 2560.050 83.830 ;
        RECT 2608.725 83.815 2609.055 83.830 ;
        RECT 2632.645 84.130 2632.975 84.145 ;
        RECT 2669.230 84.130 2669.530 84.510 ;
        RECT 2632.645 83.830 2669.530 84.130 ;
        RECT 2739.150 84.130 2739.450 84.510 ;
        RECT 2787.910 84.510 2836.050 84.810 ;
        RECT 2739.150 83.830 2787.290 84.130 ;
        RECT 2632.645 83.815 2632.975 83.830 ;
        RECT 2510.990 83.150 2560.050 83.450 ;
        RECT 2786.990 83.450 2787.290 83.830 ;
        RECT 2787.910 83.450 2788.210 84.510 ;
        RECT 2835.750 84.130 2836.050 84.510 ;
        RECT 2916.710 84.130 2917.010 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
        RECT 2835.750 83.830 2883.890 84.130 ;
        RECT 2786.990 83.150 2788.210 83.450 ;
        RECT 2883.590 83.450 2883.890 83.830 ;
        RECT 2884.510 83.830 2917.010 84.130 ;
        RECT 2884.510 83.450 2884.810 83.830 ;
        RECT 2883.590 83.150 2884.810 83.450 ;
        RECT 2076.505 83.135 2076.835 83.150 ;
        RECT 1883.510 82.470 1931.690 82.770 ;
        RECT 2269.910 82.770 2270.290 82.780 ;
        RECT 2304.205 82.770 2304.535 82.785 ;
        RECT 2269.910 82.470 2304.535 82.770 ;
        RECT 1883.510 82.460 1883.890 82.470 ;
        RECT 2269.910 82.460 2270.290 82.470 ;
        RECT 2304.205 82.455 2304.535 82.470 ;
      LAYER via3 ;
        RECT 1158.580 2497.820 1158.900 2498.140 ;
        RECT 1338.900 84.500 1339.220 84.820 ;
        RECT 1158.580 83.140 1158.900 83.460 ;
        RECT 1338.900 83.140 1339.220 83.460 ;
        RECT 1883.540 84.500 1883.860 84.820 ;
        RECT 1883.540 82.460 1883.860 82.780 ;
        RECT 2269.940 83.820 2270.260 84.140 ;
        RECT 2269.940 82.460 2270.260 82.780 ;
      LAYER met4 ;
        RECT 1158.575 2497.815 1158.905 2498.145 ;
        RECT 1158.590 83.465 1158.890 2497.815 ;
        RECT 1338.895 84.495 1339.225 84.825 ;
        RECT 1883.535 84.495 1883.865 84.825 ;
        RECT 1338.910 83.465 1339.210 84.495 ;
        RECT 1158.575 83.135 1158.905 83.465 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1338.895 83.135 1339.225 83.465 ;
        RECT 1883.550 82.785 1883.850 84.495 ;
        RECT 2269.935 83.815 2270.265 84.145 ;
        RECT 2269.950 82.785 2270.250 83.815 ;
        RECT 1883.535 82.455 1883.865 82.785 ;
        RECT 2269.935 82.455 2270.265 82.785 ;
>>>>>>> re-updated local openlane
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1348.330 2499.240 1348.650 2499.300 ;
        RECT 2135.390 2499.240 2135.710 2499.300 ;
        RECT 1348.330 2499.100 2135.710 2499.240 ;
        RECT 1348.330 2499.040 1348.650 2499.100 ;
        RECT 2135.390 2499.040 2135.710 2499.100 ;
        RECT 2135.390 2435.660 2135.710 2435.720 ;
        RECT 2900.830 2435.660 2901.150 2435.720 ;
        RECT 2135.390 2435.520 2901.150 2435.660 ;
        RECT 2135.390 2435.460 2135.710 2435.520 ;
        RECT 2900.830 2435.460 2901.150 2435.520 ;
      LAYER via ;
        RECT 1348.360 2499.040 1348.620 2499.300 ;
        RECT 2135.420 2499.040 2135.680 2499.300 ;
        RECT 2135.420 2435.460 2135.680 2435.720 ;
        RECT 2900.860 2435.460 2901.120 2435.720 ;
      LAYER met2 ;
        RECT 1346.510 2499.410 1346.790 2500.000 ;
        RECT 1346.510 2499.330 1348.560 2499.410 ;
        RECT 1346.510 2499.270 1348.620 2499.330 ;
        RECT 1346.510 2496.000 1346.790 2499.270 ;
        RECT 1348.360 2499.010 1348.620 2499.270 ;
        RECT 2135.420 2499.010 2135.680 2499.330 ;
        RECT 2135.480 2435.750 2135.620 2499.010 ;
        RECT 2135.420 2435.430 2135.680 2435.750 ;
        RECT 2900.860 2435.430 2901.120 2435.750 ;
        RECT 2900.920 2434.245 2901.060 2435.430 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 2433.460 2924.800 2434.660 ;
=======
        RECT 2901.745 2434.210 2902.075 2434.225 ;
=======
        RECT 2900.825 2434.210 2901.155 2434.225 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1365.810 2663.800 1366.130 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 1365.810 2663.660 2901.150 2663.800 ;
        RECT 1365.810 2663.600 1366.130 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
      LAYER via ;
        RECT 1365.840 2663.600 1366.100 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 1365.840 2663.570 1366.100 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 1365.900 2500.000 1366.040 2663.570 ;
        RECT 1365.830 2496.000 1366.110 2500.000 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2668.740 2924.800 2669.940 ;
=======
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1386.510 2898.400 1386.830 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 1386.510 2898.260 2901.150 2898.400 ;
        RECT 1386.510 2898.200 1386.830 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
      LAYER via ;
        RECT 1386.540 2898.200 1386.800 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 1386.540 2898.170 1386.800 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 1385.150 2499.410 1385.430 2500.000 ;
        RECT 1386.600 2499.410 1386.740 2898.170 ;
        RECT 1385.150 2499.270 1386.740 2499.410 ;
        RECT 1385.150 2496.000 1385.430 2499.270 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2903.340 2924.800 2904.540 ;
=======
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1407.210 3133.000 1407.530 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 1407.210 3132.860 2901.150 3133.000 ;
        RECT 1407.210 3132.800 1407.530 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 1407.240 3132.800 1407.500 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 1407.240 3132.770 1407.500 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 1404.470 2498.730 1404.750 2500.000 ;
        RECT 1407.300 2498.730 1407.440 3132.770 ;
        RECT 1404.470 2498.590 1407.440 2498.730 ;
        RECT 1404.470 2496.000 1404.750 2498.590 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3137.940 2924.800 3139.140 ;
=======
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1427.910 3367.600 1428.230 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1427.910 3367.460 2901.150 3367.600 ;
        RECT 1427.910 3367.400 1428.230 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 1424.230 2515.900 1424.550 2515.960 ;
        RECT 1427.910 2515.900 1428.230 2515.960 ;
        RECT 1424.230 2515.760 1428.230 2515.900 ;
        RECT 1424.230 2515.700 1424.550 2515.760 ;
        RECT 1427.910 2515.700 1428.230 2515.760 ;
      LAYER via ;
        RECT 1427.940 3367.400 1428.200 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 1424.260 2515.700 1424.520 2515.960 ;
        RECT 1427.940 2515.700 1428.200 2515.960 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1427.940 3367.370 1428.200 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1428.000 2515.990 1428.140 3367.370 ;
        RECT 1424.260 2515.670 1424.520 2515.990 ;
        RECT 1427.940 2515.670 1428.200 2515.990 ;
        RECT 1424.320 2500.000 1424.460 2515.670 ;
        RECT 1424.250 2496.000 1424.530 2500.000 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3372.540 2924.800 3373.740 ;
=======
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3422.355 ;
        RECT 2795.565 3104.965 2795.735 3139.475 ;
        RECT 2796.945 2959.445 2797.115 3035.775 ;
        RECT 2795.105 2753.065 2795.275 2801.175 ;
      LAYER mcon ;
        RECT 2796.485 3422.185 2796.655 3422.355 ;
        RECT 2795.565 3139.305 2795.735 3139.475 ;
        RECT 2796.945 3035.605 2797.115 3035.775 ;
        RECT 2795.105 2801.005 2795.275 2801.175 ;
      LAYER met1 ;
        RECT 2795.490 3443.080 2795.810 3443.140 ;
        RECT 2798.250 3443.080 2798.570 3443.140 ;
        RECT 2795.490 3442.940 2798.570 3443.080 ;
        RECT 2795.490 3442.880 2795.810 3442.940 ;
        RECT 2798.250 3442.880 2798.570 3442.940 ;
        RECT 2795.030 3422.340 2795.350 3422.400 ;
        RECT 2796.425 3422.340 2796.715 3422.385 ;
        RECT 2795.030 3422.200 2796.715 3422.340 ;
        RECT 2795.030 3422.140 2795.350 3422.200 ;
        RECT 2796.425 3422.155 2796.715 3422.200 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.490 3139.460 2795.810 3139.520 ;
        RECT 2795.295 3139.320 2795.810 3139.460 ;
        RECT 2795.490 3139.260 2795.810 3139.320 ;
        RECT 2795.505 3105.120 2795.795 3105.165 ;
        RECT 2796.410 3105.120 2796.730 3105.180 ;
        RECT 2795.505 3104.980 2796.730 3105.120 ;
        RECT 2795.505 3104.935 2795.795 3104.980 ;
        RECT 2796.410 3104.920 2796.730 3104.980 ;
        RECT 2796.410 3056.640 2796.730 3056.900 ;
        RECT 2796.500 3056.160 2796.640 3056.640 ;
        RECT 2796.870 3056.160 2797.190 3056.220 ;
        RECT 2796.500 3056.020 2797.190 3056.160 ;
        RECT 2796.870 3055.960 2797.190 3056.020 ;
        RECT 2796.870 3035.760 2797.190 3035.820 ;
        RECT 2796.675 3035.620 2797.190 3035.760 ;
        RECT 2796.870 3035.560 2797.190 3035.620 ;
        RECT 2796.870 2959.600 2797.190 2959.660 ;
        RECT 2796.675 2959.460 2797.190 2959.600 ;
        RECT 2796.870 2959.400 2797.190 2959.460 ;
        RECT 2796.870 2912.340 2797.190 2912.400 ;
        RECT 2796.500 2912.200 2797.190 2912.340 ;
        RECT 2796.500 2911.720 2796.640 2912.200 ;
        RECT 2796.870 2912.140 2797.190 2912.200 ;
        RECT 2796.410 2911.460 2796.730 2911.720 ;
        RECT 2795.030 2815.580 2795.350 2815.840 ;
        RECT 2795.120 2815.160 2795.260 2815.580 ;
        RECT 2795.030 2814.900 2795.350 2815.160 ;
        RECT 2795.030 2801.160 2795.350 2801.220 ;
        RECT 2794.835 2801.020 2795.350 2801.160 ;
        RECT 2795.030 2800.960 2795.350 2801.020 ;
        RECT 2795.045 2753.220 2795.335 2753.265 ;
        RECT 2795.950 2753.220 2796.270 2753.280 ;
        RECT 2795.045 2753.080 2796.270 2753.220 ;
        RECT 2795.045 2753.035 2795.335 2753.080 ;
        RECT 2795.950 2753.020 2796.270 2753.080 ;
        RECT 2795.030 2718.200 2795.350 2718.260 ;
        RECT 2795.950 2718.200 2796.270 2718.260 ;
        RECT 2795.030 2718.060 2796.270 2718.200 ;
        RECT 2795.030 2718.000 2795.350 2718.060 ;
        RECT 2795.950 2718.000 2796.270 2718.060 ;
        RECT 2795.030 2670.260 2795.350 2670.320 ;
        RECT 2795.950 2670.260 2796.270 2670.320 ;
        RECT 2795.030 2670.120 2796.270 2670.260 ;
        RECT 2795.030 2670.060 2795.350 2670.120 ;
        RECT 2795.950 2670.060 2796.270 2670.120 ;
        RECT 2795.950 2622.120 2796.270 2622.380 ;
        RECT 2796.040 2621.980 2796.180 2622.120 ;
        RECT 2796.410 2621.980 2796.730 2622.040 ;
        RECT 2796.040 2621.840 2796.730 2621.980 ;
        RECT 2796.410 2621.780 2796.730 2621.840 ;
        RECT 2795.490 2560.100 2795.810 2560.160 ;
        RECT 2796.870 2560.100 2797.190 2560.160 ;
        RECT 2795.490 2559.960 2797.190 2560.100 ;
        RECT 2795.490 2559.900 2795.810 2559.960 ;
        RECT 2796.870 2559.900 2797.190 2559.960 ;
        RECT 1443.550 2516.240 1443.870 2516.300 ;
        RECT 1443.550 2516.100 1456.200 2516.240 ;
        RECT 1443.550 2516.040 1443.870 2516.100 ;
        RECT 1456.060 2515.900 1456.200 2516.100 ;
        RECT 2796.870 2515.900 2797.190 2515.960 ;
        RECT 1456.060 2515.760 2797.190 2515.900 ;
        RECT 2796.870 2515.700 2797.190 2515.760 ;
      LAYER via ;
        RECT 2795.520 3442.880 2795.780 3443.140 ;
        RECT 2798.280 3442.880 2798.540 3443.140 ;
        RECT 2795.060 3422.140 2795.320 3422.400 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.520 3139.260 2795.780 3139.520 ;
        RECT 2796.440 3104.920 2796.700 3105.180 ;
        RECT 2796.440 3056.640 2796.700 3056.900 ;
        RECT 2796.900 3055.960 2797.160 3056.220 ;
        RECT 2796.900 3035.560 2797.160 3035.820 ;
        RECT 2796.900 2959.400 2797.160 2959.660 ;
        RECT 2796.900 2912.140 2797.160 2912.400 ;
        RECT 2796.440 2911.460 2796.700 2911.720 ;
        RECT 2795.060 2815.580 2795.320 2815.840 ;
        RECT 2795.060 2814.900 2795.320 2815.160 ;
        RECT 2795.060 2800.960 2795.320 2801.220 ;
        RECT 2795.980 2753.020 2796.240 2753.280 ;
        RECT 2795.060 2718.000 2795.320 2718.260 ;
        RECT 2795.980 2718.000 2796.240 2718.260 ;
        RECT 2795.060 2670.060 2795.320 2670.320 ;
        RECT 2795.980 2670.060 2796.240 2670.320 ;
        RECT 2795.980 2622.120 2796.240 2622.380 ;
        RECT 2796.440 2621.780 2796.700 2622.040 ;
        RECT 2795.520 2559.900 2795.780 2560.160 ;
        RECT 2796.900 2559.900 2797.160 2560.160 ;
        RECT 1443.580 2516.040 1443.840 2516.300 ;
        RECT 2796.900 2515.700 2797.160 2515.960 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2798.130 3519.700 2798.690 3524.800 ;
=======
        RECT 2798.130 3517.600 2798.690 3524.800 ;
<<<<<<< HEAD
        RECT 2798.340 3501.990 2798.480 3517.600 ;
        RECT 1455.540 3501.670 1455.800 3501.990 ;
        RECT 2798.280 3501.670 2798.540 3501.990 ;
        RECT 1455.600 2514.970 1455.740 3501.670 ;
        RECT 1450.480 2514.650 1450.740 2514.970 ;
        RECT 1455.540 2514.650 1455.800 2514.970 ;
        RECT 1450.540 2500.000 1450.680 2514.650 ;
        RECT 1450.470 2496.000 1450.750 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2798.340 3443.170 2798.480 3517.600 ;
        RECT 2795.520 3442.850 2795.780 3443.170 ;
        RECT 2798.280 3442.850 2798.540 3443.170 ;
        RECT 2795.580 3429.650 2795.720 3442.850 ;
        RECT 2795.120 3429.510 2795.720 3429.650 ;
        RECT 2795.120 3422.430 2795.260 3429.510 ;
        RECT 2795.060 3422.110 2795.320 3422.430 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3236.450 2796.180 3298.270 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3139.550 2795.720 3152.750 ;
        RECT 2795.520 3139.230 2795.780 3139.550 ;
        RECT 2796.440 3104.890 2796.700 3105.210 ;
        RECT 2796.500 3056.930 2796.640 3104.890 ;
        RECT 2796.440 3056.610 2796.700 3056.930 ;
        RECT 2796.900 3055.930 2797.160 3056.250 ;
        RECT 2796.960 3035.850 2797.100 3055.930 ;
        RECT 2796.900 3035.530 2797.160 3035.850 ;
        RECT 2796.900 2959.370 2797.160 2959.690 ;
        RECT 2796.960 2912.430 2797.100 2959.370 ;
        RECT 2796.900 2912.110 2797.160 2912.430 ;
        RECT 2796.440 2911.430 2796.700 2911.750 ;
        RECT 2796.500 2863.210 2796.640 2911.430 ;
        RECT 2795.580 2863.070 2796.640 2863.210 ;
        RECT 2795.580 2849.610 2795.720 2863.070 ;
        RECT 2795.120 2849.470 2795.720 2849.610 ;
        RECT 2795.120 2815.870 2795.260 2849.470 ;
        RECT 2795.060 2815.550 2795.320 2815.870 ;
        RECT 2795.060 2814.870 2795.320 2815.190 ;
        RECT 2795.120 2801.250 2795.260 2814.870 ;
        RECT 2795.060 2800.930 2795.320 2801.250 ;
        RECT 2795.980 2752.990 2796.240 2753.310 ;
        RECT 2796.040 2718.290 2796.180 2752.990 ;
        RECT 2795.060 2717.970 2795.320 2718.290 ;
        RECT 2795.980 2717.970 2796.240 2718.290 ;
        RECT 2795.120 2670.350 2795.260 2717.970 ;
        RECT 2795.060 2670.030 2795.320 2670.350 ;
        RECT 2795.980 2670.030 2796.240 2670.350 ;
        RECT 2796.040 2622.410 2796.180 2670.030 ;
        RECT 2795.980 2622.090 2796.240 2622.410 ;
        RECT 2796.440 2621.750 2796.700 2622.070 ;
        RECT 2796.500 2608.325 2796.640 2621.750 ;
        RECT 2795.510 2607.955 2795.790 2608.325 ;
        RECT 2796.430 2607.955 2796.710 2608.325 ;
        RECT 2795.580 2560.190 2795.720 2607.955 ;
        RECT 2795.520 2559.870 2795.780 2560.190 ;
        RECT 2796.900 2559.870 2797.160 2560.190 ;
        RECT 1443.580 2516.010 1443.840 2516.330 ;
        RECT 1443.640 2500.000 1443.780 2516.010 ;
        RECT 2796.960 2515.990 2797.100 2559.870 ;
        RECT 2796.900 2515.670 2797.160 2515.990 ;
        RECT 1443.570 2496.000 1443.850 2500.000 ;
      LAYER via2 ;
        RECT 2795.510 2608.000 2795.790 2608.280 ;
        RECT 2796.430 2608.000 2796.710 2608.280 ;
      LAYER met3 ;
        RECT 2795.485 2608.290 2795.815 2608.305 ;
        RECT 2796.405 2608.290 2796.735 2608.305 ;
        RECT 2795.485 2607.990 2796.735 2608.290 ;
        RECT 2795.485 2607.975 2795.815 2607.990 ;
        RECT 2796.405 2607.975 2796.735 2607.990 ;
>>>>>>> re-updated local openlane
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
        RECT 2470.805 2815.285 2470.975 2849.455 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
        RECT 2470.805 2849.285 2470.975 2849.455 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 2981.020 2470.590 2981.080 ;
        RECT 2471.190 2981.020 2471.510 2981.080 ;
        RECT 2470.270 2980.880 2471.510 2981.020 ;
        RECT 2470.270 2980.820 2470.590 2980.880 ;
        RECT 2471.190 2980.820 2471.510 2980.880 ;
        RECT 2469.350 2946.340 2469.670 2946.400 ;
        RECT 2470.730 2946.340 2471.050 2946.400 ;
        RECT 2469.350 2946.200 2471.050 2946.340 ;
        RECT 2469.350 2946.140 2469.670 2946.200 ;
        RECT 2470.730 2946.140 2471.050 2946.200 ;
        RECT 2470.730 2849.440 2471.050 2849.500 ;
        RECT 2470.535 2849.300 2471.050 2849.440 ;
        RECT 2470.730 2849.240 2471.050 2849.300 ;
        RECT 2470.745 2815.440 2471.035 2815.485 ;
        RECT 2471.650 2815.440 2471.970 2815.500 ;
        RECT 2470.745 2815.300 2471.970 2815.440 ;
        RECT 2470.745 2815.255 2471.035 2815.300 ;
        RECT 2471.650 2815.240 2471.970 2815.300 ;
        RECT 2470.730 2753.220 2471.050 2753.280 ;
        RECT 2472.110 2753.220 2472.430 2753.280 ;
        RECT 2470.730 2753.080 2472.430 2753.220 ;
        RECT 2470.730 2753.020 2471.050 2753.080 ;
        RECT 2472.110 2753.020 2472.430 2753.080 ;
        RECT 2472.110 2719.220 2472.430 2719.280 ;
        RECT 2471.740 2719.080 2472.430 2719.220 ;
        RECT 2471.740 2718.600 2471.880 2719.080 ;
        RECT 2472.110 2719.020 2472.430 2719.080 ;
        RECT 2471.650 2718.340 2471.970 2718.600 ;
        RECT 2471.650 2670.400 2471.970 2670.660 ;
        RECT 2471.740 2669.920 2471.880 2670.400 ;
        RECT 2472.110 2669.920 2472.430 2669.980 ;
        RECT 2471.740 2669.780 2472.430 2669.920 ;
        RECT 2472.110 2669.720 2472.430 2669.780 ;
        RECT 2472.110 2649.520 2472.430 2649.580 ;
        RECT 2473.030 2649.520 2473.350 2649.580 ;
        RECT 2472.110 2649.380 2473.350 2649.520 ;
        RECT 2472.110 2649.320 2472.430 2649.380 ;
        RECT 2473.030 2649.320 2473.350 2649.380 ;
        RECT 2472.110 2573.360 2472.430 2573.420 ;
        RECT 2473.030 2573.360 2473.350 2573.420 ;
        RECT 2472.110 2573.220 2473.350 2573.360 ;
        RECT 2472.110 2573.160 2472.430 2573.220 ;
        RECT 2473.030 2573.160 2473.350 2573.220 ;
        RECT 1462.870 2516.240 1463.190 2516.300 ;
        RECT 2472.110 2516.240 2472.430 2516.300 ;
        RECT 1462.870 2516.100 2472.430 2516.240 ;
        RECT 1462.870 2516.040 1463.190 2516.100 ;
        RECT 2472.110 2516.040 2472.430 2516.100 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 2980.820 2470.560 2981.080 ;
        RECT 2471.220 2980.820 2471.480 2981.080 ;
        RECT 2469.380 2946.140 2469.640 2946.400 ;
        RECT 2470.760 2946.140 2471.020 2946.400 ;
        RECT 2470.760 2849.240 2471.020 2849.500 ;
        RECT 2471.680 2815.240 2471.940 2815.500 ;
        RECT 2470.760 2753.020 2471.020 2753.280 ;
        RECT 2472.140 2753.020 2472.400 2753.280 ;
        RECT 2472.140 2719.020 2472.400 2719.280 ;
        RECT 2471.680 2718.340 2471.940 2718.600 ;
        RECT 2471.680 2670.400 2471.940 2670.660 ;
        RECT 2472.140 2669.720 2472.400 2669.980 ;
        RECT 2472.140 2649.320 2472.400 2649.580 ;
        RECT 2473.060 2649.320 2473.320 2649.580 ;
        RECT 2472.140 2573.160 2472.400 2573.420 ;
        RECT 2473.060 2573.160 2473.320 2573.420 ;
        RECT 1462.900 2516.040 1463.160 2516.300 ;
        RECT 2472.140 2516.040 2472.400 2516.300 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2473.830 3519.700 2474.390 3524.800 ;
=======
        RECT 2473.830 3517.600 2474.390 3524.800 ;
<<<<<<< HEAD
        RECT 2474.040 3503.690 2474.180 3517.600 ;
        RECT 1476.240 3503.370 1476.500 3503.690 ;
        RECT 2473.980 3503.370 2474.240 3503.690 ;
        RECT 1476.300 2514.970 1476.440 3503.370 ;
        RECT 1470.260 2514.650 1470.520 2514.970 ;
        RECT 1476.240 2514.650 1476.500 2514.970 ;
        RECT 1470.320 2500.000 1470.460 2514.650 ;
        RECT 1470.250 2496.000 1470.530 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3430.445 2474.640 3517.230 ;
        RECT 2474.430 3430.075 2474.710 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3298.410 2470.960 3332.690 ;
        RECT 2470.820 3298.270 2471.420 3298.410 ;
        RECT 2471.280 3270.790 2471.420 3298.270 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3222.250 2470.500 3270.470 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 2981.110 2471.420 3125.550 ;
        RECT 2470.300 2980.850 2470.560 2981.110 ;
        RECT 2470.300 2980.790 2470.960 2980.850 ;
        RECT 2471.220 2980.790 2471.480 2981.110 ;
        RECT 2470.360 2980.710 2470.960 2980.790 ;
        RECT 2470.820 2980.170 2470.960 2980.710 ;
        RECT 2470.820 2980.030 2471.420 2980.170 ;
        RECT 2471.280 2959.770 2471.420 2980.030 ;
        RECT 2470.820 2959.630 2471.420 2959.770 ;
        RECT 2470.820 2946.430 2470.960 2959.630 ;
        RECT 2469.380 2946.110 2469.640 2946.430 ;
        RECT 2470.760 2946.110 2471.020 2946.430 ;
        RECT 2469.440 2898.685 2469.580 2946.110 ;
        RECT 2469.370 2898.315 2469.650 2898.685 ;
        RECT 2470.290 2898.315 2470.570 2898.685 ;
        RECT 2470.360 2863.210 2470.500 2898.315 ;
        RECT 2470.360 2863.070 2470.960 2863.210 ;
        RECT 2470.820 2849.530 2470.960 2863.070 ;
        RECT 2470.760 2849.210 2471.020 2849.530 ;
        RECT 2471.680 2815.210 2471.940 2815.530 ;
        RECT 2471.740 2801.445 2471.880 2815.210 ;
        RECT 2470.750 2801.075 2471.030 2801.445 ;
        RECT 2471.670 2801.075 2471.950 2801.445 ;
        RECT 2470.820 2753.310 2470.960 2801.075 ;
        RECT 2470.760 2752.990 2471.020 2753.310 ;
        RECT 2472.140 2752.990 2472.400 2753.310 ;
        RECT 2472.200 2719.310 2472.340 2752.990 ;
        RECT 2472.140 2718.990 2472.400 2719.310 ;
        RECT 2471.680 2718.310 2471.940 2718.630 ;
        RECT 2471.740 2670.690 2471.880 2718.310 ;
        RECT 2471.680 2670.370 2471.940 2670.690 ;
        RECT 2472.140 2669.690 2472.400 2670.010 ;
        RECT 2472.200 2649.610 2472.340 2669.690 ;
        RECT 2472.140 2649.290 2472.400 2649.610 ;
        RECT 2473.060 2649.290 2473.320 2649.610 ;
        RECT 2473.120 2573.450 2473.260 2649.290 ;
        RECT 2472.140 2573.130 2472.400 2573.450 ;
        RECT 2473.060 2573.130 2473.320 2573.450 ;
        RECT 2472.200 2516.330 2472.340 2573.130 ;
        RECT 1462.900 2516.010 1463.160 2516.330 ;
        RECT 2472.140 2516.010 2472.400 2516.330 ;
        RECT 1462.960 2500.000 1463.100 2516.010 ;
        RECT 1462.890 2496.000 1463.170 2500.000 ;
      LAYER via2 ;
        RECT 2474.430 3430.120 2474.710 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
        RECT 2469.370 2898.360 2469.650 2898.640 ;
        RECT 2470.290 2898.360 2470.570 2898.640 ;
        RECT 2470.750 2801.120 2471.030 2801.400 ;
        RECT 2471.670 2801.120 2471.950 2801.400 ;
      LAYER met3 ;
        RECT 2474.405 3430.410 2474.735 3430.425 ;
        RECT 2470.510 3430.110 2474.735 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.405 3430.095 2474.735 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
        RECT 2469.345 2898.650 2469.675 2898.665 ;
        RECT 2470.265 2898.650 2470.595 2898.665 ;
        RECT 2469.345 2898.350 2470.595 2898.650 ;
        RECT 2469.345 2898.335 2469.675 2898.350 ;
        RECT 2470.265 2898.335 2470.595 2898.350 ;
        RECT 2470.725 2801.410 2471.055 2801.425 ;
        RECT 2471.645 2801.410 2471.975 2801.425 ;
        RECT 2470.725 2801.110 2471.975 2801.410 ;
        RECT 2470.725 2801.095 2471.055 2801.110 ;
        RECT 2471.645 2801.095 2471.975 2801.110 ;
>>>>>>> re-updated local openlane
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3422.355 ;
        RECT 2146.965 3104.965 2147.135 3139.475 ;
        RECT 2146.505 2753.065 2146.675 2801.175 ;
      LAYER mcon ;
        RECT 2147.885 3422.185 2148.055 3422.355 ;
        RECT 2146.965 3139.305 2147.135 3139.475 ;
        RECT 2146.505 2801.005 2146.675 2801.175 ;
      LAYER met1 ;
        RECT 2146.890 3443.080 2147.210 3443.140 ;
        RECT 2149.190 3443.080 2149.510 3443.140 ;
        RECT 2146.890 3442.940 2149.510 3443.080 ;
        RECT 2146.890 3442.880 2147.210 3442.940 ;
        RECT 2149.190 3442.880 2149.510 3442.940 ;
        RECT 2146.430 3422.340 2146.750 3422.400 ;
        RECT 2147.825 3422.340 2148.115 3422.385 ;
        RECT 2146.430 3422.200 2148.115 3422.340 ;
        RECT 2146.430 3422.140 2146.750 3422.200 ;
        RECT 2147.825 3422.155 2148.115 3422.200 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2146.890 3139.460 2147.210 3139.520 ;
        RECT 2146.695 3139.320 2147.210 3139.460 ;
        RECT 2146.890 3139.260 2147.210 3139.320 ;
        RECT 2146.905 3105.120 2147.195 3105.165 ;
        RECT 2147.810 3105.120 2148.130 3105.180 ;
        RECT 2146.905 3104.980 2148.130 3105.120 ;
        RECT 2146.905 3104.935 2147.195 3104.980 ;
        RECT 2147.810 3104.920 2148.130 3104.980 ;
        RECT 2147.810 3056.640 2148.130 3056.900 ;
        RECT 2147.900 3056.160 2148.040 3056.640 ;
        RECT 2148.270 3056.160 2148.590 3056.220 ;
        RECT 2147.900 3056.020 2148.590 3056.160 ;
        RECT 2148.270 3055.960 2148.590 3056.020 ;
        RECT 2148.270 2912.340 2148.590 2912.400 ;
        RECT 2147.900 2912.200 2148.590 2912.340 ;
        RECT 2147.900 2911.720 2148.040 2912.200 ;
        RECT 2148.270 2912.140 2148.590 2912.200 ;
        RECT 2147.810 2911.460 2148.130 2911.720 ;
        RECT 2146.430 2815.580 2146.750 2815.840 ;
        RECT 2146.520 2815.160 2146.660 2815.580 ;
        RECT 2146.430 2814.900 2146.750 2815.160 ;
        RECT 2146.430 2801.160 2146.750 2801.220 ;
        RECT 2146.235 2801.020 2146.750 2801.160 ;
        RECT 2146.430 2800.960 2146.750 2801.020 ;
        RECT 2146.445 2753.220 2146.735 2753.265 ;
        RECT 2147.350 2753.220 2147.670 2753.280 ;
        RECT 2146.445 2753.080 2147.670 2753.220 ;
        RECT 2146.445 2753.035 2146.735 2753.080 ;
        RECT 2147.350 2753.020 2147.670 2753.080 ;
        RECT 2146.430 2718.200 2146.750 2718.260 ;
        RECT 2147.350 2718.200 2147.670 2718.260 ;
        RECT 2146.430 2718.060 2147.670 2718.200 ;
        RECT 2146.430 2718.000 2146.750 2718.060 ;
        RECT 2147.350 2718.000 2147.670 2718.060 ;
        RECT 2146.430 2670.260 2146.750 2670.320 ;
        RECT 2147.350 2670.260 2147.670 2670.320 ;
        RECT 2146.430 2670.120 2147.670 2670.260 ;
        RECT 2146.430 2670.060 2146.750 2670.120 ;
        RECT 2147.350 2670.060 2147.670 2670.120 ;
        RECT 2147.350 2622.120 2147.670 2622.380 ;
        RECT 2147.440 2621.980 2147.580 2622.120 ;
        RECT 2147.810 2621.980 2148.130 2622.040 ;
        RECT 2147.440 2621.840 2148.130 2621.980 ;
        RECT 2147.810 2621.780 2148.130 2621.840 ;
        RECT 2146.890 2560.100 2147.210 2560.160 ;
        RECT 2148.270 2560.100 2148.590 2560.160 ;
        RECT 2146.890 2559.960 2148.590 2560.100 ;
        RECT 2146.890 2559.900 2147.210 2559.960 ;
        RECT 2148.270 2559.900 2148.590 2559.960 ;
        RECT 1482.190 2516.580 1482.510 2516.640 ;
        RECT 2148.270 2516.580 2148.590 2516.640 ;
        RECT 1482.190 2516.440 2148.590 2516.580 ;
        RECT 1482.190 2516.380 1482.510 2516.440 ;
        RECT 2148.270 2516.380 2148.590 2516.440 ;
      LAYER via ;
        RECT 2146.920 3442.880 2147.180 3443.140 ;
        RECT 2149.220 3442.880 2149.480 3443.140 ;
        RECT 2146.460 3422.140 2146.720 3422.400 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.920 3139.260 2147.180 3139.520 ;
        RECT 2147.840 3104.920 2148.100 3105.180 ;
        RECT 2147.840 3056.640 2148.100 3056.900 ;
        RECT 2148.300 3055.960 2148.560 3056.220 ;
        RECT 2148.300 2912.140 2148.560 2912.400 ;
        RECT 2147.840 2911.460 2148.100 2911.720 ;
        RECT 2146.460 2815.580 2146.720 2815.840 ;
        RECT 2146.460 2814.900 2146.720 2815.160 ;
        RECT 2146.460 2800.960 2146.720 2801.220 ;
        RECT 2147.380 2753.020 2147.640 2753.280 ;
        RECT 2146.460 2718.000 2146.720 2718.260 ;
        RECT 2147.380 2718.000 2147.640 2718.260 ;
        RECT 2146.460 2670.060 2146.720 2670.320 ;
        RECT 2147.380 2670.060 2147.640 2670.320 ;
        RECT 2147.380 2622.120 2147.640 2622.380 ;
        RECT 2147.840 2621.780 2148.100 2622.040 ;
        RECT 2146.920 2559.900 2147.180 2560.160 ;
        RECT 2148.300 2559.900 2148.560 2560.160 ;
        RECT 1482.220 2516.380 1482.480 2516.640 ;
        RECT 2148.300 2516.380 2148.560 2516.640 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2149.070 3519.700 2149.630 3524.800 ;
=======
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3443.170 2149.420 3517.600 ;
        RECT 2146.920 3442.850 2147.180 3443.170 ;
        RECT 2149.220 3442.850 2149.480 3443.170 ;
        RECT 2146.980 3429.650 2147.120 3442.850 ;
        RECT 2146.520 3429.510 2147.120 3429.650 ;
        RECT 2146.520 3422.430 2146.660 3429.510 ;
        RECT 2146.460 3422.110 2146.720 3422.430 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3236.450 2147.580 3298.270 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3139.550 2147.120 3152.750 ;
        RECT 2146.920 3139.230 2147.180 3139.550 ;
        RECT 2147.840 3104.890 2148.100 3105.210 ;
        RECT 2147.900 3056.930 2148.040 3104.890 ;
        RECT 2147.840 3056.610 2148.100 3056.930 ;
        RECT 2148.300 3055.930 2148.560 3056.250 ;
        RECT 2148.360 3036.045 2148.500 3055.930 ;
        RECT 2148.290 3035.675 2148.570 3036.045 ;
        RECT 2148.290 2959.515 2148.570 2959.885 ;
        RECT 2148.360 2912.430 2148.500 2959.515 ;
        RECT 2148.300 2912.110 2148.560 2912.430 ;
        RECT 2147.840 2911.430 2148.100 2911.750 ;
        RECT 2147.900 2863.210 2148.040 2911.430 ;
        RECT 2146.980 2863.070 2148.040 2863.210 ;
        RECT 2146.980 2849.610 2147.120 2863.070 ;
        RECT 2146.520 2849.470 2147.120 2849.610 ;
        RECT 2146.520 2815.870 2146.660 2849.470 ;
        RECT 2146.460 2815.550 2146.720 2815.870 ;
        RECT 2146.460 2814.870 2146.720 2815.190 ;
        RECT 2146.520 2801.250 2146.660 2814.870 ;
        RECT 2146.460 2800.930 2146.720 2801.250 ;
        RECT 2147.380 2752.990 2147.640 2753.310 ;
        RECT 2147.440 2718.290 2147.580 2752.990 ;
        RECT 2146.460 2717.970 2146.720 2718.290 ;
        RECT 2147.380 2717.970 2147.640 2718.290 ;
        RECT 2146.520 2670.350 2146.660 2717.970 ;
        RECT 2146.460 2670.030 2146.720 2670.350 ;
        RECT 2147.380 2670.030 2147.640 2670.350 ;
        RECT 2147.440 2622.410 2147.580 2670.030 ;
        RECT 2147.380 2622.090 2147.640 2622.410 ;
        RECT 2147.840 2621.750 2148.100 2622.070 ;
        RECT 2147.900 2608.325 2148.040 2621.750 ;
        RECT 2146.910 2607.955 2147.190 2608.325 ;
        RECT 2147.830 2607.955 2148.110 2608.325 ;
        RECT 2146.980 2560.190 2147.120 2607.955 ;
        RECT 2146.920 2559.870 2147.180 2560.190 ;
        RECT 2148.300 2559.870 2148.560 2560.190 ;
        RECT 2148.360 2516.670 2148.500 2559.870 ;
        RECT 1482.220 2516.350 1482.480 2516.670 ;
        RECT 2148.300 2516.350 2148.560 2516.670 ;
        RECT 1482.280 2500.000 1482.420 2516.350 ;
        RECT 1482.210 2496.000 1482.490 2500.000 ;
      LAYER via2 ;
        RECT 2148.290 3035.720 2148.570 3036.000 ;
        RECT 2148.290 2959.560 2148.570 2959.840 ;
        RECT 2146.910 2608.000 2147.190 2608.280 ;
        RECT 2147.830 2608.000 2148.110 2608.280 ;
      LAYER met3 ;
        RECT 2147.550 3036.010 2147.930 3036.020 ;
        RECT 2148.265 3036.010 2148.595 3036.025 ;
        RECT 2147.550 3035.710 2148.595 3036.010 ;
        RECT 2147.550 3035.700 2147.930 3035.710 ;
        RECT 2148.265 3035.695 2148.595 3035.710 ;
        RECT 2147.550 2959.850 2147.930 2959.860 ;
        RECT 2148.265 2959.850 2148.595 2959.865 ;
        RECT 2147.550 2959.550 2148.595 2959.850 ;
        RECT 2147.550 2959.540 2147.930 2959.550 ;
        RECT 2148.265 2959.535 2148.595 2959.550 ;
        RECT 2146.885 2608.290 2147.215 2608.305 ;
        RECT 2147.805 2608.290 2148.135 2608.305 ;
        RECT 2146.885 2607.990 2148.135 2608.290 ;
        RECT 2146.885 2607.975 2147.215 2607.990 ;
        RECT 2147.805 2607.975 2148.135 2607.990 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via3 ;
        RECT 2147.580 3035.700 2147.900 3036.020 ;
        RECT 2147.580 2959.540 2147.900 2959.860 ;
      LAYER met4 ;
        RECT 2147.575 3035.695 2147.905 3036.025 ;
        RECT 2147.590 2959.865 2147.890 3035.695 ;
        RECT 2147.575 2959.535 2147.905 2959.865 ;
>>>>>>> re-updated local openlane
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1821.745 3332.765 1821.915 3380.875 ;
        RECT 1822.205 2815.285 1822.375 2849.455 ;
      LAYER mcon ;
        RECT 1821.745 3380.705 1821.915 3380.875 ;
        RECT 1822.205 2849.285 1822.375 2849.455 ;
      LAYER met1 ;
        RECT 1821.670 3380.860 1821.990 3380.920 ;
        RECT 1821.475 3380.720 1821.990 3380.860 ;
        RECT 1821.670 3380.660 1821.990 3380.720 ;
        RECT 1821.685 3332.920 1821.975 3332.965 ;
        RECT 1822.130 3332.920 1822.450 3332.980 ;
        RECT 1821.685 3332.780 1822.450 3332.920 ;
        RECT 1821.685 3332.735 1821.975 3332.780 ;
        RECT 1822.130 3332.720 1822.450 3332.780 ;
        RECT 1821.670 3270.700 1821.990 3270.760 ;
        RECT 1822.590 3270.700 1822.910 3270.760 ;
        RECT 1821.670 3270.560 1822.910 3270.700 ;
        RECT 1821.670 3270.500 1821.990 3270.560 ;
        RECT 1822.590 3270.500 1822.910 3270.560 ;
        RECT 1821.670 3174.140 1821.990 3174.200 ;
        RECT 1822.590 3174.140 1822.910 3174.200 ;
        RECT 1821.670 3174.000 1822.910 3174.140 ;
        RECT 1821.670 3173.940 1821.990 3174.000 ;
        RECT 1822.590 3173.940 1822.910 3174.000 ;
        RECT 1821.670 3077.580 1821.990 3077.640 ;
        RECT 1822.590 3077.580 1822.910 3077.640 ;
        RECT 1821.670 3077.440 1822.910 3077.580 ;
        RECT 1821.670 3077.380 1821.990 3077.440 ;
        RECT 1822.590 3077.380 1822.910 3077.440 ;
        RECT 1821.670 2981.020 1821.990 2981.080 ;
        RECT 1822.590 2981.020 1822.910 2981.080 ;
        RECT 1821.670 2980.880 1822.910 2981.020 ;
        RECT 1821.670 2980.820 1821.990 2980.880 ;
        RECT 1822.590 2980.820 1822.910 2980.880 ;
        RECT 1820.750 2946.340 1821.070 2946.400 ;
        RECT 1822.130 2946.340 1822.450 2946.400 ;
        RECT 1820.750 2946.200 1822.450 2946.340 ;
        RECT 1820.750 2946.140 1821.070 2946.200 ;
        RECT 1822.130 2946.140 1822.450 2946.200 ;
        RECT 1822.130 2849.440 1822.450 2849.500 ;
        RECT 1821.935 2849.300 1822.450 2849.440 ;
        RECT 1822.130 2849.240 1822.450 2849.300 ;
        RECT 1822.145 2815.440 1822.435 2815.485 ;
        RECT 1823.050 2815.440 1823.370 2815.500 ;
        RECT 1822.145 2815.300 1823.370 2815.440 ;
        RECT 1822.145 2815.255 1822.435 2815.300 ;
        RECT 1823.050 2815.240 1823.370 2815.300 ;
        RECT 1822.130 2753.220 1822.450 2753.280 ;
        RECT 1823.510 2753.220 1823.830 2753.280 ;
        RECT 1822.130 2753.080 1823.830 2753.220 ;
        RECT 1822.130 2753.020 1822.450 2753.080 ;
        RECT 1823.510 2753.020 1823.830 2753.080 ;
        RECT 1823.510 2719.220 1823.830 2719.280 ;
        RECT 1823.140 2719.080 1823.830 2719.220 ;
        RECT 1823.140 2718.600 1823.280 2719.080 ;
        RECT 1823.510 2719.020 1823.830 2719.080 ;
        RECT 1823.050 2718.340 1823.370 2718.600 ;
        RECT 1822.130 2656.660 1822.450 2656.720 ;
        RECT 1823.510 2656.660 1823.830 2656.720 ;
        RECT 1822.130 2656.520 1823.830 2656.660 ;
        RECT 1822.130 2656.460 1822.450 2656.520 ;
        RECT 1823.510 2656.460 1823.830 2656.520 ;
        RECT 1822.590 2608.380 1822.910 2608.440 ;
        RECT 1823.510 2608.380 1823.830 2608.440 ;
        RECT 1822.590 2608.240 1823.830 2608.380 ;
        RECT 1822.590 2608.180 1822.910 2608.240 ;
        RECT 1823.510 2608.180 1823.830 2608.240 ;
        RECT 1821.670 2560.100 1821.990 2560.160 ;
        RECT 1822.130 2560.100 1822.450 2560.160 ;
        RECT 1821.670 2559.960 1822.450 2560.100 ;
        RECT 1821.670 2559.900 1821.990 2559.960 ;
        RECT 1822.130 2559.900 1822.450 2559.960 ;
        RECT 1821.670 2517.940 1821.990 2518.000 ;
        RECT 1535.180 2517.800 1821.990 2517.940 ;
        RECT 1501.510 2517.600 1501.830 2517.660 ;
        RECT 1535.180 2517.600 1535.320 2517.800 ;
        RECT 1821.670 2517.740 1821.990 2517.800 ;
        RECT 1501.510 2517.460 1535.320 2517.600 ;
        RECT 1501.510 2517.400 1501.830 2517.460 ;
      LAYER via ;
        RECT 1821.700 3380.660 1821.960 3380.920 ;
        RECT 1822.160 3332.720 1822.420 3332.980 ;
        RECT 1821.700 3270.500 1821.960 3270.760 ;
        RECT 1822.620 3270.500 1822.880 3270.760 ;
        RECT 1821.700 3173.940 1821.960 3174.200 ;
        RECT 1822.620 3173.940 1822.880 3174.200 ;
        RECT 1821.700 3077.380 1821.960 3077.640 ;
        RECT 1822.620 3077.380 1822.880 3077.640 ;
        RECT 1821.700 2980.820 1821.960 2981.080 ;
        RECT 1822.620 2980.820 1822.880 2981.080 ;
        RECT 1820.780 2946.140 1821.040 2946.400 ;
        RECT 1822.160 2946.140 1822.420 2946.400 ;
        RECT 1822.160 2849.240 1822.420 2849.500 ;
        RECT 1823.080 2815.240 1823.340 2815.500 ;
        RECT 1822.160 2753.020 1822.420 2753.280 ;
        RECT 1823.540 2753.020 1823.800 2753.280 ;
        RECT 1823.540 2719.020 1823.800 2719.280 ;
        RECT 1823.080 2718.340 1823.340 2718.600 ;
        RECT 1822.160 2656.460 1822.420 2656.720 ;
        RECT 1823.540 2656.460 1823.800 2656.720 ;
        RECT 1822.620 2608.180 1822.880 2608.440 ;
        RECT 1823.540 2608.180 1823.800 2608.440 ;
        RECT 1821.700 2559.900 1821.960 2560.160 ;
        RECT 1822.160 2559.900 1822.420 2560.160 ;
        RECT 1501.540 2517.400 1501.800 2517.660 ;
        RECT 1821.700 2517.740 1821.960 2518.000 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1824.770 3519.700 1825.330 3524.800 ;
=======
        RECT 1824.770 3517.600 1825.330 3524.800 ;
<<<<<<< HEAD
        RECT 1824.980 3499.950 1825.120 3517.600 ;
        RECT 1510.740 3499.630 1511.000 3499.950 ;
        RECT 1824.920 3499.630 1825.180 3499.950 ;
        RECT 1510.270 2499.410 1510.550 2500.000 ;
        RECT 1510.800 2499.410 1510.940 3499.630 ;
        RECT 1510.270 2499.270 1510.940 2499.410 ;
        RECT 1510.270 2496.000 1510.550 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3430.445 1825.580 3517.230 ;
        RECT 1825.370 3430.075 1825.650 3430.445 ;
        RECT 1822.610 3429.395 1822.890 3429.765 ;
        RECT 1822.680 3394.970 1822.820 3429.395 ;
        RECT 1821.760 3394.830 1822.820 3394.970 ;
        RECT 1821.760 3380.950 1821.900 3394.830 ;
        RECT 1821.700 3380.630 1821.960 3380.950 ;
        RECT 1822.160 3332.690 1822.420 3333.010 ;
        RECT 1822.220 3298.410 1822.360 3332.690 ;
        RECT 1822.220 3298.270 1822.820 3298.410 ;
        RECT 1822.680 3270.790 1822.820 3298.270 ;
        RECT 1821.700 3270.470 1821.960 3270.790 ;
        RECT 1822.620 3270.470 1822.880 3270.790 ;
        RECT 1821.760 3222.250 1821.900 3270.470 ;
        RECT 1821.760 3222.110 1822.820 3222.250 ;
        RECT 1822.680 3174.230 1822.820 3222.110 ;
        RECT 1821.700 3173.910 1821.960 3174.230 ;
        RECT 1822.620 3173.910 1822.880 3174.230 ;
        RECT 1821.760 3125.690 1821.900 3173.910 ;
        RECT 1821.760 3125.550 1822.820 3125.690 ;
        RECT 1822.680 3077.670 1822.820 3125.550 ;
        RECT 1821.700 3077.350 1821.960 3077.670 ;
        RECT 1822.620 3077.350 1822.880 3077.670 ;
        RECT 1821.760 3029.130 1821.900 3077.350 ;
        RECT 1821.760 3028.990 1822.820 3029.130 ;
        RECT 1822.680 2981.110 1822.820 3028.990 ;
        RECT 1821.700 2980.850 1821.960 2981.110 ;
        RECT 1821.700 2980.790 1822.360 2980.850 ;
        RECT 1822.620 2980.790 1822.880 2981.110 ;
        RECT 1821.760 2980.710 1822.360 2980.790 ;
        RECT 1822.220 2980.170 1822.360 2980.710 ;
        RECT 1822.220 2980.030 1822.820 2980.170 ;
        RECT 1822.680 2959.770 1822.820 2980.030 ;
        RECT 1822.220 2959.630 1822.820 2959.770 ;
        RECT 1822.220 2946.430 1822.360 2959.630 ;
        RECT 1820.780 2946.110 1821.040 2946.430 ;
        RECT 1822.160 2946.110 1822.420 2946.430 ;
        RECT 1820.840 2898.685 1820.980 2946.110 ;
        RECT 1820.770 2898.315 1821.050 2898.685 ;
        RECT 1821.690 2898.315 1821.970 2898.685 ;
        RECT 1821.760 2863.210 1821.900 2898.315 ;
        RECT 1821.760 2863.070 1822.360 2863.210 ;
        RECT 1822.220 2849.530 1822.360 2863.070 ;
        RECT 1822.160 2849.210 1822.420 2849.530 ;
        RECT 1823.080 2815.210 1823.340 2815.530 ;
        RECT 1823.140 2801.445 1823.280 2815.210 ;
        RECT 1822.150 2801.075 1822.430 2801.445 ;
        RECT 1823.070 2801.075 1823.350 2801.445 ;
        RECT 1822.220 2753.310 1822.360 2801.075 ;
        RECT 1822.160 2752.990 1822.420 2753.310 ;
        RECT 1823.540 2752.990 1823.800 2753.310 ;
        RECT 1823.600 2719.310 1823.740 2752.990 ;
        RECT 1823.540 2718.990 1823.800 2719.310 ;
        RECT 1823.080 2718.310 1823.340 2718.630 ;
        RECT 1823.140 2704.885 1823.280 2718.310 ;
        RECT 1822.150 2704.515 1822.430 2704.885 ;
        RECT 1823.070 2704.515 1823.350 2704.885 ;
        RECT 1822.220 2656.750 1822.360 2704.515 ;
        RECT 1822.160 2656.430 1822.420 2656.750 ;
        RECT 1823.540 2656.430 1823.800 2656.750 ;
        RECT 1823.600 2608.470 1823.740 2656.430 ;
        RECT 1822.620 2608.325 1822.880 2608.470 ;
        RECT 1821.690 2607.955 1821.970 2608.325 ;
        RECT 1822.610 2607.955 1822.890 2608.325 ;
        RECT 1823.540 2608.150 1823.800 2608.470 ;
        RECT 1821.760 2560.190 1821.900 2607.955 ;
        RECT 1821.700 2559.870 1821.960 2560.190 ;
        RECT 1822.160 2559.870 1822.420 2560.190 ;
        RECT 1822.220 2525.930 1822.360 2559.870 ;
        RECT 1821.760 2525.790 1822.360 2525.930 ;
        RECT 1821.760 2518.030 1821.900 2525.790 ;
        RECT 1821.700 2517.710 1821.960 2518.030 ;
        RECT 1501.540 2517.370 1501.800 2517.690 ;
        RECT 1501.600 2500.000 1501.740 2517.370 ;
        RECT 1501.530 2496.000 1501.810 2500.000 ;
      LAYER via2 ;
        RECT 1825.370 3430.120 1825.650 3430.400 ;
        RECT 1822.610 3429.440 1822.890 3429.720 ;
        RECT 1820.770 2898.360 1821.050 2898.640 ;
        RECT 1821.690 2898.360 1821.970 2898.640 ;
        RECT 1822.150 2801.120 1822.430 2801.400 ;
        RECT 1823.070 2801.120 1823.350 2801.400 ;
        RECT 1822.150 2704.560 1822.430 2704.840 ;
        RECT 1823.070 2704.560 1823.350 2704.840 ;
        RECT 1821.690 2608.000 1821.970 2608.280 ;
        RECT 1822.610 2608.000 1822.890 2608.280 ;
      LAYER met3 ;
        RECT 1825.345 3430.410 1825.675 3430.425 ;
        RECT 1821.910 3430.110 1825.675 3430.410 ;
        RECT 1821.910 3429.730 1822.210 3430.110 ;
        RECT 1825.345 3430.095 1825.675 3430.110 ;
        RECT 1822.585 3429.730 1822.915 3429.745 ;
        RECT 1821.910 3429.430 1822.915 3429.730 ;
        RECT 1822.585 3429.415 1822.915 3429.430 ;
        RECT 1820.745 2898.650 1821.075 2898.665 ;
        RECT 1821.665 2898.650 1821.995 2898.665 ;
        RECT 1820.745 2898.350 1821.995 2898.650 ;
        RECT 1820.745 2898.335 1821.075 2898.350 ;
        RECT 1821.665 2898.335 1821.995 2898.350 ;
        RECT 1822.125 2801.410 1822.455 2801.425 ;
        RECT 1823.045 2801.410 1823.375 2801.425 ;
        RECT 1822.125 2801.110 1823.375 2801.410 ;
        RECT 1822.125 2801.095 1822.455 2801.110 ;
        RECT 1823.045 2801.095 1823.375 2801.110 ;
        RECT 1822.125 2704.850 1822.455 2704.865 ;
        RECT 1823.045 2704.850 1823.375 2704.865 ;
        RECT 1822.125 2704.550 1823.375 2704.850 ;
        RECT 1822.125 2704.535 1822.455 2704.550 ;
        RECT 1823.045 2704.535 1823.375 2704.550 ;
        RECT 1821.665 2608.290 1821.995 2608.305 ;
        RECT 1822.585 2608.290 1822.915 2608.305 ;
        RECT 1821.665 2607.990 1822.915 2608.290 ;
        RECT 1821.665 2607.975 1821.995 2607.990 ;
        RECT 1822.585 2607.975 1822.915 2607.990 ;
>>>>>>> re-updated local openlane
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3504.620 1500.910 3504.680 ;
        RECT 1503.810 3504.620 1504.130 3504.680 ;
        RECT 1500.590 3504.480 1504.130 3504.620 ;
        RECT 1500.590 3504.420 1500.910 3504.480 ;
        RECT 1503.810 3504.420 1504.130 3504.480 ;
        RECT 1503.810 2517.940 1504.130 2518.000 ;
        RECT 1520.830 2517.940 1521.150 2518.000 ;
        RECT 1503.810 2517.800 1521.150 2517.940 ;
        RECT 1503.810 2517.740 1504.130 2517.800 ;
        RECT 1520.830 2517.740 1521.150 2517.800 ;
      LAYER via ;
        RECT 1500.620 3504.420 1500.880 3504.680 ;
        RECT 1503.840 3504.420 1504.100 3504.680 ;
        RECT 1503.840 2517.740 1504.100 2518.000 ;
        RECT 1520.860 2517.740 1521.120 2518.000 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1500.470 3519.700 1501.030 3524.800 ;
=======
        RECT 1500.470 3517.600 1501.030 3524.800 ;
<<<<<<< HEAD
        RECT 1500.680 3499.270 1500.820 3517.600 ;
        RECT 1500.620 3498.950 1500.880 3499.270 ;
        RECT 1525.000 3498.950 1525.260 3499.270 ;
        RECT 1525.060 2498.730 1525.200 3498.950 ;
        RECT 1530.050 2498.730 1530.330 2500.000 ;
        RECT 1525.060 2498.590 1530.330 2498.730 ;
        RECT 1530.050 2496.000 1530.330 2498.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1500.680 3504.710 1500.820 3517.600 ;
        RECT 1500.620 3504.390 1500.880 3504.710 ;
        RECT 1503.840 3504.390 1504.100 3504.710 ;
        RECT 1503.900 2518.030 1504.040 3504.390 ;
        RECT 1503.840 2517.710 1504.100 2518.030 ;
        RECT 1520.860 2517.710 1521.120 2518.030 ;
        RECT 1520.920 2500.000 1521.060 2517.710 ;
        RECT 1520.850 2496.000 1521.130 2500.000 ;
>>>>>>> re-updated local openlane
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1172.610 2507.400 1172.930 2507.460 ;
        RECT 1955.990 2507.400 1956.310 2507.460 ;
        RECT 1172.610 2507.260 1956.310 2507.400 ;
        RECT 1172.610 2507.200 1172.930 2507.260 ;
        RECT 1955.990 2507.200 1956.310 2507.260 ;
        RECT 1955.990 324.260 1956.310 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 1955.990 324.120 2899.310 324.260 ;
        RECT 1955.990 324.060 1956.310 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 1172.640 2507.200 1172.900 2507.460 ;
        RECT 1956.020 2507.200 1956.280 2507.460 ;
        RECT 1956.020 324.060 1956.280 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 1172.640 2507.170 1172.900 2507.490 ;
        RECT 1956.020 2507.170 1956.280 2507.490 ;
        RECT 1172.700 2500.000 1172.840 2507.170 ;
        RECT 1172.630 2496.000 1172.910 2500.000 ;
        RECT 1956.080 324.350 1956.220 2507.170 ;
        RECT 1956.020 324.030 1956.280 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 322.060 2924.800 323.260 ;
=======
        RECT 1174.445 2498.810 1174.775 2498.825 ;
        RECT 1178.790 2498.810 1179.170 2498.820 ;
        RECT 1174.445 2498.510 1179.170 2498.810 ;
        RECT 1174.445 2498.495 1174.775 2498.510 ;
        RECT 1178.790 2498.500 1179.170 2498.510 ;
=======
        RECT 2898.985 322.810 2899.315 322.825 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
<<<<<<< HEAD
        RECT 2835.750 318.430 2883.890 318.730 ;
        RECT 2786.990 317.750 2788.210 318.050 ;
        RECT 2883.590 318.050 2883.890 318.430 ;
        RECT 2884.510 318.430 2917.010 318.730 ;
        RECT 2884.510 318.050 2884.810 318.430 ;
        RECT 2883.590 317.750 2884.810 318.050 ;
        RECT 2052.585 317.735 2052.915 317.750 ;
        RECT 1895.265 316.390 1931.690 316.690 ;
        RECT 1895.265 316.375 1895.595 316.390 ;
      LAYER via3 ;
        RECT 1178.820 2498.500 1179.140 2498.820 ;
        RECT 1178.820 319.100 1179.140 319.420 ;
        RECT 1248.740 319.100 1249.060 319.420 ;
        RECT 1248.740 317.740 1249.060 318.060 ;
        RECT 1980.140 320.460 1980.460 320.780 ;
        RECT 1980.140 319.100 1980.460 319.420 ;
      LAYER met4 ;
        RECT 1178.815 2498.495 1179.145 2498.825 ;
        RECT 1178.830 319.425 1179.130 2498.495 ;
        RECT 1980.135 320.455 1980.465 320.785 ;
        RECT 1980.150 319.425 1980.450 320.455 ;
        RECT 1178.815 319.095 1179.145 319.425 ;
        RECT 1248.735 319.095 1249.065 319.425 ;
        RECT 1980.135 319.095 1980.465 319.425 ;
        RECT 1248.750 318.065 1249.050 319.095 ;
        RECT 1248.735 317.735 1249.065 318.065 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1249.045 2517.445 1249.215 2518.295 ;
        RECT 1345.645 2517.785 1345.815 2518.635 ;
        RECT 1393.485 2517.445 1393.655 2518.635 ;
        RECT 1400.845 2517.445 1401.015 2518.295 ;
        RECT 1462.485 2517.785 1462.655 2519.315 ;
        RECT 1496.985 2518.125 1497.155 2519.315 ;
      LAYER mcon ;
        RECT 1462.485 2519.145 1462.655 2519.315 ;
        RECT 1345.645 2518.465 1345.815 2518.635 ;
        RECT 1249.045 2518.125 1249.215 2518.295 ;
        RECT 1393.485 2518.465 1393.655 2518.635 ;
        RECT 1400.845 2518.125 1401.015 2518.295 ;
        RECT 1496.985 2519.145 1497.155 2519.315 ;
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1462.425 2519.300 1462.715 2519.345 ;
        RECT 1496.925 2519.300 1497.215 2519.345 ;
        RECT 1462.425 2519.160 1497.215 2519.300 ;
        RECT 1462.425 2519.115 1462.715 2519.160 ;
        RECT 1496.925 2519.115 1497.215 2519.160 ;
        RECT 1345.585 2518.620 1345.875 2518.665 ;
        RECT 1393.425 2518.620 1393.715 2518.665 ;
        RECT 1345.585 2518.480 1393.715 2518.620 ;
        RECT 1345.585 2518.435 1345.875 2518.480 ;
        RECT 1393.425 2518.435 1393.715 2518.480 ;
        RECT 1248.985 2518.280 1249.275 2518.325 ;
        RECT 1220.540 2518.140 1249.275 2518.280 ;
        RECT 1179.510 2517.600 1179.830 2517.660 ;
        RECT 1220.540 2517.600 1220.680 2518.140 ;
        RECT 1248.985 2518.095 1249.275 2518.140 ;
        RECT 1400.785 2518.280 1401.075 2518.325 ;
        RECT 1496.925 2518.280 1497.215 2518.325 ;
        RECT 1540.150 2518.280 1540.470 2518.340 ;
        RECT 1400.785 2518.140 1415.260 2518.280 ;
        RECT 1400.785 2518.095 1401.075 2518.140 ;
        RECT 1345.585 2517.940 1345.875 2517.985 ;
        RECT 1270.220 2517.800 1345.875 2517.940 ;
        RECT 1415.120 2517.940 1415.260 2518.140 ;
        RECT 1496.925 2518.140 1540.470 2518.280 ;
        RECT 1496.925 2518.095 1497.215 2518.140 ;
        RECT 1540.150 2518.080 1540.470 2518.140 ;
        RECT 1462.425 2517.940 1462.715 2517.985 ;
        RECT 1415.120 2517.800 1462.715 2517.940 ;
        RECT 1179.510 2517.460 1220.680 2517.600 ;
        RECT 1248.985 2517.600 1249.275 2517.645 ;
        RECT 1270.220 2517.600 1270.360 2517.800 ;
        RECT 1345.585 2517.755 1345.875 2517.800 ;
        RECT 1462.425 2517.755 1462.715 2517.800 ;
        RECT 1248.985 2517.460 1270.360 2517.600 ;
        RECT 1393.425 2517.600 1393.715 2517.645 ;
        RECT 1400.785 2517.600 1401.075 2517.645 ;
        RECT 1393.425 2517.460 1401.075 2517.600 ;
        RECT 1179.510 2517.400 1179.830 2517.460 ;
        RECT 1248.985 2517.415 1249.275 2517.460 ;
        RECT 1393.425 2517.415 1393.715 2517.460 ;
        RECT 1400.785 2517.415 1401.075 2517.460 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 2517.400 1179.800 2517.660 ;
        RECT 1540.180 2518.080 1540.440 2518.340 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1175.710 3519.700 1176.270 3524.800 ;
=======
        RECT 1175.710 3517.600 1176.270 3524.800 ;
<<<<<<< HEAD
        RECT 1175.920 3500.290 1176.060 3517.600 ;
        RECT 1175.860 3499.970 1176.120 3500.290 ;
        RECT 1545.700 3499.970 1545.960 3500.290 ;
        RECT 1545.760 2498.730 1545.900 3499.970 ;
        RECT 1549.830 2498.730 1550.110 2500.000 ;
        RECT 1545.760 2498.590 1550.110 2498.730 ;
        RECT 1549.830 2496.000 1550.110 2498.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 2517.690 1179.740 3498.270 ;
        RECT 1540.180 2518.050 1540.440 2518.370 ;
        RECT 1179.540 2517.370 1179.800 2517.690 ;
        RECT 1540.240 2500.000 1540.380 2518.050 ;
        RECT 1540.170 2496.000 1540.450 2500.000 ;
>>>>>>> re-updated local openlane
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 1559.930 3501.220 1560.250 3501.280 ;
        RECT 851.530 3501.080 1560.250 3501.220 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
        RECT 1559.930 3501.020 1560.250 3501.080 ;
      LAYER via ;
        RECT 851.560 3501.020 851.820 3501.280 ;
        RECT 1559.960 3501.020 1560.220 3501.280 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 851.410 3519.700 851.970 3524.800 ;
=======
        RECT 851.410 3517.600 851.970 3524.800 ;
<<<<<<< HEAD
        RECT 851.620 3505.050 851.760 3517.600 ;
        RECT 851.560 3504.730 851.820 3505.050 ;
        RECT 1566.400 3504.730 1566.660 3505.050 ;
        RECT 1566.460 2498.730 1566.600 3504.730 ;
        RECT 1569.610 2498.730 1569.890 2500.000 ;
        RECT 1566.460 2498.590 1569.890 2498.730 ;
        RECT 1569.610 2496.000 1569.890 2498.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 1559.960 3500.990 1560.220 3501.310 ;
        RECT 1559.490 2499.410 1559.770 2500.000 ;
        RECT 1560.020 2499.410 1560.160 3500.990 ;
        RECT 1559.490 2499.270 1560.160 2499.410 ;
        RECT 1559.490 2496.000 1559.770 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.230 3503.600 527.550 3503.660 ;
        RECT 1573.270 3503.600 1573.590 3503.660 ;
        RECT 527.230 3503.460 1573.590 3503.600 ;
        RECT 527.230 3503.400 527.550 3503.460 ;
        RECT 1573.270 3503.400 1573.590 3503.460 ;
      LAYER via ;
        RECT 527.260 3503.400 527.520 3503.660 ;
        RECT 1573.300 3503.400 1573.560 3503.660 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 527.110 3519.700 527.670 3524.800 ;
=======
        RECT 527.110 3517.600 527.670 3524.800 ;
<<<<<<< HEAD
        RECT 527.320 3503.350 527.460 3517.600 ;
        RECT 527.260 3503.030 527.520 3503.350 ;
        RECT 1587.100 3503.030 1587.360 3503.350 ;
        RECT 1587.160 2499.410 1587.300 3503.030 ;
        RECT 1589.390 2499.410 1589.670 2500.000 ;
        RECT 1587.160 2499.270 1589.670 2499.410 ;
        RECT 1589.390 2496.000 1589.670 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 527.320 3503.690 527.460 3517.600 ;
        RECT 527.260 3503.370 527.520 3503.690 ;
        RECT 1573.300 3503.370 1573.560 3503.690 ;
        RECT 1573.360 2500.770 1573.500 3503.370 ;
        RECT 1573.360 2500.630 1576.720 2500.770 ;
        RECT 1576.580 2499.410 1576.720 2500.630 ;
        RECT 1578.810 2499.410 1579.090 2500.000 ;
        RECT 1576.580 2499.270 1579.090 2499.410 ;
        RECT 1578.810 2496.000 1579.090 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 1593.970 3501.900 1594.290 3501.960 ;
        RECT 202.470 3501.760 1594.290 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 1593.970 3501.700 1594.290 3501.760 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 1594.000 3501.700 1594.260 3501.960 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 202.350 3519.700 202.910 3524.800 ;
=======
        RECT 202.350 3517.600 202.910 3524.800 ;
<<<<<<< HEAD
        RECT 202.560 3501.650 202.700 3517.600 ;
        RECT 202.500 3501.330 202.760 3501.650 ;
        RECT 1607.800 3501.330 1608.060 3501.650 ;
        RECT 1607.860 2499.410 1608.000 3501.330 ;
        RECT 1609.170 2499.410 1609.450 2500.000 ;
        RECT 1607.860 2499.270 1609.450 2499.410 ;
        RECT 1609.170 2496.000 1609.450 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 1594.000 3501.670 1594.260 3501.990 ;
        RECT 1594.060 2499.410 1594.200 3501.670 ;
        RECT 1598.130 2499.410 1598.410 2500.000 ;
        RECT 1594.060 2499.270 1598.410 2499.410 ;
        RECT 1598.130 2496.000 1598.410 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 1614.670 3408.740 1614.990 3408.800 ;
        RECT 17.550 3408.600 1614.990 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 1614.670 3408.540 1614.990 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 1614.700 3408.540 1614.960 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 1614.700 3408.510 1614.960 3408.830 ;
        RECT 1614.760 2498.730 1614.900 3408.510 ;
        RECT 1617.450 2498.730 1617.730 2500.000 ;
        RECT 1614.760 2498.590 1617.730 2498.730 ;
        RECT 1617.450 2496.000 1617.730 2498.590 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3410.620 0.300 3411.820 ;
=======
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 3119.060 16.490 3119.120 ;
        RECT 1635.370 3119.060 1635.690 3119.120 ;
        RECT 16.170 3118.920 1635.690 3119.060 ;
        RECT 16.170 3118.860 16.490 3118.920 ;
        RECT 1635.370 3118.860 1635.690 3118.920 ;
      LAYER via ;
        RECT 16.200 3118.860 16.460 3119.120 ;
        RECT 1635.400 3118.860 1635.660 3119.120 ;
      LAYER met2 ;
        RECT 16.190 3124.075 16.470 3124.445 ;
        RECT 16.260 3119.150 16.400 3124.075 ;
        RECT 16.200 3118.830 16.460 3119.150 ;
        RECT 1635.400 3118.830 1635.660 3119.150 ;
        RECT 1635.460 2499.410 1635.600 3118.830 ;
        RECT 1636.770 2499.410 1637.050 2500.000 ;
        RECT 1635.460 2499.270 1637.050 2499.410 ;
        RECT 1636.770 2496.000 1637.050 2499.270 ;
      LAYER via2 ;
        RECT 16.190 3124.120 16.470 3124.400 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3123.660 0.300 3124.860 ;
=======
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 16.165 3124.410 16.495 3124.425 ;
        RECT -4.800 3124.110 16.495 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
<<<<<<< HEAD
        RECT 17.085 3124.095 17.415 3124.110 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.165 3124.095 16.495 3124.110 ;
>>>>>>> re-updated local openlane
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2836.180 16.950 2836.240 ;
        RECT 1656.070 2836.180 1656.390 2836.240 ;
        RECT 16.630 2836.040 1656.390 2836.180 ;
        RECT 16.630 2835.980 16.950 2836.040 ;
        RECT 1656.070 2835.980 1656.390 2836.040 ;
      LAYER via ;
        RECT 16.660 2835.980 16.920 2836.240 ;
        RECT 1656.100 2835.980 1656.360 2836.240 ;
      LAYER met2 ;
        RECT 16.650 2836.435 16.930 2836.805 ;
        RECT 16.720 2836.270 16.860 2836.435 ;
        RECT 16.660 2835.950 16.920 2836.270 ;
        RECT 1656.100 2835.950 1656.360 2836.270 ;
        RECT 1656.160 2500.000 1656.300 2835.950 ;
        RECT 1656.090 2496.000 1656.370 2500.000 ;
      LAYER via2 ;
        RECT 16.650 2836.480 16.930 2836.760 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2836.020 0.300 2837.220 ;
=======
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 16.625 2836.770 16.955 2836.785 ;
        RECT -4.800 2836.470 16.955 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
<<<<<<< HEAD
        RECT 17.085 2836.455 17.415 2836.470 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 2836.455 16.955 2836.470 ;
>>>>>>> re-updated local openlane
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2546.500 16.030 2546.560 ;
        RECT 1669.870 2546.500 1670.190 2546.560 ;
        RECT 15.710 2546.360 1670.190 2546.500 ;
        RECT 15.710 2546.300 16.030 2546.360 ;
        RECT 1669.870 2546.300 1670.190 2546.360 ;
      LAYER via ;
        RECT 15.740 2546.300 16.000 2546.560 ;
        RECT 1669.900 2546.300 1670.160 2546.560 ;
      LAYER met2 ;
        RECT 15.730 2549.475 16.010 2549.845 ;
        RECT 15.800 2546.590 15.940 2549.475 ;
        RECT 15.740 2546.270 16.000 2546.590 ;
        RECT 1669.900 2546.270 1670.160 2546.590 ;
        RECT 1669.960 2500.090 1670.100 2546.270 ;
        RECT 1669.960 2499.950 1673.780 2500.090 ;
        RECT 1673.640 2499.410 1673.780 2499.950 ;
        RECT 1675.410 2499.410 1675.690 2500.000 ;
        RECT 1673.640 2499.270 1675.690 2499.410 ;
        RECT 1675.410 2496.000 1675.690 2499.270 ;
      LAYER via2 ;
        RECT 15.730 2549.520 16.010 2549.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2549.060 0.300 2550.260 ;
=======
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 15.705 2549.810 16.035 2549.825 ;
        RECT -4.800 2549.510 16.035 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 15.705 2549.495 16.035 2549.510 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 879.590 2498.220 879.910 2498.280 ;
        RECT 1693.790 2498.220 1694.110 2498.280 ;
        RECT 879.590 2498.080 1694.110 2498.220 ;
        RECT 879.590 2498.020 879.910 2498.080 ;
        RECT 1693.790 2498.020 1694.110 2498.080 ;
        RECT 15.710 2262.940 16.030 2263.000 ;
        RECT 879.590 2262.940 879.910 2263.000 ;
        RECT 15.710 2262.800 879.910 2262.940 ;
        RECT 15.710 2262.740 16.030 2262.800 ;
        RECT 879.590 2262.740 879.910 2262.800 ;
      LAYER via ;
        RECT 879.620 2498.020 879.880 2498.280 ;
        RECT 1693.820 2498.020 1694.080 2498.280 ;
        RECT 15.740 2262.740 16.000 2263.000 ;
        RECT 879.620 2262.740 879.880 2263.000 ;
      LAYER met2 ;
        RECT 879.620 2497.990 879.880 2498.310 ;
        RECT 1693.820 2498.050 1694.080 2498.310 ;
        RECT 1695.190 2498.050 1695.470 2500.000 ;
        RECT 1693.820 2497.990 1695.470 2498.050 ;
        RECT 879.680 2263.030 879.820 2497.990 ;
        RECT 1693.880 2497.910 1695.470 2497.990 ;
        RECT 1695.190 2496.000 1695.470 2497.910 ;
        RECT 15.740 2262.710 16.000 2263.030 ;
        RECT 879.620 2262.710 879.880 2263.030 ;
        RECT 15.800 2262.205 15.940 2262.710 ;
        RECT 15.730 2261.835 16.010 2262.205 ;
      LAYER via2 ;
        RECT 15.730 2261.880 16.010 2262.160 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT -4.800 2261.420 0.300 2262.620 ;
=======
        RECT 1272.630 2514.450 1273.010 2514.460 ;
        RECT 1708.505 2514.450 1708.835 2514.465 ;
        RECT 1272.630 2514.150 1708.835 2514.450 ;
        RECT 1272.630 2514.140 1273.010 2514.150 ;
        RECT 1708.505 2514.135 1708.835 2514.150 ;
=======
>>>>>>> re-updated local openlane
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 15.705 2262.170 16.035 2262.185 ;
        RECT -4.800 2261.870 16.035 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
<<<<<<< HEAD
        RECT 19.590 2261.860 19.970 2261.870 ;
      LAYER via3 ;
        RECT 1272.660 2514.140 1272.980 2514.460 ;
        RECT 19.620 2261.860 19.940 2262.180 ;
      LAYER met4 ;
        RECT 1272.655 2514.135 1272.985 2514.465 ;
        RECT 1272.670 2273.490 1272.970 2514.135 ;
        RECT 1272.230 2272.310 1273.410 2273.490 ;
        RECT 19.190 2265.510 20.370 2266.690 ;
        RECT 19.630 2262.185 19.930 2265.510 ;
        RECT 19.615 2261.855 19.945 2262.185 ;
      LAYER met5 ;
        RECT 82.460 2272.100 130.980 2273.700 ;
        RECT 82.460 2266.900 84.060 2272.100 ;
        RECT 18.980 2265.300 84.060 2266.900 ;
        RECT 129.380 2266.900 130.980 2272.100 ;
        RECT 179.060 2272.100 227.580 2273.700 ;
        RECT 179.060 2266.900 180.660 2272.100 ;
        RECT 129.380 2265.300 180.660 2266.900 ;
        RECT 225.980 2266.900 227.580 2272.100 ;
        RECT 275.660 2272.100 324.180 2273.700 ;
        RECT 275.660 2266.900 277.260 2272.100 ;
        RECT 225.980 2265.300 277.260 2266.900 ;
        RECT 322.580 2266.900 324.180 2272.100 ;
        RECT 372.260 2272.100 420.780 2273.700 ;
        RECT 372.260 2266.900 373.860 2272.100 ;
        RECT 322.580 2265.300 373.860 2266.900 ;
        RECT 419.180 2266.900 420.780 2272.100 ;
        RECT 468.860 2272.100 517.380 2273.700 ;
        RECT 468.860 2266.900 470.460 2272.100 ;
        RECT 419.180 2265.300 470.460 2266.900 ;
        RECT 515.780 2266.900 517.380 2272.100 ;
        RECT 565.460 2272.100 613.980 2273.700 ;
        RECT 565.460 2266.900 567.060 2272.100 ;
        RECT 515.780 2265.300 567.060 2266.900 ;
        RECT 612.380 2266.900 613.980 2272.100 ;
        RECT 662.060 2272.100 710.580 2273.700 ;
        RECT 662.060 2266.900 663.660 2272.100 ;
        RECT 612.380 2265.300 663.660 2266.900 ;
        RECT 708.980 2266.900 710.580 2272.100 ;
        RECT 758.660 2272.100 807.180 2273.700 ;
        RECT 758.660 2266.900 760.260 2272.100 ;
        RECT 708.980 2265.300 760.260 2266.900 ;
        RECT 805.580 2266.900 807.180 2272.100 ;
        RECT 855.260 2272.100 903.780 2273.700 ;
        RECT 855.260 2266.900 856.860 2272.100 ;
        RECT 805.580 2265.300 856.860 2266.900 ;
        RECT 902.180 2266.900 903.780 2272.100 ;
        RECT 951.860 2272.100 1000.380 2273.700 ;
        RECT 951.860 2266.900 953.460 2272.100 ;
        RECT 902.180 2265.300 953.460 2266.900 ;
        RECT 998.780 2266.900 1000.380 2272.100 ;
        RECT 1048.460 2272.100 1096.980 2273.700 ;
        RECT 1048.460 2266.900 1050.060 2272.100 ;
        RECT 998.780 2265.300 1050.060 2266.900 ;
        RECT 1095.380 2266.900 1096.980 2272.100 ;
        RECT 1145.060 2272.100 1193.580 2273.700 ;
        RECT 1145.060 2266.900 1146.660 2272.100 ;
        RECT 1095.380 2265.300 1146.660 2266.900 ;
        RECT 1191.980 2266.900 1193.580 2272.100 ;
        RECT 1241.660 2272.100 1273.620 2273.700 ;
        RECT 1241.660 2266.900 1243.260 2272.100 ;
        RECT 1191.980 2265.300 1243.260 2266.900 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 15.705 2261.855 16.035 2261.870 ;
>>>>>>> re-updated local openlane
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 886.490 2506.380 886.810 2506.440 ;
        RECT 1714.490 2506.380 1714.810 2506.440 ;
        RECT 886.490 2506.240 1714.810 2506.380 ;
        RECT 886.490 2506.180 886.810 2506.240 ;
        RECT 1714.490 2506.180 1714.810 2506.240 ;
        RECT 14.790 1980.060 15.110 1980.120 ;
        RECT 886.490 1980.060 886.810 1980.120 ;
        RECT 14.790 1979.920 886.810 1980.060 ;
        RECT 14.790 1979.860 15.110 1979.920 ;
        RECT 886.490 1979.860 886.810 1979.920 ;
      LAYER via ;
        RECT 886.520 2506.180 886.780 2506.440 ;
        RECT 1714.520 2506.180 1714.780 2506.440 ;
        RECT 14.820 1979.860 15.080 1980.120 ;
        RECT 886.520 1979.860 886.780 1980.120 ;
      LAYER met2 ;
        RECT 886.520 2506.150 886.780 2506.470 ;
        RECT 1714.520 2506.150 1714.780 2506.470 ;
        RECT 886.580 1980.150 886.720 2506.150 ;
        RECT 1714.580 2500.000 1714.720 2506.150 ;
        RECT 1714.510 2496.000 1714.790 2500.000 ;
        RECT 14.820 1979.830 15.080 1980.150 ;
        RECT 886.520 1979.830 886.780 1980.150 ;
        RECT 14.880 1975.245 15.020 1979.830 ;
        RECT 14.810 1974.875 15.090 1975.245 ;
      LAYER via2 ;
        RECT 14.810 1974.920 15.090 1975.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1974.460 0.300 1975.660 ;
=======
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 14.785 1975.210 15.115 1975.225 ;
        RECT -4.800 1974.910 15.115 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 14.785 1974.895 15.115 1974.910 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1193.310 2499.580 1193.630 2499.640 ;
        RECT 1969.790 2499.580 1970.110 2499.640 ;
        RECT 1193.310 2499.440 1970.110 2499.580 ;
        RECT 1193.310 2499.380 1193.630 2499.440 ;
        RECT 1969.790 2499.380 1970.110 2499.440 ;
        RECT 1969.790 558.860 1970.110 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 1969.790 558.720 2899.310 558.860 ;
        RECT 1969.790 558.660 1970.110 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 1193.340 2499.380 1193.600 2499.640 ;
        RECT 1969.820 2499.380 1970.080 2499.640 ;
        RECT 1969.820 558.660 1970.080 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 1191.950 2499.410 1192.230 2500.000 ;
        RECT 1193.340 2499.410 1193.600 2499.670 ;
        RECT 1191.950 2499.350 1193.600 2499.410 ;
        RECT 1969.820 2499.350 1970.080 2499.670 ;
        RECT 1191.950 2499.270 1193.540 2499.350 ;
        RECT 1191.950 2496.000 1192.230 2499.270 ;
        RECT 1969.880 558.950 1970.020 2499.350 ;
        RECT 1969.820 558.630 1970.080 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 556.660 2924.800 557.860 ;
=======
        RECT 1190.750 2498.130 1191.130 2498.140 ;
        RECT 1191.465 2498.130 1191.795 2498.145 ;
        RECT 1190.750 2497.830 1191.795 2498.130 ;
        RECT 1190.750 2497.820 1191.130 2497.830 ;
        RECT 1191.465 2497.815 1191.795 2497.830 ;
=======
        RECT 2898.985 557.410 2899.315 557.425 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
<<<<<<< HEAD
        RECT 2835.750 553.030 2883.890 553.330 ;
        RECT 2786.990 552.350 2788.210 552.650 ;
        RECT 2883.590 552.650 2883.890 553.030 ;
        RECT 2884.510 553.030 2917.010 553.330 ;
        RECT 2884.510 552.650 2884.810 553.030 ;
        RECT 2883.590 552.350 2884.810 552.650 ;
        RECT 2052.585 552.335 2052.915 552.350 ;
        RECT 1895.265 550.990 1931.690 551.290 ;
        RECT 1895.265 550.975 1895.595 550.990 ;
      LAYER via3 ;
        RECT 1190.780 2497.820 1191.100 2498.140 ;
        RECT 1980.140 555.060 1980.460 555.380 ;
        RECT 1190.780 554.380 1191.100 554.700 ;
        RECT 1980.140 553.700 1980.460 554.020 ;
      LAYER met4 ;
        RECT 1190.775 2497.815 1191.105 2498.145 ;
        RECT 1190.790 554.705 1191.090 2497.815 ;
        RECT 1980.135 555.055 1980.465 555.385 ;
        RECT 1190.775 554.375 1191.105 554.705 ;
        RECT 1980.150 554.025 1980.450 555.055 ;
        RECT 1980.135 553.695 1980.465 554.025 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 72.750 2505.700 73.070 2505.760 ;
        RECT 1733.810 2505.700 1734.130 2505.760 ;
        RECT 72.750 2505.560 1734.130 2505.700 ;
        RECT 72.750 2505.500 73.070 2505.560 ;
        RECT 1733.810 2505.500 1734.130 2505.560 ;
        RECT 18.930 1690.040 19.250 1690.100 ;
        RECT 72.750 1690.040 73.070 1690.100 ;
        RECT 18.930 1689.900 73.070 1690.040 ;
        RECT 18.930 1689.840 19.250 1689.900 ;
        RECT 72.750 1689.840 73.070 1689.900 ;
      LAYER via ;
        RECT 72.780 2505.500 73.040 2505.760 ;
        RECT 1733.840 2505.500 1734.100 2505.760 ;
        RECT 18.960 1689.840 19.220 1690.100 ;
        RECT 72.780 1689.840 73.040 1690.100 ;
      LAYER met2 ;
        RECT 72.780 2505.470 73.040 2505.790 ;
        RECT 1733.840 2505.470 1734.100 2505.790 ;
        RECT 72.840 1690.130 72.980 2505.470 ;
        RECT 1733.900 2500.000 1734.040 2505.470 ;
        RECT 1733.830 2496.000 1734.110 2500.000 ;
        RECT 18.960 1689.810 19.220 1690.130 ;
        RECT 72.780 1689.810 73.040 1690.130 ;
        RECT 19.020 1687.605 19.160 1689.810 ;
        RECT 18.950 1687.235 19.230 1687.605 ;
      LAYER via2 ;
        RECT 18.950 1687.280 19.230 1687.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1686.820 0.300 1688.020 ;
=======
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 18.925 1687.570 19.255 1687.585 ;
        RECT -4.800 1687.270 19.255 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
<<<<<<< HEAD
        RECT 16.165 1687.255 16.495 1687.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 18.925 1687.255 19.255 1687.270 ;
>>>>>>> re-updated local openlane
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1128.450 2502.300 1128.770 2502.360 ;
        RECT 1753.130 2502.300 1753.450 2502.360 ;
        RECT 1128.450 2502.160 1753.450 2502.300 ;
        RECT 1128.450 2502.100 1128.770 2502.160 ;
        RECT 1753.130 2502.100 1753.450 2502.160 ;
        RECT 16.630 1476.520 16.950 1476.580 ;
        RECT 1128.450 1476.520 1128.770 1476.580 ;
        RECT 16.630 1476.380 1128.770 1476.520 ;
        RECT 16.630 1476.320 16.950 1476.380 ;
        RECT 1128.450 1476.320 1128.770 1476.380 ;
      LAYER via ;
        RECT 1128.480 2502.100 1128.740 2502.360 ;
        RECT 1753.160 2502.100 1753.420 2502.360 ;
        RECT 16.660 1476.320 16.920 1476.580 ;
        RECT 1128.480 1476.320 1128.740 1476.580 ;
      LAYER met2 ;
        RECT 1128.480 2502.070 1128.740 2502.390 ;
        RECT 1753.160 2502.070 1753.420 2502.390 ;
        RECT 1128.540 1476.610 1128.680 2502.070 ;
        RECT 1753.220 2500.000 1753.360 2502.070 ;
        RECT 1753.150 2496.000 1753.430 2500.000 ;
        RECT 16.660 1476.290 16.920 1476.610 ;
        RECT 1128.480 1476.290 1128.740 1476.610 ;
        RECT 16.720 1472.045 16.860 1476.290 ;
        RECT 16.650 1471.675 16.930 1472.045 ;
      LAYER via2 ;
        RECT 16.650 1471.720 16.930 1472.000 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1471.260 0.300 1472.460 ;
=======
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 16.625 1472.010 16.955 1472.025 ;
        RECT -4.800 1471.710 16.955 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
<<<<<<< HEAD
        RECT 20.305 1471.695 20.635 1471.710 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 1471.695 16.955 1471.710 ;
>>>>>>> re-updated local openlane
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1114.650 2509.440 1114.970 2509.500 ;
        RECT 1772.450 2509.440 1772.770 2509.500 ;
        RECT 1114.650 2509.300 1772.770 2509.440 ;
        RECT 1114.650 2509.240 1114.970 2509.300 ;
        RECT 1772.450 2509.240 1772.770 2509.300 ;
        RECT 15.710 1262.660 16.030 1262.720 ;
        RECT 1114.650 1262.660 1114.970 1262.720 ;
        RECT 15.710 1262.520 1114.970 1262.660 ;
        RECT 15.710 1262.460 16.030 1262.520 ;
        RECT 1114.650 1262.460 1114.970 1262.520 ;
      LAYER via ;
        RECT 1114.680 2509.240 1114.940 2509.500 ;
        RECT 1772.480 2509.240 1772.740 2509.500 ;
        RECT 15.740 1262.460 16.000 1262.720 ;
        RECT 1114.680 1262.460 1114.940 1262.720 ;
      LAYER met2 ;
        RECT 1114.680 2509.210 1114.940 2509.530 ;
        RECT 1772.480 2509.210 1772.740 2509.530 ;
        RECT 1114.740 1262.750 1114.880 2509.210 ;
        RECT 1772.540 2500.000 1772.680 2509.210 ;
        RECT 1772.470 2496.000 1772.750 2500.000 ;
        RECT 15.740 1262.430 16.000 1262.750 ;
        RECT 1114.680 1262.430 1114.940 1262.750 ;
        RECT 15.800 1256.485 15.940 1262.430 ;
        RECT 15.730 1256.115 16.010 1256.485 ;
      LAYER via2 ;
        RECT 15.730 1256.160 16.010 1256.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1255.700 0.300 1256.900 ;
=======
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 15.705 1256.450 16.035 1256.465 ;
        RECT -4.800 1256.150 16.035 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
<<<<<<< HEAD
        RECT 19.845 1256.135 20.175 1256.150 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 15.705 1256.135 16.035 1256.150 ;
>>>>>>> re-updated local openlane
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1093.950 2501.960 1094.270 2502.020 ;
        RECT 1791.770 2501.960 1792.090 2502.020 ;
        RECT 1093.950 2501.820 1792.090 2501.960 ;
        RECT 1093.950 2501.760 1094.270 2501.820 ;
        RECT 1791.770 2501.760 1792.090 2501.820 ;
        RECT 15.710 1041.660 16.030 1041.720 ;
        RECT 1093.950 1041.660 1094.270 1041.720 ;
        RECT 15.710 1041.520 1094.270 1041.660 ;
        RECT 15.710 1041.460 16.030 1041.520 ;
        RECT 1093.950 1041.460 1094.270 1041.520 ;
      LAYER via ;
        RECT 1093.980 2501.760 1094.240 2502.020 ;
        RECT 1791.800 2501.760 1792.060 2502.020 ;
        RECT 15.740 1041.460 16.000 1041.720 ;
        RECT 1093.980 1041.460 1094.240 1041.720 ;
      LAYER met2 ;
        RECT 1093.980 2501.730 1094.240 2502.050 ;
        RECT 1791.800 2501.730 1792.060 2502.050 ;
        RECT 1094.040 1041.750 1094.180 2501.730 ;
        RECT 1791.860 2500.000 1792.000 2501.730 ;
        RECT 1791.790 2496.000 1792.070 2500.000 ;
        RECT 15.740 1041.430 16.000 1041.750 ;
        RECT 1093.980 1041.430 1094.240 1041.750 ;
        RECT 15.800 1040.925 15.940 1041.430 ;
        RECT 15.730 1040.555 16.010 1040.925 ;
      LAYER via2 ;
        RECT 15.730 1040.600 16.010 1040.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1040.140 0.300 1041.340 ;
=======
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 15.705 1040.890 16.035 1040.905 ;
        RECT -4.800 1040.590 16.035 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
<<<<<<< HEAD
        RECT 19.385 1040.575 19.715 1040.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 15.705 1040.575 16.035 1040.590 ;
>>>>>>> re-updated local openlane
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1809.710 2496.320 1810.030 2496.580 ;
        RECT 1809.800 2495.500 1809.940 2496.320 ;
        RECT 1632.700 2495.360 1680.220 2495.500 ;
        RECT 1127.990 2495.160 1128.310 2495.220 ;
        RECT 1632.700 2495.160 1632.840 2495.360 ;
        RECT 1127.990 2495.020 1632.840 2495.160 ;
        RECT 1680.080 2495.160 1680.220 2495.360 ;
        RECT 1725.160 2495.360 1809.940 2495.500 ;
        RECT 1725.160 2495.160 1725.300 2495.360 ;
        RECT 1680.080 2495.020 1725.300 2495.160 ;
        RECT 1127.990 2494.960 1128.310 2495.020 ;
        RECT 14.790 827.800 15.110 827.860 ;
        RECT 1127.990 827.800 1128.310 827.860 ;
        RECT 14.790 827.660 1128.310 827.800 ;
        RECT 14.790 827.600 15.110 827.660 ;
        RECT 1127.990 827.600 1128.310 827.660 ;
      LAYER via ;
        RECT 1809.740 2496.320 1810.000 2496.580 ;
        RECT 1128.020 2494.960 1128.280 2495.220 ;
        RECT 14.820 827.600 15.080 827.860 ;
        RECT 1128.020 827.600 1128.280 827.860 ;
      LAYER met2 ;
        RECT 1811.110 2496.690 1811.390 2500.000 ;
        RECT 1809.800 2496.610 1811.390 2496.690 ;
        RECT 1809.740 2496.550 1811.390 2496.610 ;
        RECT 1809.740 2496.290 1810.000 2496.550 ;
        RECT 1811.110 2496.000 1811.390 2496.550 ;
        RECT 1128.020 2494.930 1128.280 2495.250 ;
        RECT 1128.080 827.890 1128.220 2494.930 ;
        RECT 14.820 827.570 15.080 827.890 ;
        RECT 1128.020 827.570 1128.280 827.890 ;
        RECT 14.880 825.365 15.020 827.570 ;
        RECT 14.810 824.995 15.090 825.365 ;
      LAYER via2 ;
        RECT 14.810 825.040 15.090 825.320 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 824.580 0.300 825.780 ;
=======
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 14.785 825.330 15.115 825.345 ;
        RECT -4.800 825.030 15.115 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
<<<<<<< HEAD
        RECT 18.925 825.015 19.255 825.030 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 14.785 825.015 15.115 825.030 ;
>>>>>>> re-updated local openlane
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1072.790 2508.080 1073.110 2508.140 ;
        RECT 1830.410 2508.080 1830.730 2508.140 ;
        RECT 1072.790 2507.940 1830.730 2508.080 ;
        RECT 1072.790 2507.880 1073.110 2507.940 ;
        RECT 1830.410 2507.880 1830.730 2507.940 ;
        RECT 14.790 613.940 15.110 614.000 ;
        RECT 1072.790 613.940 1073.110 614.000 ;
        RECT 14.790 613.800 1073.110 613.940 ;
        RECT 14.790 613.740 15.110 613.800 ;
        RECT 1072.790 613.740 1073.110 613.800 ;
      LAYER via ;
        RECT 1072.820 2507.880 1073.080 2508.140 ;
        RECT 1830.440 2507.880 1830.700 2508.140 ;
        RECT 14.820 613.740 15.080 614.000 ;
        RECT 1072.820 613.740 1073.080 614.000 ;
      LAYER met2 ;
        RECT 1072.820 2507.850 1073.080 2508.170 ;
        RECT 1830.440 2507.850 1830.700 2508.170 ;
        RECT 1072.880 614.030 1073.020 2507.850 ;
        RECT 1830.500 2500.000 1830.640 2507.850 ;
        RECT 1830.430 2496.000 1830.710 2500.000 ;
        RECT 14.820 613.710 15.080 614.030 ;
        RECT 1072.820 613.710 1073.080 614.030 ;
        RECT 14.880 610.485 15.020 613.710 ;
        RECT 14.810 610.115 15.090 610.485 ;
      LAYER via2 ;
        RECT 14.810 610.160 15.090 610.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 609.700 0.300 610.900 ;
=======
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 14.785 610.450 15.115 610.465 ;
        RECT -4.800 610.150 15.115 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
<<<<<<< HEAD
        RECT 18.005 610.135 18.335 610.150 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 14.785 610.135 15.115 610.150 ;
>>>>>>> re-updated local openlane
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1114.190 2500.260 1114.510 2500.320 ;
        RECT 1849.270 2500.260 1849.590 2500.320 ;
        RECT 1114.190 2500.120 1849.590 2500.260 ;
        RECT 1114.190 2500.060 1114.510 2500.120 ;
        RECT 1849.270 2500.060 1849.590 2500.120 ;
        RECT 16.170 400.080 16.490 400.140 ;
        RECT 1114.190 400.080 1114.510 400.140 ;
        RECT 16.170 399.940 1114.510 400.080 ;
        RECT 16.170 399.880 16.490 399.940 ;
        RECT 1114.190 399.880 1114.510 399.940 ;
      LAYER via ;
        RECT 1114.220 2500.060 1114.480 2500.320 ;
        RECT 1849.300 2500.060 1849.560 2500.320 ;
        RECT 16.200 399.880 16.460 400.140 ;
        RECT 1114.220 399.880 1114.480 400.140 ;
      LAYER met2 ;
        RECT 1114.220 2500.030 1114.480 2500.350 ;
        RECT 1849.300 2500.030 1849.560 2500.350 ;
        RECT 1114.280 400.170 1114.420 2500.030 ;
        RECT 1849.360 2499.410 1849.500 2500.030 ;
        RECT 1849.750 2499.410 1850.030 2500.000 ;
        RECT 1849.360 2499.270 1850.030 2499.410 ;
        RECT 1849.750 2496.000 1850.030 2499.270 ;
        RECT 16.200 399.850 16.460 400.170 ;
        RECT 1114.220 399.850 1114.480 400.170 ;
        RECT 16.260 394.925 16.400 399.850 ;
        RECT 16.190 394.555 16.470 394.925 ;
      LAYER via2 ;
        RECT 16.190 394.600 16.470 394.880 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT -4.800 394.140 0.300 395.340 ;
=======
        RECT 1252.390 2513.770 1252.770 2513.780 ;
        RECT 1867.205 2513.770 1867.535 2513.785 ;
        RECT 1252.390 2513.470 1867.535 2513.770 ;
        RECT 1252.390 2513.460 1252.770 2513.470 ;
        RECT 1867.205 2513.455 1867.535 2513.470 ;
        RECT 17.545 400.330 17.875 400.345 ;
        RECT 1252.390 400.330 1252.770 400.340 ;
        RECT 17.545 400.030 1252.770 400.330 ;
        RECT 17.545 400.015 17.875 400.030 ;
        RECT 1252.390 400.020 1252.770 400.030 ;
=======
>>>>>>> re-updated local openlane
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 16.165 394.890 16.495 394.905 ;
        RECT -4.800 394.590 16.495 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
<<<<<<< HEAD
        RECT 17.545 394.575 17.875 394.590 ;
      LAYER via3 ;
        RECT 1252.420 2513.460 1252.740 2513.780 ;
        RECT 1252.420 400.020 1252.740 400.340 ;
      LAYER met4 ;
        RECT 1252.415 2513.455 1252.745 2513.785 ;
        RECT 1252.430 400.345 1252.730 2513.455 ;
        RECT 1252.415 400.015 1252.745 400.345 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.165 394.575 16.495 394.590 ;
>>>>>>> re-updated local openlane
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1867.745 2493.645 1867.915 2496.535 ;
      LAYER mcon ;
        RECT 1867.745 2496.365 1867.915 2496.535 ;
      LAYER met1 ;
        RECT 1867.670 2496.520 1867.990 2496.580 ;
        RECT 1867.475 2496.380 1867.990 2496.520 ;
        RECT 1867.670 2496.320 1867.990 2496.380 ;
        RECT 1093.490 2493.800 1093.810 2493.860 ;
        RECT 1867.685 2493.800 1867.975 2493.845 ;
        RECT 1093.490 2493.660 1867.975 2493.800 ;
        RECT 1093.490 2493.600 1093.810 2493.660 ;
        RECT 1867.685 2493.615 1867.975 2493.660 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 1093.490 179.420 1093.810 179.480 ;
        RECT 17.090 179.280 1093.810 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 1093.490 179.220 1093.810 179.280 ;
      LAYER via ;
        RECT 1867.700 2496.320 1867.960 2496.580 ;
        RECT 1093.520 2493.600 1093.780 2493.860 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 1093.520 179.220 1093.780 179.480 ;
      LAYER met2 ;
        RECT 1869.070 2496.690 1869.350 2500.000 ;
        RECT 1867.760 2496.610 1869.350 2496.690 ;
        RECT 1867.700 2496.550 1869.350 2496.610 ;
        RECT 1867.700 2496.290 1867.960 2496.550 ;
        RECT 1869.070 2496.000 1869.350 2496.550 ;
        RECT 1093.520 2493.570 1093.780 2493.890 ;
        RECT 1093.580 179.510 1093.720 2493.570 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 1093.520 179.190 1093.780 179.510 ;
      LAYER via2 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT -4.800 178.580 0.300 179.780 ;
=======
        RECT 1251.470 2513.090 1251.850 2513.100 ;
        RECT 1886.985 2513.090 1887.315 2513.105 ;
        RECT 1251.470 2512.790 1887.315 2513.090 ;
        RECT 1251.470 2512.780 1251.850 2512.790 ;
        RECT 1886.985 2512.775 1887.315 2512.790 ;
=======
>>>>>>> re-updated local openlane
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
<<<<<<< HEAD
        RECT 1251.470 179.020 1251.850 179.030 ;
      LAYER via3 ;
        RECT 1251.500 2512.780 1251.820 2513.100 ;
        RECT 1251.500 179.020 1251.820 179.340 ;
      LAYER met4 ;
        RECT 1251.495 2512.775 1251.825 2513.105 ;
        RECT 1251.510 179.345 1251.810 2512.775 ;
        RECT 1251.495 179.015 1251.825 179.345 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 17.085 179.015 17.415 179.030 ;
>>>>>>> re-updated local openlane
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1211.250 2507.740 1211.570 2507.800 ;
        RECT 1990.490 2507.740 1990.810 2507.800 ;
        RECT 1211.250 2507.600 1990.810 2507.740 ;
        RECT 1211.250 2507.540 1211.570 2507.600 ;
        RECT 1990.490 2507.540 1990.810 2507.600 ;
        RECT 1990.490 793.460 1990.810 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 1990.490 793.320 2899.310 793.460 ;
        RECT 1990.490 793.260 1990.810 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 1211.280 2507.540 1211.540 2507.800 ;
        RECT 1990.520 2507.540 1990.780 2507.800 ;
        RECT 1990.520 793.260 1990.780 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 1211.280 2507.510 1211.540 2507.830 ;
        RECT 1990.520 2507.510 1990.780 2507.830 ;
        RECT 1211.340 2500.000 1211.480 2507.510 ;
        RECT 1211.270 2496.000 1211.550 2500.000 ;
        RECT 1990.580 793.550 1990.720 2507.510 ;
        RECT 1990.520 793.230 1990.780 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 791.260 2924.800 792.460 ;
=======
        RECT 1213.545 2498.140 1213.875 2498.145 ;
        RECT 1213.545 2498.130 1214.130 2498.140 ;
        RECT 1213.545 2497.830 1214.330 2498.130 ;
        RECT 1213.545 2497.820 1214.130 2497.830 ;
        RECT 1213.545 2497.815 1213.875 2497.820 ;
=======
        RECT 2898.985 792.010 2899.315 792.025 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
<<<<<<< HEAD
        RECT 2835.750 787.630 2883.890 787.930 ;
        RECT 2786.990 786.950 2788.210 787.250 ;
        RECT 2883.590 787.250 2883.890 787.630 ;
        RECT 2884.510 787.630 2917.010 787.930 ;
        RECT 2884.510 787.250 2884.810 787.630 ;
        RECT 2883.590 786.950 2884.810 787.250 ;
        RECT 2052.585 786.935 2052.915 786.950 ;
        RECT 1895.265 785.590 1931.690 785.890 ;
        RECT 1895.265 785.575 1895.595 785.590 ;
      LAYER via3 ;
        RECT 1213.780 2497.820 1214.100 2498.140 ;
        RECT 1980.140 789.660 1980.460 789.980 ;
        RECT 1213.780 786.940 1214.100 787.260 ;
        RECT 1980.140 788.300 1980.460 788.620 ;
      LAYER met4 ;
        RECT 1213.775 2497.815 1214.105 2498.145 ;
        RECT 1213.790 787.265 1214.090 2497.815 ;
        RECT 1980.135 789.655 1980.465 789.985 ;
        RECT 1980.150 788.625 1980.450 789.655 ;
        RECT 1980.135 788.295 1980.465 788.625 ;
        RECT 1213.775 786.935 1214.105 787.265 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1232.485 2493.305 1232.655 2496.535 ;
      LAYER mcon ;
        RECT 1232.485 2496.365 1232.655 2496.535 ;
      LAYER met1 ;
        RECT 1232.410 2496.520 1232.730 2496.580 ;
        RECT 1232.215 2496.380 1232.730 2496.520 ;
        RECT 1232.410 2496.320 1232.730 2496.380 ;
        RECT 1232.425 2493.460 1232.715 2493.505 ;
        RECT 2045.690 2493.460 2046.010 2493.520 ;
        RECT 1232.425 2493.320 2046.010 2493.460 ;
        RECT 1232.425 2493.275 1232.715 2493.320 ;
        RECT 2045.690 2493.260 2046.010 2493.320 ;
        RECT 2045.690 1028.060 2046.010 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 2045.690 1027.920 2899.310 1028.060 ;
        RECT 2045.690 1027.860 2046.010 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 1232.440 2496.320 1232.700 2496.580 ;
        RECT 2045.720 2493.260 2045.980 2493.520 ;
        RECT 2045.720 1027.860 2045.980 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 1230.590 2496.690 1230.870 2500.000 ;
        RECT 1230.590 2496.610 1232.640 2496.690 ;
        RECT 1230.590 2496.550 1232.700 2496.610 ;
        RECT 1230.590 2496.000 1230.870 2496.550 ;
        RECT 1232.440 2496.290 1232.700 2496.550 ;
        RECT 2045.720 2493.230 2045.980 2493.550 ;
        RECT 2045.780 1028.150 2045.920 2493.230 ;
        RECT 2045.720 1027.830 2045.980 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1025.860 2924.800 1027.060 ;
=======
        RECT 1233.785 2498.140 1234.115 2498.145 ;
        RECT 1233.785 2498.130 1234.370 2498.140 ;
        RECT 1233.785 2497.830 1234.570 2498.130 ;
        RECT 1233.785 2497.820 1234.370 2497.830 ;
        RECT 1233.785 2497.815 1234.115 2497.820 ;
=======
        RECT 2898.985 1026.610 2899.315 1026.625 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
<<<<<<< HEAD
        RECT 2835.750 1022.230 2883.890 1022.530 ;
        RECT 2786.990 1021.550 2788.210 1021.850 ;
        RECT 2883.590 1021.850 2883.890 1022.230 ;
        RECT 2884.510 1022.230 2917.010 1022.530 ;
        RECT 2884.510 1021.850 2884.810 1022.230 ;
        RECT 2883.590 1021.550 2884.810 1021.850 ;
        RECT 2052.585 1021.535 2052.915 1021.550 ;
        RECT 1895.265 1020.190 1931.690 1020.490 ;
        RECT 1895.265 1020.175 1895.595 1020.190 ;
      LAYER via3 ;
        RECT 1234.020 2497.820 1234.340 2498.140 ;
        RECT 1234.020 1023.580 1234.340 1023.900 ;
        RECT 1980.140 1024.260 1980.460 1024.580 ;
        RECT 1441.940 1023.580 1442.260 1023.900 ;
        RECT 1441.940 1022.220 1442.260 1022.540 ;
        RECT 1980.140 1022.900 1980.460 1023.220 ;
      LAYER met4 ;
        RECT 1234.015 2497.815 1234.345 2498.145 ;
        RECT 1234.030 1023.905 1234.330 2497.815 ;
        RECT 1980.135 1024.255 1980.465 1024.585 ;
        RECT 1234.015 1023.575 1234.345 1023.905 ;
        RECT 1441.935 1023.575 1442.265 1023.905 ;
        RECT 1441.950 1022.545 1442.250 1023.575 ;
        RECT 1980.150 1023.225 1980.450 1024.255 ;
        RECT 1980.135 1022.895 1980.465 1023.225 ;
        RECT 1441.935 1022.215 1442.265 1022.545 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2186.910 1257.560 2187.230 1257.620 ;
        RECT 2221.410 1257.560 2221.730 1257.620 ;
        RECT 2186.910 1257.420 2221.730 1257.560 ;
        RECT 2186.910 1257.360 2187.230 1257.420 ;
        RECT 2221.410 1257.360 2221.730 1257.420 ;
        RECT 2456.470 1257.560 2456.790 1257.620 ;
        RECT 2504.310 1257.560 2504.630 1257.620 ;
        RECT 2456.470 1257.420 2504.630 1257.560 ;
        RECT 2456.470 1257.360 2456.790 1257.420 ;
        RECT 2504.310 1257.360 2504.630 1257.420 ;
        RECT 1799.130 1257.220 1799.450 1257.280 ;
        RECT 1800.970 1257.220 1801.290 1257.280 ;
        RECT 1799.130 1257.080 1801.290 1257.220 ;
        RECT 1799.130 1257.020 1799.450 1257.080 ;
        RECT 1800.970 1257.020 1801.290 1257.080 ;
        RECT 1883.770 1257.220 1884.090 1257.280 ;
        RECT 1929.770 1257.220 1930.090 1257.280 ;
        RECT 1883.770 1257.080 1930.090 1257.220 ;
        RECT 1883.770 1257.020 1884.090 1257.080 ;
        RECT 1929.770 1257.020 1930.090 1257.080 ;
        RECT 1932.070 1257.220 1932.390 1257.280 ;
        RECT 1970.250 1257.220 1970.570 1257.280 ;
        RECT 1932.070 1257.080 1970.570 1257.220 ;
        RECT 1932.070 1257.020 1932.390 1257.080 ;
        RECT 1970.250 1257.020 1970.570 1257.080 ;
        RECT 2621.610 1256.880 2621.930 1256.940 ;
        RECT 2622.530 1256.880 2622.850 1256.940 ;
        RECT 2621.610 1256.740 2622.850 1256.880 ;
        RECT 2621.610 1256.680 2621.930 1256.740 ;
        RECT 2622.530 1256.680 2622.850 1256.740 ;
        RECT 1606.390 1256.540 1606.710 1256.600 ;
        RECT 1639.970 1256.540 1640.290 1256.600 ;
        RECT 1606.390 1256.400 1640.290 1256.540 ;
        RECT 1606.390 1256.340 1606.710 1256.400 ;
        RECT 1639.970 1256.340 1640.290 1256.400 ;
        RECT 1642.270 1256.540 1642.590 1256.600 ;
        RECT 1690.110 1256.540 1690.430 1256.600 ;
        RECT 1642.270 1256.400 1690.430 1256.540 ;
        RECT 1642.270 1256.340 1642.590 1256.400 ;
        RECT 1690.110 1256.340 1690.430 1256.400 ;
        RECT 2649.670 1256.540 2649.990 1256.600 ;
        RECT 2697.510 1256.540 2697.830 1256.600 ;
        RECT 2649.670 1256.400 2697.830 1256.540 ;
        RECT 2649.670 1256.340 2649.990 1256.400 ;
        RECT 2697.510 1256.340 2697.830 1256.400 ;
      LAYER via ;
        RECT 2186.940 1257.360 2187.200 1257.620 ;
        RECT 2221.440 1257.360 2221.700 1257.620 ;
        RECT 2456.500 1257.360 2456.760 1257.620 ;
        RECT 2504.340 1257.360 2504.600 1257.620 ;
        RECT 1799.160 1257.020 1799.420 1257.280 ;
        RECT 1801.000 1257.020 1801.260 1257.280 ;
        RECT 1883.800 1257.020 1884.060 1257.280 ;
        RECT 1929.800 1257.020 1930.060 1257.280 ;
        RECT 1932.100 1257.020 1932.360 1257.280 ;
        RECT 1970.280 1257.020 1970.540 1257.280 ;
        RECT 2621.640 1256.680 2621.900 1256.940 ;
        RECT 2622.560 1256.680 2622.820 1256.940 ;
        RECT 1606.420 1256.340 1606.680 1256.600 ;
        RECT 1640.000 1256.340 1640.260 1256.600 ;
        RECT 1642.300 1256.340 1642.560 1256.600 ;
        RECT 1690.140 1256.340 1690.400 1256.600 ;
        RECT 2649.700 1256.340 2649.960 1256.600 ;
        RECT 2697.540 1256.340 2697.800 1256.600 ;
      LAYER met2 ;
        RECT 1249.910 2498.050 1250.190 2500.000 ;
        RECT 1251.750 2498.050 1252.030 2498.165 ;
        RECT 1249.910 2497.910 1252.030 2498.050 ;
        RECT 1249.910 2496.000 1250.190 2497.910 ;
        RECT 1251.750 2497.795 1252.030 2497.910 ;
        RECT 1562.710 1258.835 1562.990 1259.205 ;
        RECT 2304.230 1258.835 2304.510 1259.205 ;
        RECT 1562.780 1257.845 1562.920 1258.835 ;
        RECT 1970.270 1258.155 1970.550 1258.525 ;
        RECT 1562.710 1257.475 1562.990 1257.845 ;
        RECT 1690.130 1257.475 1690.410 1257.845 ;
        RECT 1883.790 1257.475 1884.070 1257.845 ;
        RECT 1606.410 1256.795 1606.690 1257.165 ;
        RECT 1606.480 1256.630 1606.620 1256.795 ;
        RECT 1606.420 1256.310 1606.680 1256.630 ;
        RECT 1639.990 1256.285 1640.270 1256.655 ;
        RECT 1690.200 1256.630 1690.340 1257.475 ;
        RECT 1883.860 1257.310 1884.000 1257.475 ;
        RECT 1799.160 1257.165 1799.420 1257.310 ;
        RECT 1801.000 1257.165 1801.260 1257.310 ;
        RECT 1799.150 1256.795 1799.430 1257.165 ;
        RECT 1800.990 1256.795 1801.270 1257.165 ;
        RECT 1883.800 1256.990 1884.060 1257.310 ;
        RECT 1929.790 1256.965 1930.070 1257.335 ;
        RECT 1970.340 1257.310 1970.480 1258.155 ;
        RECT 2304.300 1257.845 2304.440 1258.835 ;
        RECT 2186.930 1257.475 2187.210 1257.845 ;
        RECT 2221.430 1257.475 2221.710 1257.845 ;
        RECT 2304.230 1257.475 2304.510 1257.845 ;
        RECT 2186.940 1257.330 2187.200 1257.475 ;
        RECT 2221.440 1257.330 2221.700 1257.475 ;
        RECT 2456.500 1257.330 2456.760 1257.650 ;
        RECT 2504.330 1257.475 2504.610 1257.845 ;
        RECT 2697.530 1257.475 2697.810 1257.845 ;
        RECT 2504.340 1257.330 2504.600 1257.475 ;
        RECT 1932.100 1257.165 1932.360 1257.310 ;
        RECT 1932.090 1256.795 1932.370 1257.165 ;
        RECT 1970.280 1256.990 1970.540 1257.310 ;
        RECT 2456.560 1257.165 2456.700 1257.330 ;
        RECT 1993.730 1257.050 1994.010 1257.165 ;
        RECT 1994.650 1257.050 1994.930 1257.165 ;
        RECT 1993.730 1256.910 1994.930 1257.050 ;
        RECT 1993.730 1256.795 1994.010 1256.910 ;
        RECT 1994.650 1256.795 1994.930 1256.910 ;
        RECT 2456.490 1256.795 2456.770 1257.165 ;
        RECT 2574.250 1257.050 2574.530 1257.165 ;
        RECT 2573.400 1256.910 2574.530 1257.050 ;
        RECT 1642.300 1256.485 1642.560 1256.630 ;
        RECT 1642.290 1256.115 1642.570 1256.485 ;
        RECT 1690.140 1256.310 1690.400 1256.630 ;
        RECT 2573.400 1256.485 2573.540 1256.910 ;
        RECT 2574.250 1256.795 2574.530 1256.910 ;
        RECT 2621.630 1256.795 2621.910 1257.165 ;
        RECT 2621.640 1256.650 2621.900 1256.795 ;
        RECT 2622.560 1256.650 2622.820 1256.970 ;
        RECT 2622.620 1256.485 2622.760 1256.650 ;
        RECT 2697.600 1256.630 2697.740 1257.475 ;
        RECT 2649.700 1256.485 2649.960 1256.630 ;
        RECT 2573.330 1256.115 2573.610 1256.485 ;
        RECT 2622.550 1256.115 2622.830 1256.485 ;
        RECT 2649.690 1256.115 2649.970 1256.485 ;
        RECT 2697.540 1256.310 2697.800 1256.630 ;
      LAYER via2 ;
        RECT 1251.750 2497.840 1252.030 2498.120 ;
        RECT 1562.710 1258.880 1562.990 1259.160 ;
        RECT 2304.230 1258.880 2304.510 1259.160 ;
        RECT 1970.270 1258.200 1970.550 1258.480 ;
        RECT 1562.710 1257.520 1562.990 1257.800 ;
        RECT 1690.130 1257.520 1690.410 1257.800 ;
        RECT 1883.790 1257.520 1884.070 1257.800 ;
        RECT 1606.410 1256.840 1606.690 1257.120 ;
        RECT 1799.150 1256.840 1799.430 1257.120 ;
        RECT 1800.990 1256.840 1801.270 1257.120 ;
        RECT 2186.930 1257.520 2187.210 1257.800 ;
        RECT 2221.430 1257.520 2221.710 1257.800 ;
        RECT 2304.230 1257.520 2304.510 1257.800 ;
        RECT 2504.330 1257.520 2504.610 1257.800 ;
        RECT 2697.530 1257.520 2697.810 1257.800 ;
        RECT 1929.790 1257.010 1930.070 1257.290 ;
        RECT 1932.090 1256.840 1932.370 1257.120 ;
        RECT 1993.730 1256.840 1994.010 1257.120 ;
        RECT 1994.650 1256.840 1994.930 1257.120 ;
        RECT 2456.490 1256.840 2456.770 1257.120 ;
        RECT 1639.990 1256.330 1640.270 1256.610 ;
        RECT 1642.290 1256.160 1642.570 1256.440 ;
        RECT 2574.250 1256.840 2574.530 1257.120 ;
        RECT 2621.630 1256.840 2621.910 1257.120 ;
        RECT 2573.330 1256.160 2573.610 1256.440 ;
        RECT 2622.550 1256.160 2622.830 1256.440 ;
        RECT 2649.690 1256.160 2649.970 1256.440 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1260.460 2924.800 1261.660 ;
=======
        RECT 1253.565 2498.130 1253.895 2498.145 ;
=======
        RECT 1251.725 2498.130 1252.055 2498.145 ;
>>>>>>> re-updated local openlane
        RECT 1255.150 2498.130 1255.530 2498.140 ;
        RECT 1251.725 2497.830 1255.530 2498.130 ;
        RECT 1251.725 2497.815 1252.055 2497.830 ;
        RECT 1255.150 2497.820 1255.530 2497.830 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2916.710 1260.910 2924.800 1261.210 ;
        RECT 1538.510 1259.170 1538.890 1259.180 ;
        RECT 1562.685 1259.170 1563.015 1259.185 ;
        RECT 1538.510 1258.870 1563.015 1259.170 ;
        RECT 1538.510 1258.860 1538.890 1258.870 ;
        RECT 1562.685 1258.855 1563.015 1258.870 ;
        RECT 2269.910 1259.170 2270.290 1259.180 ;
        RECT 2304.205 1259.170 2304.535 1259.185 ;
        RECT 2269.910 1258.870 2304.535 1259.170 ;
        RECT 2269.910 1258.860 2270.290 1258.870 ;
        RECT 2304.205 1258.855 2304.535 1258.870 ;
        RECT 1970.245 1258.490 1970.575 1258.505 ;
        RECT 1980.110 1258.490 1980.490 1258.500 ;
        RECT 1970.245 1258.190 1980.490 1258.490 ;
        RECT 1970.245 1258.175 1970.575 1258.190 ;
        RECT 1980.110 1258.180 1980.490 1258.190 ;
        RECT 1441.910 1257.810 1442.290 1257.820 ;
        RECT 1538.510 1257.810 1538.890 1257.820 ;
        RECT 1280.030 1257.510 1318.970 1257.810 ;
        RECT 1255.150 1257.130 1255.530 1257.140 ;
        RECT 1255.150 1256.830 1269.290 1257.130 ;
        RECT 1255.150 1256.820 1255.530 1256.830 ;
        RECT 1268.990 1256.450 1269.290 1256.830 ;
        RECT 1280.030 1256.450 1280.330 1257.510 ;
        RECT 1268.990 1256.150 1280.330 1256.450 ;
        RECT 1318.670 1256.450 1318.970 1257.510 ;
        RECT 1365.590 1257.510 1366.810 1257.810 ;
        RECT 1365.590 1256.450 1365.890 1257.510 ;
        RECT 1366.510 1257.130 1366.810 1257.510 ;
        RECT 1441.910 1257.510 1538.890 1257.810 ;
        RECT 1441.910 1257.500 1442.290 1257.510 ;
        RECT 1538.510 1257.500 1538.890 1257.510 ;
        RECT 1562.685 1257.810 1563.015 1257.825 ;
        RECT 1690.105 1257.810 1690.435 1257.825 ;
        RECT 1883.765 1257.810 1884.095 1257.825 ;
        RECT 2186.905 1257.810 2187.235 1257.825 ;
        RECT 1562.685 1257.510 1586.690 1257.810 ;
        RECT 1562.685 1257.495 1563.015 1257.510 ;
        RECT 1586.390 1257.130 1586.690 1257.510 ;
        RECT 1690.105 1257.510 1704.450 1257.810 ;
        RECT 1690.105 1257.495 1690.435 1257.510 ;
        RECT 1606.385 1257.130 1606.715 1257.145 ;
        RECT 1366.510 1256.830 1424.770 1257.130 ;
        RECT 1586.390 1256.830 1606.715 1257.130 ;
        RECT 1318.670 1256.150 1365.890 1256.450 ;
        RECT 1424.470 1256.450 1424.770 1256.830 ;
        RECT 1606.385 1256.815 1606.715 1256.830 ;
        RECT 1639.965 1256.620 1640.295 1256.635 ;
        RECT 1441.910 1256.450 1442.290 1256.460 ;
        RECT 1424.470 1256.150 1442.290 1256.450 ;
        RECT 1639.965 1256.450 1641.890 1256.620 ;
        RECT 1642.265 1256.450 1642.595 1256.465 ;
        RECT 1639.965 1256.320 1642.595 1256.450 ;
        RECT 1639.965 1256.305 1640.295 1256.320 ;
        RECT 1641.590 1256.150 1642.595 1256.320 ;
        RECT 1704.150 1256.450 1704.450 1257.510 ;
        RECT 1849.510 1257.510 1884.095 1257.810 ;
        RECT 1799.125 1257.130 1799.455 1257.145 ;
        RECT 1752.910 1256.830 1799.455 1257.130 ;
        RECT 1752.910 1256.450 1753.210 1256.830 ;
        RECT 1799.125 1256.815 1799.455 1256.830 ;
        RECT 1800.965 1257.130 1801.295 1257.145 ;
        RECT 1800.965 1256.830 1835.090 1257.130 ;
        RECT 1800.965 1256.815 1801.295 1256.830 ;
        RECT 1704.150 1256.150 1753.210 1256.450 ;
        RECT 1834.790 1256.450 1835.090 1256.830 ;
        RECT 1849.510 1256.450 1849.810 1257.510 ;
        RECT 1883.765 1257.495 1884.095 1257.510 ;
        RECT 2062.950 1257.510 2111.090 1257.810 ;
        RECT 1929.765 1257.300 1930.095 1257.315 ;
        RECT 1929.765 1257.130 1931.690 1257.300 ;
        RECT 1932.065 1257.130 1932.395 1257.145 ;
        RECT 1929.765 1257.000 1932.395 1257.130 ;
        RECT 1929.765 1256.985 1930.095 1257.000 ;
        RECT 1931.390 1256.830 1932.395 1257.000 ;
        RECT 1932.065 1256.815 1932.395 1256.830 ;
        RECT 1980.110 1257.130 1980.490 1257.140 ;
        RECT 1993.705 1257.130 1994.035 1257.145 ;
        RECT 1980.110 1256.830 1994.035 1257.130 ;
        RECT 1980.110 1256.820 1980.490 1256.830 ;
        RECT 1993.705 1256.815 1994.035 1256.830 ;
        RECT 1994.625 1257.130 1994.955 1257.145 ;
        RECT 1994.625 1256.830 2042.090 1257.130 ;
        RECT 1994.625 1256.815 1994.955 1256.830 ;
        RECT 1834.790 1256.150 1849.810 1256.450 ;
        RECT 2041.790 1256.450 2042.090 1256.830 ;
        RECT 2062.950 1256.450 2063.250 1257.510 ;
        RECT 2041.790 1256.150 2063.250 1256.450 ;
        RECT 2110.790 1256.450 2111.090 1257.510 ;
        RECT 2111.710 1257.510 2187.235 1257.810 ;
        RECT 2111.710 1256.450 2112.010 1257.510 ;
        RECT 2186.905 1257.495 2187.235 1257.510 ;
        RECT 2221.405 1257.810 2221.735 1257.825 ;
        RECT 2304.205 1257.810 2304.535 1257.825 ;
        RECT 2504.305 1257.810 2504.635 1257.825 ;
        RECT 2697.505 1257.810 2697.835 1257.825 ;
        RECT 2221.405 1257.510 2235.290 1257.810 ;
        RECT 2221.405 1257.495 2221.735 1257.510 ;
        RECT 2110.790 1256.150 2112.010 1256.450 ;
        RECT 2234.990 1256.450 2235.290 1257.510 ;
        RECT 2304.205 1257.510 2353.050 1257.810 ;
        RECT 2304.205 1257.495 2304.535 1257.510 ;
        RECT 2269.910 1257.130 2270.290 1257.140 ;
        RECT 2235.910 1256.830 2270.290 1257.130 ;
        RECT 2352.750 1257.130 2353.050 1257.510 ;
        RECT 2401.510 1257.510 2429.410 1257.810 ;
        RECT 2352.750 1256.830 2400.890 1257.130 ;
        RECT 2235.910 1256.450 2236.210 1256.830 ;
        RECT 2269.910 1256.820 2270.290 1256.830 ;
        RECT 2234.990 1256.150 2236.210 1256.450 ;
        RECT 2400.590 1256.450 2400.890 1256.830 ;
        RECT 2401.510 1256.450 2401.810 1257.510 ;
        RECT 2429.110 1257.130 2429.410 1257.510 ;
        RECT 2504.305 1257.510 2526.010 1257.810 ;
        RECT 2504.305 1257.495 2504.635 1257.510 ;
        RECT 2456.465 1257.130 2456.795 1257.145 ;
        RECT 2429.110 1256.830 2456.795 1257.130 ;
        RECT 2456.465 1256.815 2456.795 1256.830 ;
        RECT 2400.590 1256.150 2401.810 1256.450 ;
        RECT 2525.710 1256.450 2526.010 1257.510 ;
        RECT 2697.505 1257.510 2739.450 1257.810 ;
        RECT 2697.505 1257.495 2697.835 1257.510 ;
        RECT 2574.225 1257.130 2574.555 1257.145 ;
        RECT 2621.605 1257.130 2621.935 1257.145 ;
        RECT 2574.225 1256.830 2621.935 1257.130 ;
        RECT 2739.150 1257.130 2739.450 1257.510 ;
        RECT 2787.910 1257.510 2836.050 1257.810 ;
        RECT 2739.150 1256.830 2787.290 1257.130 ;
        RECT 2574.225 1256.815 2574.555 1256.830 ;
        RECT 2621.605 1256.815 2621.935 1256.830 ;
        RECT 2573.305 1256.450 2573.635 1256.465 ;
        RECT 2525.710 1256.150 2573.635 1256.450 ;
        RECT 1441.910 1256.140 1442.290 1256.150 ;
        RECT 1642.265 1256.135 1642.595 1256.150 ;
        RECT 2573.305 1256.135 2573.635 1256.150 ;
        RECT 2622.525 1256.450 2622.855 1256.465 ;
        RECT 2649.665 1256.450 2649.995 1256.465 ;
        RECT 2622.525 1256.150 2649.995 1256.450 ;
        RECT 2786.990 1256.450 2787.290 1256.830 ;
        RECT 2787.910 1256.450 2788.210 1257.510 ;
        RECT 2835.750 1257.130 2836.050 1257.510 ;
        RECT 2916.710 1257.130 2917.010 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2835.750 1256.830 2883.890 1257.130 ;
        RECT 2786.990 1256.150 2788.210 1256.450 ;
        RECT 2883.590 1256.450 2883.890 1256.830 ;
        RECT 2884.510 1256.830 2917.010 1257.130 ;
        RECT 2884.510 1256.450 2884.810 1256.830 ;
        RECT 2883.590 1256.150 2884.810 1256.450 ;
        RECT 2622.525 1256.135 2622.855 1256.150 ;
        RECT 2649.665 1256.135 2649.995 1256.150 ;
      LAYER via3 ;
        RECT 1255.180 2497.820 1255.500 2498.140 ;
        RECT 1538.540 1258.860 1538.860 1259.180 ;
        RECT 2269.940 1258.860 2270.260 1259.180 ;
        RECT 1980.140 1258.180 1980.460 1258.500 ;
        RECT 1255.180 1256.820 1255.500 1257.140 ;
        RECT 1441.940 1257.500 1442.260 1257.820 ;
        RECT 1538.540 1257.500 1538.860 1257.820 ;
        RECT 1441.940 1256.140 1442.260 1256.460 ;
        RECT 1980.140 1256.820 1980.460 1257.140 ;
        RECT 2269.940 1256.820 2270.260 1257.140 ;
      LAYER met4 ;
        RECT 1255.175 2497.815 1255.505 2498.145 ;
<<<<<<< HEAD
        RECT 1255.190 1256.465 1255.490 2497.815 ;
        RECT 1442.855 1257.495 1443.185 1257.825 ;
        RECT 1255.175 1256.135 1255.505 1256.465 ;
        RECT 1441.935 1256.450 1442.265 1256.465 ;
        RECT 1442.870 1256.450 1443.170 1257.495 ;
        RECT 1441.935 1256.150 1443.170 1256.450 ;
        RECT 1441.935 1256.135 1442.265 1256.150 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1255.190 1257.145 1255.490 2497.815 ;
        RECT 1538.535 1258.855 1538.865 1259.185 ;
        RECT 2269.935 1258.855 2270.265 1259.185 ;
        RECT 1538.550 1257.825 1538.850 1258.855 ;
        RECT 1980.135 1258.175 1980.465 1258.505 ;
        RECT 1441.935 1257.495 1442.265 1257.825 ;
        RECT 1538.535 1257.495 1538.865 1257.825 ;
        RECT 1255.175 1256.815 1255.505 1257.145 ;
        RECT 1441.950 1256.465 1442.250 1257.495 ;
        RECT 1980.150 1257.145 1980.450 1258.175 ;
        RECT 2269.950 1257.145 2270.250 1258.855 ;
        RECT 1980.135 1256.815 1980.465 1257.145 ;
        RECT 2269.935 1256.815 2270.265 1257.145 ;
        RECT 1441.935 1256.135 1442.265 1256.465 ;
>>>>>>> re-updated local openlane
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1269.210 2500.600 1269.530 2500.660 ;
        RECT 1997.850 2500.600 1998.170 2500.660 ;
        RECT 1269.210 2500.460 1998.170 2500.600 ;
        RECT 1269.210 2500.400 1269.530 2500.460 ;
        RECT 1997.850 2500.400 1998.170 2500.460 ;
        RECT 1997.850 1497.260 1998.170 1497.320 ;
        RECT 2898.990 1497.260 2899.310 1497.320 ;
        RECT 1997.850 1497.120 2899.310 1497.260 ;
        RECT 1997.850 1497.060 1998.170 1497.120 ;
        RECT 2898.990 1497.060 2899.310 1497.120 ;
      LAYER via ;
        RECT 1269.240 2500.400 1269.500 2500.660 ;
        RECT 1997.880 2500.400 1998.140 2500.660 ;
        RECT 1997.880 1497.060 1998.140 1497.320 ;
        RECT 2899.020 1497.060 2899.280 1497.320 ;
      LAYER met2 ;
        RECT 1269.240 2500.370 1269.500 2500.690 ;
        RECT 1997.880 2500.370 1998.140 2500.690 ;
        RECT 1269.300 2500.000 1269.440 2500.370 ;
        RECT 1269.230 2496.000 1269.510 2500.000 ;
        RECT 1997.940 1497.350 1998.080 2500.370 ;
        RECT 1997.880 1497.030 1998.140 1497.350 ;
        RECT 2899.020 1497.030 2899.280 1497.350 ;
        RECT 2899.080 1495.845 2899.220 1497.030 ;
        RECT 2899.010 1495.475 2899.290 1495.845 ;
      LAYER via2 ;
        RECT 2899.010 1495.520 2899.290 1495.800 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1495.060 2924.800 1496.260 ;
=======
        RECT 1273.805 2498.130 1274.135 2498.145 ;
        RECT 1275.390 2498.130 1275.770 2498.140 ;
        RECT 1273.805 2497.830 1275.770 2498.130 ;
        RECT 1273.805 2497.815 1274.135 2497.830 ;
        RECT 1275.390 2497.820 1275.770 2497.830 ;
=======
        RECT 2898.985 1495.810 2899.315 1495.825 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.985 1495.510 2924.800 1495.810 ;
        RECT 2898.985 1495.495 2899.315 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
<<<<<<< HEAD
        RECT 2835.750 1491.430 2883.890 1491.730 ;
        RECT 2786.990 1490.750 2788.210 1491.050 ;
        RECT 2883.590 1491.050 2883.890 1491.430 ;
        RECT 2884.510 1491.430 2917.010 1491.730 ;
        RECT 2884.510 1491.050 2884.810 1491.430 ;
        RECT 2883.590 1490.750 2884.810 1491.050 ;
        RECT 2052.585 1490.735 2052.915 1490.750 ;
        RECT 1895.265 1489.390 1931.690 1489.690 ;
        RECT 1895.265 1489.375 1895.595 1489.390 ;
      LAYER via3 ;
        RECT 1275.420 2497.820 1275.740 2498.140 ;
        RECT 1980.140 1493.460 1980.460 1493.780 ;
        RECT 1435.500 1492.780 1435.820 1493.100 ;
        RECT 1275.420 1492.100 1275.740 1492.420 ;
        RECT 1435.500 1491.420 1435.820 1491.740 ;
        RECT 1980.140 1492.100 1980.460 1492.420 ;
      LAYER met4 ;
        RECT 1275.415 2497.815 1275.745 2498.145 ;
        RECT 1275.430 1492.425 1275.730 2497.815 ;
        RECT 1980.135 1493.455 1980.465 1493.785 ;
        RECT 1435.495 1492.775 1435.825 1493.105 ;
        RECT 1275.415 1492.095 1275.745 1492.425 ;
        RECT 1435.510 1491.745 1435.810 1492.775 ;
        RECT 1980.150 1492.425 1980.450 1493.455 ;
        RECT 1980.135 1492.095 1980.465 1492.425 ;
        RECT 1435.495 1491.415 1435.825 1491.745 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1288.530 2508.760 1288.850 2508.820 ;
        RECT 2011.650 2508.760 2011.970 2508.820 ;
        RECT 1288.530 2508.620 2011.970 2508.760 ;
        RECT 1288.530 2508.560 1288.850 2508.620 ;
        RECT 2011.650 2508.560 2011.970 2508.620 ;
        RECT 2011.650 1731.860 2011.970 1731.920 ;
        RECT 2900.830 1731.860 2901.150 1731.920 ;
        RECT 2011.650 1731.720 2901.150 1731.860 ;
        RECT 2011.650 1731.660 2011.970 1731.720 ;
        RECT 2900.830 1731.660 2901.150 1731.720 ;
      LAYER via ;
        RECT 1288.560 2508.560 1288.820 2508.820 ;
        RECT 2011.680 2508.560 2011.940 2508.820 ;
        RECT 2011.680 1731.660 2011.940 1731.920 ;
        RECT 2900.860 1731.660 2901.120 1731.920 ;
      LAYER met2 ;
        RECT 1288.560 2508.530 1288.820 2508.850 ;
        RECT 2011.680 2508.530 2011.940 2508.850 ;
        RECT 1288.620 2500.000 1288.760 2508.530 ;
        RECT 1288.550 2496.000 1288.830 2500.000 ;
        RECT 2011.740 1731.950 2011.880 2508.530 ;
        RECT 2011.680 1731.630 2011.940 1731.950 ;
        RECT 2900.860 1731.630 2901.120 1731.950 ;
        RECT 2900.920 1730.445 2901.060 1731.630 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1729.660 2924.800 1730.860 ;
=======
        RECT 2901.285 1730.410 2901.615 1730.425 ;
=======
        RECT 2900.825 1730.410 2901.155 1730.425 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1309.765 2494.325 1309.935 2496.535 ;
      LAYER mcon ;
        RECT 1309.765 2496.365 1309.935 2496.535 ;
      LAYER met1 ;
        RECT 1309.690 2496.520 1310.010 2496.580 ;
        RECT 1309.495 2496.380 1310.010 2496.520 ;
        RECT 1309.690 2496.320 1310.010 2496.380 ;
        RECT 1309.705 2494.480 1309.995 2494.525 ;
        RECT 2052.590 2494.480 2052.910 2494.540 ;
        RECT 1309.705 2494.340 2052.910 2494.480 ;
        RECT 1309.705 2494.295 1309.995 2494.340 ;
        RECT 2052.590 2494.280 2052.910 2494.340 ;
        RECT 2052.590 1966.460 2052.910 1966.520 ;
        RECT 2900.830 1966.460 2901.150 1966.520 ;
        RECT 2052.590 1966.320 2901.150 1966.460 ;
        RECT 2052.590 1966.260 2052.910 1966.320 ;
        RECT 2900.830 1966.260 2901.150 1966.320 ;
      LAYER via ;
        RECT 1309.720 2496.320 1309.980 2496.580 ;
        RECT 2052.620 2494.280 2052.880 2494.540 ;
        RECT 2052.620 1966.260 2052.880 1966.520 ;
        RECT 2900.860 1966.260 2901.120 1966.520 ;
      LAYER met2 ;
        RECT 1307.870 2496.690 1308.150 2500.000 ;
        RECT 1307.870 2496.610 1309.920 2496.690 ;
        RECT 1307.870 2496.550 1309.980 2496.610 ;
        RECT 1307.870 2496.000 1308.150 2496.550 ;
        RECT 1309.720 2496.290 1309.980 2496.550 ;
        RECT 2052.620 2494.250 2052.880 2494.570 ;
        RECT 2052.680 1966.550 2052.820 2494.250 ;
        RECT 2052.620 1966.230 2052.880 1966.550 ;
        RECT 2900.860 1966.230 2901.120 1966.550 ;
        RECT 2900.920 1965.045 2901.060 1966.230 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1964.260 2924.800 1965.460 ;
=======
        RECT 2898.065 1965.010 2898.395 1965.025 ;
=======
        RECT 2900.825 1965.010 2901.155 1965.025 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1327.170 2501.620 1327.490 2501.680 ;
        RECT 2032.350 2501.620 2032.670 2501.680 ;
        RECT 1327.170 2501.480 2032.670 2501.620 ;
        RECT 1327.170 2501.420 1327.490 2501.480 ;
        RECT 2032.350 2501.420 2032.670 2501.480 ;
        RECT 2032.350 2201.060 2032.670 2201.120 ;
        RECT 2900.830 2201.060 2901.150 2201.120 ;
        RECT 2032.350 2200.920 2901.150 2201.060 ;
        RECT 2032.350 2200.860 2032.670 2200.920 ;
        RECT 2900.830 2200.860 2901.150 2200.920 ;
      LAYER via ;
        RECT 1327.200 2501.420 1327.460 2501.680 ;
        RECT 2032.380 2501.420 2032.640 2501.680 ;
        RECT 2032.380 2200.860 2032.640 2201.120 ;
        RECT 2900.860 2200.860 2901.120 2201.120 ;
      LAYER met2 ;
        RECT 1327.200 2501.390 1327.460 2501.710 ;
        RECT 2032.380 2501.390 2032.640 2501.710 ;
        RECT 1327.260 2500.000 1327.400 2501.390 ;
        RECT 1327.190 2496.000 1327.470 2500.000 ;
        RECT 2032.440 2201.150 2032.580 2501.390 ;
        RECT 2032.380 2200.830 2032.640 2201.150 ;
        RECT 2900.860 2200.830 2901.120 2201.150 ;
        RECT 2900.920 2199.645 2901.060 2200.830 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 2198.860 2924.800 2200.060 ;
=======
        RECT 2898.065 2199.610 2898.395 2199.625 ;
=======
        RECT 2900.825 2199.610 2901.155 2199.625 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1883.770 201.860 1884.090 201.920 ;
        RECT 1897.570 201.860 1897.890 201.920 ;
        RECT 1883.770 201.720 1897.890 201.860 ;
        RECT 1883.770 201.660 1884.090 201.720 ;
        RECT 1897.570 201.660 1897.890 201.720 ;
        RECT 1242.070 201.520 1242.390 201.580 ;
        RECT 1249.890 201.520 1250.210 201.580 ;
        RECT 1242.070 201.380 1250.210 201.520 ;
        RECT 1242.070 201.320 1242.390 201.380 ;
        RECT 1249.890 201.320 1250.210 201.380 ;
        RECT 1799.130 201.180 1799.450 201.240 ;
        RECT 1805.570 201.180 1805.890 201.240 ;
        RECT 1799.130 201.040 1805.890 201.180 ;
        RECT 1799.130 200.980 1799.450 201.040 ;
        RECT 1805.570 200.980 1805.890 201.040 ;
        RECT 1944.950 200.840 1945.270 200.900 ;
        RECT 1955.990 200.840 1956.310 200.900 ;
        RECT 1944.950 200.700 1956.310 200.840 ;
        RECT 1944.950 200.640 1945.270 200.700 ;
        RECT 1955.990 200.640 1956.310 200.700 ;
        RECT 2456.470 200.840 2456.790 200.900 ;
        RECT 2504.310 200.840 2504.630 200.900 ;
        RECT 2456.470 200.700 2504.630 200.840 ;
        RECT 2456.470 200.640 2456.790 200.700 ;
        RECT 2504.310 200.640 2504.630 200.700 ;
        RECT 2621.610 200.840 2621.930 200.900 ;
        RECT 2622.530 200.840 2622.850 200.900 ;
        RECT 2621.610 200.700 2622.850 200.840 ;
        RECT 2621.610 200.640 2621.930 200.700 ;
        RECT 2622.530 200.640 2622.850 200.700 ;
        RECT 1642.270 200.500 1642.590 200.560 ;
        RECT 1690.110 200.500 1690.430 200.560 ;
        RECT 1642.270 200.360 1690.430 200.500 ;
        RECT 1642.270 200.300 1642.590 200.360 ;
        RECT 1690.110 200.300 1690.430 200.360 ;
        RECT 2070.070 200.500 2070.390 200.560 ;
        RECT 2117.910 200.500 2118.230 200.560 ;
        RECT 2070.070 200.360 2118.230 200.500 ;
        RECT 2070.070 200.300 2070.390 200.360 ;
        RECT 2117.910 200.300 2118.230 200.360 ;
        RECT 2649.670 200.500 2649.990 200.560 ;
        RECT 2697.510 200.500 2697.830 200.560 ;
        RECT 2649.670 200.360 2697.830 200.500 ;
        RECT 2649.670 200.300 2649.990 200.360 ;
        RECT 2697.510 200.300 2697.830 200.360 ;
      LAYER via ;
        RECT 1883.800 201.660 1884.060 201.920 ;
        RECT 1897.600 201.660 1897.860 201.920 ;
        RECT 1242.100 201.320 1242.360 201.580 ;
        RECT 1249.920 201.320 1250.180 201.580 ;
        RECT 1799.160 200.980 1799.420 201.240 ;
        RECT 1805.600 200.980 1805.860 201.240 ;
        RECT 1944.980 200.640 1945.240 200.900 ;
        RECT 1956.020 200.640 1956.280 200.900 ;
        RECT 2456.500 200.640 2456.760 200.900 ;
        RECT 2504.340 200.640 2504.600 200.900 ;
        RECT 2621.640 200.640 2621.900 200.900 ;
        RECT 2622.560 200.640 2622.820 200.900 ;
        RECT 1642.300 200.300 1642.560 200.560 ;
        RECT 1690.140 200.300 1690.400 200.560 ;
        RECT 2070.100 200.300 2070.360 200.560 ;
        RECT 2117.940 200.300 2118.200 200.560 ;
        RECT 2649.700 200.300 2649.960 200.560 ;
        RECT 2697.540 200.300 2697.800 200.560 ;
      LAYER met2 ;
        RECT 1159.750 2498.050 1160.030 2500.000 ;
        RECT 1161.590 2498.050 1161.870 2498.165 ;
        RECT 1159.750 2497.910 1161.870 2498.050 ;
        RECT 1159.750 2496.000 1160.030 2497.910 ;
        RECT 1161.590 2497.795 1161.870 2497.910 ;
        RECT 1883.800 201.805 1884.060 201.950 ;
        RECT 1897.600 201.805 1897.860 201.950 ;
        RECT 1242.090 201.435 1242.370 201.805 ;
        RECT 1242.100 201.290 1242.360 201.435 ;
        RECT 1249.920 201.290 1250.180 201.610 ;
        RECT 1524.530 201.435 1524.810 201.805 ;
        RECT 1690.130 201.435 1690.410 201.805 ;
        RECT 1883.790 201.435 1884.070 201.805 ;
        RECT 1897.590 201.435 1897.870 201.805 ;
        RECT 2117.930 201.435 2118.210 201.805 ;
        RECT 2234.310 201.690 2234.590 201.805 ;
        RECT 2235.230 201.690 2235.510 201.805 ;
        RECT 2234.310 201.550 2235.510 201.690 ;
        RECT 2234.310 201.435 2234.590 201.550 ;
        RECT 2235.230 201.435 2235.510 201.550 ;
        RECT 2304.230 201.435 2304.510 201.805 ;
        RECT 2427.510 201.690 2427.790 201.805 ;
        RECT 2428.430 201.690 2428.710 201.805 ;
        RECT 2427.510 201.550 2428.710 201.690 ;
        RECT 2427.510 201.435 2427.790 201.550 ;
        RECT 2428.430 201.435 2428.710 201.550 ;
        RECT 2573.330 201.435 2573.610 201.805 ;
        RECT 2697.530 201.435 2697.810 201.805 ;
        RECT 1249.980 200.445 1250.120 201.290 ;
        RECT 1379.630 200.755 1379.910 201.125 ;
        RECT 1427.930 200.755 1428.210 201.125 ;
        RECT 1476.230 200.755 1476.510 201.125 ;
        RECT 1249.910 200.075 1250.190 200.445 ;
        RECT 1379.700 197.725 1379.840 200.755 ;
        RECT 1428.000 199.765 1428.140 200.755 ;
        RECT 1427.930 199.395 1428.210 199.765 ;
        RECT 1476.300 199.085 1476.440 200.755 ;
        RECT 1476.230 198.715 1476.510 199.085 ;
        RECT 1524.600 197.725 1524.740 201.435 ;
        RECT 1606.410 200.755 1606.690 201.125 ;
        RECT 1606.480 199.085 1606.620 200.755 ;
        RECT 1690.200 200.590 1690.340 201.435 ;
        RECT 1799.160 201.125 1799.420 201.270 ;
        RECT 1805.600 201.125 1805.860 201.270 ;
        RECT 1799.150 200.755 1799.430 201.125 ;
        RECT 1805.590 200.755 1805.870 201.125 ;
        RECT 1944.970 200.755 1945.250 201.125 ;
        RECT 1944.980 200.610 1945.240 200.755 ;
        RECT 1956.020 200.610 1956.280 200.930 ;
        RECT 1642.300 200.445 1642.560 200.590 ;
        RECT 1642.290 200.075 1642.570 200.445 ;
        RECT 1690.140 200.270 1690.400 200.590 ;
        RECT 1956.080 200.445 1956.220 200.610 ;
        RECT 2118.000 200.590 2118.140 201.435 ;
        RECT 2070.100 200.445 2070.360 200.590 ;
        RECT 1956.010 200.075 1956.290 200.445 ;
        RECT 2004.310 200.075 2004.590 200.445 ;
        RECT 2051.230 200.330 2051.510 200.445 ;
        RECT 2052.150 200.330 2052.430 200.445 ;
        RECT 2051.230 200.190 2052.430 200.330 ;
        RECT 2051.230 200.075 2051.510 200.190 ;
        RECT 2052.150 200.075 2052.430 200.190 ;
        RECT 2070.090 200.075 2070.370 200.445 ;
        RECT 2117.940 200.270 2118.200 200.590 ;
        RECT 2004.380 199.085 2004.520 200.075 ;
        RECT 2304.300 199.765 2304.440 201.435 ;
        RECT 2456.490 200.755 2456.770 201.125 ;
        RECT 2573.400 201.010 2573.540 201.435 ;
        RECT 2574.250 201.010 2574.530 201.125 ;
        RECT 2456.500 200.610 2456.760 200.755 ;
        RECT 2504.340 200.610 2504.600 200.930 ;
        RECT 2573.400 200.870 2574.530 201.010 ;
        RECT 2574.250 200.755 2574.530 200.870 ;
        RECT 2621.630 200.755 2621.910 201.125 ;
        RECT 2621.640 200.610 2621.900 200.755 ;
        RECT 2622.560 200.610 2622.820 200.930 ;
        RECT 2504.400 200.445 2504.540 200.610 ;
        RECT 2622.620 200.445 2622.760 200.610 ;
        RECT 2697.600 200.590 2697.740 201.435 ;
        RECT 2649.700 200.445 2649.960 200.590 ;
        RECT 2504.330 200.075 2504.610 200.445 ;
        RECT 2622.550 200.075 2622.830 200.445 ;
        RECT 2649.690 200.075 2649.970 200.445 ;
        RECT 2697.540 200.270 2697.800 200.590 ;
        RECT 2304.230 199.395 2304.510 199.765 ;
        RECT 1606.410 198.715 1606.690 199.085 ;
        RECT 2004.310 198.715 2004.590 199.085 ;
        RECT 1379.630 197.355 1379.910 197.725 ;
        RECT 1524.530 197.355 1524.810 197.725 ;
      LAYER via2 ;
        RECT 1161.590 2497.840 1161.870 2498.120 ;
        RECT 1242.090 201.480 1242.370 201.760 ;
        RECT 1524.530 201.480 1524.810 201.760 ;
        RECT 1690.130 201.480 1690.410 201.760 ;
        RECT 1883.790 201.480 1884.070 201.760 ;
        RECT 1897.590 201.480 1897.870 201.760 ;
        RECT 2117.930 201.480 2118.210 201.760 ;
        RECT 2234.310 201.480 2234.590 201.760 ;
        RECT 2235.230 201.480 2235.510 201.760 ;
        RECT 2304.230 201.480 2304.510 201.760 ;
        RECT 2427.510 201.480 2427.790 201.760 ;
        RECT 2428.430 201.480 2428.710 201.760 ;
        RECT 2573.330 201.480 2573.610 201.760 ;
        RECT 2697.530 201.480 2697.810 201.760 ;
        RECT 1379.630 200.800 1379.910 201.080 ;
        RECT 1427.930 200.800 1428.210 201.080 ;
        RECT 1476.230 200.800 1476.510 201.080 ;
        RECT 1249.910 200.120 1250.190 200.400 ;
        RECT 1427.930 199.440 1428.210 199.720 ;
        RECT 1476.230 198.760 1476.510 199.040 ;
        RECT 1606.410 200.800 1606.690 201.080 ;
        RECT 1799.150 200.800 1799.430 201.080 ;
        RECT 1805.590 200.800 1805.870 201.080 ;
        RECT 1944.970 200.800 1945.250 201.080 ;
        RECT 1642.290 200.120 1642.570 200.400 ;
        RECT 1956.010 200.120 1956.290 200.400 ;
        RECT 2004.310 200.120 2004.590 200.400 ;
        RECT 2051.230 200.120 2051.510 200.400 ;
        RECT 2052.150 200.120 2052.430 200.400 ;
        RECT 2070.090 200.120 2070.370 200.400 ;
        RECT 2456.490 200.800 2456.770 201.080 ;
        RECT 2574.250 200.800 2574.530 201.080 ;
        RECT 2621.630 200.800 2621.910 201.080 ;
        RECT 2504.330 200.120 2504.610 200.400 ;
        RECT 2622.550 200.120 2622.830 200.400 ;
        RECT 2649.690 200.120 2649.970 200.400 ;
        RECT 2304.230 199.440 2304.510 199.720 ;
        RECT 1606.410 198.760 1606.690 199.040 ;
        RECT 2004.310 198.760 2004.590 199.040 ;
        RECT 1379.630 197.400 1379.910 197.680 ;
        RECT 1524.530 197.400 1524.810 197.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 204.420 2924.800 205.620 ;
=======
        RECT 1161.565 2498.130 1161.895 2498.145 ;
        RECT 1164.990 2498.130 1165.370 2498.140 ;
        RECT 1161.565 2497.830 1165.370 2498.130 ;
        RECT 1161.565 2497.815 1161.895 2497.830 ;
        RECT 1164.990 2497.820 1165.370 2497.830 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2916.710 204.870 2924.800 205.170 ;
        RECT 1242.065 201.770 1242.395 201.785 ;
        RECT 1224.830 201.470 1242.395 201.770 ;
        RECT 1224.830 201.090 1225.130 201.470 ;
        RECT 1242.065 201.455 1242.395 201.470 ;
        RECT 1524.505 201.770 1524.835 201.785 ;
        RECT 1690.105 201.770 1690.435 201.785 ;
        RECT 1883.765 201.770 1884.095 201.785 ;
        RECT 1524.505 201.470 1559.090 201.770 ;
        RECT 1524.505 201.455 1524.835 201.470 ;
        RECT 1199.990 200.790 1225.130 201.090 ;
        RECT 1379.605 201.090 1379.935 201.105 ;
        RECT 1427.905 201.090 1428.235 201.105 ;
        RECT 1476.205 201.090 1476.535 201.105 ;
        RECT 1379.605 200.790 1380.610 201.090 ;
        RECT 1164.990 200.410 1165.370 200.420 ;
        RECT 1199.990 200.410 1200.290 200.790 ;
        RECT 1379.605 200.775 1379.935 200.790 ;
        RECT 1164.990 200.110 1200.290 200.410 ;
        RECT 1249.885 200.410 1250.215 200.425 ;
        RECT 1290.110 200.410 1290.490 200.420 ;
        RECT 1249.885 200.110 1290.490 200.410 ;
        RECT 1164.990 200.100 1165.370 200.110 ;
        RECT 1249.885 200.095 1250.215 200.110 ;
        RECT 1290.110 200.100 1290.490 200.110 ;
        RECT 1380.310 199.730 1380.610 200.790 ;
        RECT 1427.905 200.790 1476.535 201.090 ;
        RECT 1427.905 200.775 1428.235 200.790 ;
        RECT 1476.205 200.775 1476.535 200.790 ;
        RECT 1558.790 200.410 1559.090 201.470 ;
        RECT 1690.105 201.470 1704.450 201.770 ;
        RECT 1690.105 201.455 1690.435 201.470 ;
        RECT 1606.385 201.090 1606.715 201.105 ;
        RECT 1559.710 200.790 1606.715 201.090 ;
        RECT 1559.710 200.410 1560.010 200.790 ;
        RECT 1606.385 200.775 1606.715 200.790 ;
        RECT 1642.265 200.410 1642.595 200.425 ;
        RECT 1558.790 200.110 1560.010 200.410 ;
        RECT 1641.590 200.110 1642.595 200.410 ;
        RECT 1704.150 200.410 1704.450 201.470 ;
        RECT 1849.510 201.470 1884.095 201.770 ;
        RECT 1799.125 201.090 1799.455 201.105 ;
        RECT 1752.910 200.790 1799.455 201.090 ;
        RECT 1752.910 200.410 1753.210 200.790 ;
        RECT 1799.125 200.775 1799.455 200.790 ;
        RECT 1805.565 201.090 1805.895 201.105 ;
        RECT 1805.565 200.790 1835.090 201.090 ;
        RECT 1805.565 200.775 1805.895 200.790 ;
        RECT 1704.150 200.110 1753.210 200.410 ;
        RECT 1834.790 200.410 1835.090 200.790 ;
        RECT 1849.510 200.410 1849.810 201.470 ;
        RECT 1883.765 201.455 1884.095 201.470 ;
        RECT 1897.565 201.770 1897.895 201.785 ;
        RECT 2117.905 201.770 2118.235 201.785 ;
        RECT 2234.285 201.770 2234.615 201.785 ;
        RECT 1897.565 201.470 1931.690 201.770 ;
        RECT 1897.565 201.455 1897.895 201.470 ;
        RECT 1931.390 201.090 1931.690 201.470 ;
        RECT 2117.905 201.470 2234.615 201.770 ;
        RECT 2117.905 201.455 2118.235 201.470 ;
        RECT 2234.285 201.455 2234.615 201.470 ;
        RECT 2235.205 201.770 2235.535 201.785 ;
        RECT 2304.205 201.770 2304.535 201.785 ;
        RECT 2427.485 201.770 2427.815 201.785 ;
        RECT 2235.205 201.470 2246.330 201.770 ;
        RECT 2235.205 201.455 2235.535 201.470 ;
        RECT 1944.945 201.090 1945.275 201.105 ;
        RECT 1931.390 200.790 1945.275 201.090 ;
        RECT 2246.030 201.090 2246.330 201.470 ;
        RECT 2304.205 201.470 2427.815 201.770 ;
        RECT 2304.205 201.455 2304.535 201.470 ;
        RECT 2427.485 201.455 2427.815 201.470 ;
        RECT 2428.405 201.770 2428.735 201.785 ;
        RECT 2573.305 201.770 2573.635 201.785 ;
        RECT 2428.405 201.470 2456.090 201.770 ;
        RECT 2428.405 201.455 2428.735 201.470 ;
        RECT 2269.910 201.090 2270.290 201.100 ;
        RECT 2246.030 200.790 2270.290 201.090 ;
        RECT 2455.790 201.090 2456.090 201.470 ;
        RECT 2525.710 201.470 2573.635 201.770 ;
        RECT 2456.465 201.090 2456.795 201.105 ;
        RECT 2455.790 200.790 2456.795 201.090 ;
        RECT 1944.945 200.775 1945.275 200.790 ;
        RECT 2269.910 200.780 2270.290 200.790 ;
        RECT 2456.465 200.775 2456.795 200.790 ;
        RECT 1834.790 200.110 1849.810 200.410 ;
        RECT 1955.985 200.410 1956.315 200.425 ;
        RECT 1980.110 200.410 1980.490 200.420 ;
        RECT 1955.985 200.110 1980.490 200.410 ;
        RECT 1427.905 199.730 1428.235 199.745 ;
        RECT 1380.310 199.430 1428.235 199.730 ;
        RECT 1427.905 199.415 1428.235 199.430 ;
        RECT 1290.110 199.050 1290.490 199.060 ;
        RECT 1331.510 199.050 1331.890 199.060 ;
        RECT 1290.110 198.750 1331.890 199.050 ;
        RECT 1290.110 198.740 1290.490 198.750 ;
        RECT 1331.510 198.740 1331.890 198.750 ;
        RECT 1476.205 199.050 1476.535 199.065 ;
        RECT 1606.385 199.050 1606.715 199.065 ;
        RECT 1641.590 199.050 1641.890 200.110 ;
        RECT 1642.265 200.095 1642.595 200.110 ;
        RECT 1955.985 200.095 1956.315 200.110 ;
        RECT 1980.110 200.100 1980.490 200.110 ;
        RECT 2004.285 200.410 2004.615 200.425 ;
        RECT 2051.205 200.410 2051.535 200.425 ;
        RECT 2004.285 200.110 2051.535 200.410 ;
        RECT 2004.285 200.095 2004.615 200.110 ;
        RECT 2051.205 200.095 2051.535 200.110 ;
        RECT 2052.125 200.410 2052.455 200.425 ;
        RECT 2070.065 200.410 2070.395 200.425 ;
        RECT 2052.125 200.110 2070.395 200.410 ;
        RECT 2052.125 200.095 2052.455 200.110 ;
        RECT 2070.065 200.095 2070.395 200.110 ;
        RECT 2504.305 200.410 2504.635 200.425 ;
        RECT 2525.710 200.410 2526.010 201.470 ;
        RECT 2573.305 201.455 2573.635 201.470 ;
        RECT 2697.505 201.770 2697.835 201.785 ;
        RECT 2697.505 201.470 2739.450 201.770 ;
        RECT 2697.505 201.455 2697.835 201.470 ;
        RECT 2574.225 201.090 2574.555 201.105 ;
        RECT 2621.605 201.090 2621.935 201.105 ;
        RECT 2574.225 200.790 2621.935 201.090 ;
        RECT 2739.150 201.090 2739.450 201.470 ;
        RECT 2787.910 201.470 2836.050 201.770 ;
        RECT 2739.150 200.790 2787.290 201.090 ;
        RECT 2574.225 200.775 2574.555 200.790 ;
        RECT 2621.605 200.775 2621.935 200.790 ;
        RECT 2504.305 200.110 2526.010 200.410 ;
        RECT 2622.525 200.410 2622.855 200.425 ;
        RECT 2649.665 200.410 2649.995 200.425 ;
        RECT 2622.525 200.110 2649.995 200.410 ;
        RECT 2786.990 200.410 2787.290 200.790 ;
        RECT 2787.910 200.410 2788.210 201.470 ;
        RECT 2835.750 201.090 2836.050 201.470 ;
        RECT 2916.710 201.090 2917.010 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2835.750 200.790 2883.890 201.090 ;
        RECT 2786.990 200.110 2788.210 200.410 ;
        RECT 2883.590 200.410 2883.890 200.790 ;
        RECT 2884.510 200.790 2917.010 201.090 ;
        RECT 2884.510 200.410 2884.810 200.790 ;
        RECT 2883.590 200.110 2884.810 200.410 ;
        RECT 2504.305 200.095 2504.635 200.110 ;
        RECT 2622.525 200.095 2622.855 200.110 ;
        RECT 2649.665 200.095 2649.995 200.110 ;
        RECT 2269.910 199.730 2270.290 199.740 ;
        RECT 2304.205 199.730 2304.535 199.745 ;
        RECT 2269.910 199.430 2304.535 199.730 ;
        RECT 2269.910 199.420 2270.290 199.430 ;
        RECT 2304.205 199.415 2304.535 199.430 ;
        RECT 1476.205 198.750 1477.210 199.050 ;
        RECT 1476.205 198.735 1476.535 198.750 ;
        RECT 1331.510 197.690 1331.890 197.700 ;
        RECT 1379.605 197.690 1379.935 197.705 ;
        RECT 1331.510 197.390 1379.935 197.690 ;
        RECT 1476.910 197.690 1477.210 198.750 ;
        RECT 1606.385 198.750 1641.890 199.050 ;
        RECT 1980.110 199.050 1980.490 199.060 ;
        RECT 2004.285 199.050 2004.615 199.065 ;
        RECT 1980.110 198.750 2004.615 199.050 ;
        RECT 1606.385 198.735 1606.715 198.750 ;
        RECT 1980.110 198.740 1980.490 198.750 ;
        RECT 2004.285 198.735 2004.615 198.750 ;
        RECT 1524.505 197.690 1524.835 197.705 ;
        RECT 1476.910 197.390 1524.835 197.690 ;
        RECT 1331.510 197.380 1331.890 197.390 ;
        RECT 1379.605 197.375 1379.935 197.390 ;
        RECT 1524.505 197.375 1524.835 197.390 ;
      LAYER via3 ;
        RECT 1165.020 2497.820 1165.340 2498.140 ;
        RECT 1165.020 200.100 1165.340 200.420 ;
        RECT 1290.140 200.100 1290.460 200.420 ;
        RECT 2269.940 200.780 2270.260 201.100 ;
        RECT 1290.140 198.740 1290.460 199.060 ;
        RECT 1331.540 198.740 1331.860 199.060 ;
        RECT 1980.140 200.100 1980.460 200.420 ;
        RECT 2269.940 199.420 2270.260 199.740 ;
        RECT 1331.540 197.380 1331.860 197.700 ;
        RECT 1980.140 198.740 1980.460 199.060 ;
      LAYER met4 ;
        RECT 1165.015 2497.815 1165.345 2498.145 ;
<<<<<<< HEAD
        RECT 1165.030 218.105 1165.330 2497.815 ;
        RECT 1165.015 217.775 1165.345 218.105 ;
        RECT 1980.135 202.815 1980.465 203.145 ;
        RECT 1980.150 201.785 1980.450 202.815 ;
        RECT 1248.735 201.455 1249.065 201.785 ;
        RECT 1980.135 201.455 1980.465 201.785 ;
        RECT 1248.750 200.425 1249.050 201.455 ;
        RECT 1248.735 200.095 1249.065 200.425 ;
        RECT 1345.335 200.095 1345.665 200.425 ;
        RECT 1345.350 199.065 1345.650 200.095 ;
        RECT 1345.335 198.735 1345.665 199.065 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1165.030 200.425 1165.330 2497.815 ;
        RECT 2269.935 200.775 2270.265 201.105 ;
        RECT 1165.015 200.095 1165.345 200.425 ;
        RECT 1290.135 200.095 1290.465 200.425 ;
        RECT 1980.135 200.095 1980.465 200.425 ;
        RECT 1290.150 199.065 1290.450 200.095 ;
        RECT 1980.150 199.065 1980.450 200.095 ;
        RECT 2269.950 199.745 2270.250 200.775 ;
        RECT 2269.935 199.415 2270.265 199.745 ;
        RECT 1290.135 198.735 1290.465 199.065 ;
        RECT 1331.535 198.735 1331.865 199.065 ;
        RECT 1980.135 198.735 1980.465 199.065 ;
        RECT 1331.550 197.705 1331.850 198.735 ;
        RECT 1331.535 197.375 1331.865 197.705 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1352.470 2546.840 1352.790 2546.900 ;
        RECT 2899.450 2546.840 2899.770 2546.900 ;
        RECT 1352.470 2546.700 2899.770 2546.840 ;
        RECT 1352.470 2546.640 1352.790 2546.700 ;
        RECT 2899.450 2546.640 2899.770 2546.700 ;
      LAYER via ;
        RECT 1352.500 2546.640 1352.760 2546.900 ;
        RECT 2899.480 2546.640 2899.740 2546.900 ;
      LAYER met2 ;
        RECT 2899.470 2551.515 2899.750 2551.885 ;
        RECT 2899.540 2546.930 2899.680 2551.515 ;
        RECT 1352.500 2546.610 1352.760 2546.930 ;
        RECT 2899.480 2546.610 2899.740 2546.930 ;
        RECT 1352.560 2499.410 1352.700 2546.610 ;
        RECT 1352.950 2499.410 1353.230 2500.000 ;
        RECT 1352.560 2499.270 1353.230 2499.410 ;
        RECT 1352.950 2496.000 1353.230 2499.270 ;
      LAYER via2 ;
        RECT 2899.470 2551.560 2899.750 2551.840 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 2551.100 2924.800 2552.300 ;
=======
        RECT 2900.825 2551.850 2901.155 2551.865 ;
=======
        RECT 2899.445 2551.850 2899.775 2551.865 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2899.445 2551.550 2924.800 2551.850 ;
        RECT 2899.445 2551.535 2899.775 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1372.710 2781.100 1373.030 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 1372.710 2780.960 2901.150 2781.100 ;
        RECT 1372.710 2780.900 1373.030 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 1372.740 2780.900 1373.000 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 1372.740 2780.870 1373.000 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 1372.270 2499.410 1372.550 2500.000 ;
        RECT 1372.800 2499.410 1372.940 2780.870 ;
        RECT 1372.270 2499.270 1372.940 2499.410 ;
        RECT 1372.270 2496.000 1372.550 2499.270 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2785.700 2924.800 2786.900 ;
=======
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1393.410 3015.700 1393.730 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 1393.410 3015.560 2901.150 3015.700 ;
        RECT 1393.410 3015.500 1393.730 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 1393.440 3015.500 1393.700 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 1393.440 3015.470 1393.700 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 1391.590 2499.410 1391.870 2500.000 ;
        RECT 1393.500 2499.410 1393.640 3015.470 ;
        RECT 1391.590 2499.270 1393.640 2499.410 ;
        RECT 1391.590 2496.000 1391.870 2499.270 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3020.300 2924.800 3021.500 ;
=======
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1414.110 3250.300 1414.430 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1414.110 3250.160 2901.150 3250.300 ;
        RECT 1414.110 3250.100 1414.430 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 1414.140 3250.100 1414.400 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1414.140 3250.070 1414.400 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1410.910 2498.730 1411.190 2500.000 ;
        RECT 1414.200 2498.730 1414.340 3250.070 ;
        RECT 1410.910 2498.590 1414.340 2498.730 ;
        RECT 1410.910 2496.000 1411.190 2498.590 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3254.900 2924.800 3256.100 ;
=======
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1434.810 3484.900 1435.130 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1434.810 3484.760 2901.150 3484.900 ;
        RECT 1434.810 3484.700 1435.130 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 1430.670 2515.900 1430.990 2515.960 ;
        RECT 1434.810 2515.900 1435.130 2515.960 ;
        RECT 1430.670 2515.760 1435.130 2515.900 ;
        RECT 1430.670 2515.700 1430.990 2515.760 ;
        RECT 1434.810 2515.700 1435.130 2515.760 ;
      LAYER via ;
        RECT 1434.840 3484.700 1435.100 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 1430.700 2515.700 1430.960 2515.960 ;
        RECT 1434.840 2515.700 1435.100 2515.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1434.840 3484.670 1435.100 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1434.900 2515.990 1435.040 3484.670 ;
        RECT 1430.700 2515.670 1430.960 2515.990 ;
        RECT 1434.840 2515.670 1435.100 2515.990 ;
        RECT 1430.760 2500.000 1430.900 2515.670 ;
        RECT 1430.690 2496.000 1430.970 2500.000 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3489.500 2924.800 3490.700 ;
=======
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1455.510 3502.920 1455.830 3502.980 ;
        RECT 2635.870 3502.920 2636.190 3502.980 ;
        RECT 1455.510 3502.780 2636.190 3502.920 ;
        RECT 1455.510 3502.720 1455.830 3502.780 ;
        RECT 2635.870 3502.720 2636.190 3502.780 ;
        RECT 1449.990 2515.900 1450.310 2515.960 ;
        RECT 1455.510 2515.900 1455.830 2515.960 ;
        RECT 1449.990 2515.760 1455.830 2515.900 ;
        RECT 1449.990 2515.700 1450.310 2515.760 ;
        RECT 1455.510 2515.700 1455.830 2515.760 ;
      LAYER via ;
        RECT 1455.540 3502.720 1455.800 3502.980 ;
        RECT 2635.900 3502.720 2636.160 3502.980 ;
        RECT 1450.020 2515.700 1450.280 2515.960 ;
        RECT 1455.540 2515.700 1455.800 2515.960 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2635.750 3519.700 2636.310 3524.800 ;
=======
        RECT 2635.750 3517.600 2636.310 3524.800 ;
<<<<<<< HEAD
        RECT 2635.960 3502.670 2636.100 3517.600 ;
        RECT 1462.440 3502.350 1462.700 3502.670 ;
        RECT 2635.900 3502.350 2636.160 3502.670 ;
        RECT 1462.500 2514.970 1462.640 3502.350 ;
        RECT 1457.380 2514.650 1457.640 2514.970 ;
        RECT 1462.440 2514.650 1462.700 2514.970 ;
        RECT 1457.440 2500.000 1457.580 2514.650 ;
        RECT 1457.370 2496.000 1457.650 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2635.960 3503.010 2636.100 3517.600 ;
        RECT 1455.540 3502.690 1455.800 3503.010 ;
        RECT 2635.900 3502.690 2636.160 3503.010 ;
        RECT 1455.600 2515.990 1455.740 3502.690 ;
        RECT 1450.020 2515.670 1450.280 2515.990 ;
        RECT 1455.540 2515.670 1455.800 2515.990 ;
        RECT 1450.080 2500.000 1450.220 2515.670 ;
        RECT 1450.010 2496.000 1450.290 2500.000 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1504.345 3499.365 1504.515 3504.635 ;
      LAYER mcon ;
        RECT 1504.345 3504.465 1504.515 3504.635 ;
      LAYER met1 ;
        RECT 1504.285 3504.620 1504.575 3504.665 ;
        RECT 2311.570 3504.620 2311.890 3504.680 ;
        RECT 1504.285 3504.480 2311.890 3504.620 ;
        RECT 1504.285 3504.435 1504.575 3504.480 ;
        RECT 2311.570 3504.420 2311.890 3504.480 ;
        RECT 1469.310 3499.520 1469.630 3499.580 ;
        RECT 1504.285 3499.520 1504.575 3499.565 ;
        RECT 1469.310 3499.380 1504.575 3499.520 ;
        RECT 1469.310 3499.320 1469.630 3499.380 ;
        RECT 1504.285 3499.335 1504.575 3499.380 ;
      LAYER via ;
        RECT 2311.600 3504.420 2311.860 3504.680 ;
        RECT 1469.340 3499.320 1469.600 3499.580 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2311.450 3519.700 2312.010 3524.800 ;
=======
        RECT 2311.450 3517.600 2312.010 3524.800 ;
<<<<<<< HEAD
        RECT 2311.660 3504.370 2311.800 3517.600 ;
        RECT 1483.140 3504.050 1483.400 3504.370 ;
        RECT 2311.600 3504.050 2311.860 3504.370 ;
        RECT 1483.200 2514.970 1483.340 3504.050 ;
        RECT 1477.160 2514.650 1477.420 2514.970 ;
        RECT 1483.140 2514.650 1483.400 2514.970 ;
        RECT 1477.220 2500.000 1477.360 2514.650 ;
        RECT 1477.150 2496.000 1477.430 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2311.660 3504.710 2311.800 3517.600 ;
        RECT 2311.600 3504.390 2311.860 3504.710 ;
        RECT 1469.340 3499.290 1469.600 3499.610 ;
        RECT 1469.400 2500.000 1469.540 3499.290 ;
        RECT 1469.330 2496.000 1469.610 2500.000 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1490.010 3500.200 1490.330 3500.260 ;
        RECT 1987.270 3500.200 1987.590 3500.260 ;
        RECT 1490.010 3500.060 1987.590 3500.200 ;
        RECT 1490.010 3500.000 1490.330 3500.060 ;
        RECT 1987.270 3500.000 1987.590 3500.060 ;
      LAYER via ;
        RECT 1490.040 3500.000 1490.300 3500.260 ;
        RECT 1987.300 3500.000 1987.560 3500.260 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1987.150 3519.700 1987.710 3524.800 ;
=======
        RECT 1987.150 3517.600 1987.710 3524.800 ;
<<<<<<< HEAD
        RECT 1987.360 3500.970 1987.500 3517.600 ;
        RECT 1496.940 3500.650 1497.200 3500.970 ;
        RECT 1987.300 3500.650 1987.560 3500.970 ;
        RECT 1497.000 2500.000 1497.140 3500.650 ;
        RECT 1496.930 2496.000 1497.210 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1987.360 3500.290 1987.500 3517.600 ;
        RECT 1490.040 3499.970 1490.300 3500.290 ;
        RECT 1987.300 3499.970 1987.560 3500.290 ;
        RECT 1488.650 2499.410 1488.930 2500.000 ;
        RECT 1490.100 2499.410 1490.240 3499.970 ;
        RECT 1488.650 2499.270 1490.240 2499.410 ;
        RECT 1488.650 2496.000 1488.930 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1586.685 3481.685 1586.855 3498.855 ;
        RECT 1635.445 3498.685 1635.615 3501.235 ;
      LAYER mcon ;
        RECT 1635.445 3501.065 1635.615 3501.235 ;
        RECT 1586.685 3498.685 1586.855 3498.855 ;
      LAYER met1 ;
        RECT 1635.385 3501.220 1635.675 3501.265 ;
        RECT 1662.510 3501.220 1662.830 3501.280 ;
        RECT 1635.385 3501.080 1662.830 3501.220 ;
        RECT 1635.385 3501.035 1635.675 3501.080 ;
        RECT 1662.510 3501.020 1662.830 3501.080 ;
        RECT 1586.625 3498.840 1586.915 3498.885 ;
        RECT 1635.385 3498.840 1635.675 3498.885 ;
        RECT 1586.625 3498.700 1635.675 3498.840 ;
        RECT 1586.625 3498.655 1586.915 3498.700 ;
        RECT 1635.385 3498.655 1635.675 3498.700 ;
        RECT 1510.710 3481.840 1511.030 3481.900 ;
        RECT 1586.625 3481.840 1586.915 3481.885 ;
        RECT 1510.710 3481.700 1586.915 3481.840 ;
        RECT 1510.710 3481.640 1511.030 3481.700 ;
        RECT 1586.625 3481.655 1586.915 3481.700 ;
      LAYER via ;
        RECT 1662.540 3501.020 1662.800 3501.280 ;
        RECT 1510.740 3481.640 1511.000 3481.900 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1662.390 3519.700 1662.950 3524.800 ;
=======
        RECT 1662.390 3517.600 1662.950 3524.800 ;
<<<<<<< HEAD
        RECT 1662.600 3498.930 1662.740 3517.600 ;
        RECT 1517.640 3498.610 1517.900 3498.930 ;
        RECT 1662.540 3498.610 1662.800 3498.930 ;
        RECT 1516.710 2499.410 1516.990 2500.000 ;
        RECT 1517.700 2499.410 1517.840 3498.610 ;
        RECT 1516.710 2499.270 1517.840 2499.410 ;
        RECT 1516.710 2496.000 1516.990 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1662.600 3501.310 1662.740 3517.600 ;
        RECT 1662.540 3500.990 1662.800 3501.310 ;
        RECT 1510.740 3481.610 1511.000 3481.930 ;
        RECT 1510.800 2500.090 1510.940 3481.610 ;
        RECT 1507.970 2499.410 1508.250 2500.000 ;
        RECT 1509.420 2499.950 1510.940 2500.090 ;
        RECT 1509.420 2499.410 1509.560 2499.950 ;
        RECT 1507.970 2499.270 1509.560 2499.410 ;
        RECT 1507.970 2496.000 1508.250 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3499.180 1338.530 3499.240 ;
        RECT 1524.970 3499.180 1525.290 3499.240 ;
        RECT 1338.210 3499.040 1525.290 3499.180 ;
        RECT 1338.210 3498.980 1338.530 3499.040 ;
        RECT 1524.970 3498.980 1525.290 3499.040 ;
      LAYER via ;
        RECT 1338.240 3498.980 1338.500 3499.240 ;
        RECT 1525.000 3498.980 1525.260 3499.240 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1338.090 3519.700 1338.650 3524.800 ;
=======
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3499.270 1338.440 3517.600 ;
        RECT 1338.240 3498.950 1338.500 3499.270 ;
<<<<<<< HEAD
        RECT 1528.220 3498.950 1528.480 3499.270 ;
        RECT 1528.280 2518.370 1528.420 3498.950 ;
        RECT 1528.220 2518.050 1528.480 2518.370 ;
        RECT 1534.660 2518.050 1534.920 2518.370 ;
        RECT 1534.720 2499.410 1534.860 2518.050 ;
        RECT 1536.490 2499.410 1536.770 2500.000 ;
        RECT 1534.720 2499.270 1536.770 2499.410 ;
        RECT 1536.490 2496.000 1536.770 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1525.000 3498.950 1525.260 3499.270 ;
        RECT 1525.060 2499.410 1525.200 3498.950 ;
        RECT 1527.290 2499.410 1527.570 2500.000 ;
        RECT 1525.060 2499.270 1527.570 2499.410 ;
        RECT 1527.290 2496.000 1527.570 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1179.050 2506.720 1179.370 2506.780 ;
        RECT 1976.690 2506.720 1977.010 2506.780 ;
        RECT 1179.050 2506.580 1977.010 2506.720 ;
        RECT 1179.050 2506.520 1179.370 2506.580 ;
        RECT 1976.690 2506.520 1977.010 2506.580 ;
        RECT 1976.690 441.560 1977.010 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 1976.690 441.420 2901.150 441.560 ;
        RECT 1976.690 441.360 1977.010 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 1179.080 2506.520 1179.340 2506.780 ;
        RECT 1976.720 2506.520 1976.980 2506.780 ;
        RECT 1976.720 441.360 1976.980 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 1179.080 2506.490 1179.340 2506.810 ;
        RECT 1976.720 2506.490 1976.980 2506.810 ;
        RECT 1179.140 2500.000 1179.280 2506.490 ;
        RECT 1179.070 2496.000 1179.350 2500.000 ;
        RECT 1976.780 441.650 1976.920 2506.490 ;
        RECT 1976.720 441.330 1976.980 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 439.020 2924.800 440.220 ;
=======
        RECT 1178.125 2498.140 1178.455 2498.145 ;
        RECT 1177.870 2498.130 1178.455 2498.140 ;
        RECT 1177.670 2497.830 1178.455 2498.130 ;
        RECT 1177.870 2497.820 1178.455 2497.830 ;
        RECT 1178.125 2497.815 1178.455 2497.820 ;
=======
        RECT 2900.825 439.770 2901.155 439.785 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
<<<<<<< HEAD
        RECT 2835.750 435.390 2883.890 435.690 ;
        RECT 2786.990 434.710 2788.210 435.010 ;
        RECT 2883.590 435.010 2883.890 435.390 ;
        RECT 2884.510 435.390 2917.010 435.690 ;
        RECT 2884.510 435.010 2884.810 435.390 ;
        RECT 2883.590 434.710 2884.810 435.010 ;
        RECT 2069.605 434.695 2069.935 434.710 ;
      LAYER via3 ;
        RECT 1177.900 2497.820 1178.220 2498.140 ;
        RECT 1177.900 436.740 1178.220 437.060 ;
        RECT 1738.180 436.060 1738.500 436.380 ;
        RECT 1834.780 436.060 1835.100 436.380 ;
        RECT 1738.180 434.700 1738.500 435.020 ;
        RECT 1834.780 434.700 1835.100 435.020 ;
      LAYER met4 ;
        RECT 1177.895 2497.815 1178.225 2498.145 ;
        RECT 1177.910 437.065 1178.210 2497.815 ;
        RECT 1177.895 436.735 1178.225 437.065 ;
        RECT 1738.175 436.055 1738.505 436.385 ;
        RECT 1834.775 436.055 1835.105 436.385 ;
        RECT 1738.190 435.025 1738.490 436.055 ;
        RECT 1834.790 435.025 1835.090 436.055 ;
        RECT 1738.175 434.695 1738.505 435.025 ;
        RECT 1834.775 434.695 1835.105 435.025 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3500.540 1014.230 3500.600 ;
        RECT 1545.670 3500.540 1545.990 3500.600 ;
        RECT 1013.910 3500.400 1545.990 3500.540 ;
        RECT 1013.910 3500.340 1014.230 3500.400 ;
        RECT 1545.670 3500.340 1545.990 3500.400 ;
      LAYER via ;
        RECT 1013.940 3500.340 1014.200 3500.600 ;
        RECT 1545.700 3500.340 1545.960 3500.600 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1013.790 3519.700 1014.350 3524.800 ;
=======
        RECT 1013.790 3517.600 1014.350 3524.800 ;
<<<<<<< HEAD
        RECT 1014.000 3501.310 1014.140 3517.600 ;
        RECT 1013.940 3500.990 1014.200 3501.310 ;
        RECT 1535.120 3500.990 1535.380 3501.310 ;
        RECT 1535.180 2518.370 1535.320 3500.990 ;
        RECT 1535.120 2518.050 1535.380 2518.370 ;
        RECT 1554.900 2518.050 1555.160 2518.370 ;
        RECT 1554.960 2499.410 1555.100 2518.050 ;
        RECT 1556.270 2499.410 1556.550 2500.000 ;
        RECT 1554.960 2499.270 1556.550 2499.410 ;
        RECT 1556.270 2496.000 1556.550 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1014.000 3500.630 1014.140 3517.600 ;
        RECT 1013.940 3500.310 1014.200 3500.630 ;
        RECT 1545.700 3500.310 1545.960 3500.630 ;
        RECT 1545.760 2499.410 1545.900 3500.310 ;
        RECT 1546.610 2499.410 1546.890 2500.000 ;
        RECT 1545.760 2499.270 1546.890 2499.410 ;
        RECT 1546.610 2496.000 1546.890 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 689.150 3504.280 689.470 3504.340 ;
        RECT 1559.470 3504.280 1559.790 3504.340 ;
        RECT 689.150 3504.140 1559.790 3504.280 ;
        RECT 689.150 3504.080 689.470 3504.140 ;
        RECT 1559.470 3504.080 1559.790 3504.140 ;
        RECT 1559.470 2511.140 1559.790 2511.200 ;
        RECT 1564.070 2511.140 1564.390 2511.200 ;
        RECT 1559.470 2511.000 1564.390 2511.140 ;
        RECT 1559.470 2510.940 1559.790 2511.000 ;
        RECT 1564.070 2510.940 1564.390 2511.000 ;
      LAYER via ;
        RECT 689.180 3504.080 689.440 3504.340 ;
        RECT 1559.500 3504.080 1559.760 3504.340 ;
        RECT 1559.500 2510.940 1559.760 2511.200 ;
        RECT 1564.100 2510.940 1564.360 2511.200 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 689.030 3519.700 689.590 3524.800 ;
=======
        RECT 689.030 3517.600 689.590 3524.800 ;
<<<<<<< HEAD
        RECT 689.240 3504.030 689.380 3517.600 ;
        RECT 689.180 3503.710 689.440 3504.030 ;
        RECT 1555.820 3503.710 1556.080 3504.030 ;
        RECT 1555.880 2518.370 1556.020 3503.710 ;
        RECT 1555.820 2518.050 1556.080 2518.370 ;
        RECT 1576.060 2517.710 1576.320 2518.030 ;
        RECT 1576.120 2500.000 1576.260 2517.710 ;
        RECT 1576.050 2496.000 1576.330 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 689.240 3504.370 689.380 3517.600 ;
        RECT 689.180 3504.050 689.440 3504.370 ;
        RECT 1559.500 3504.050 1559.760 3504.370 ;
        RECT 1559.560 2511.230 1559.700 3504.050 ;
        RECT 1559.500 2510.910 1559.760 2511.230 ;
        RECT 1564.100 2510.910 1564.360 2511.230 ;
        RECT 1564.160 2499.410 1564.300 2510.910 ;
        RECT 1565.930 2499.410 1566.210 2500.000 ;
        RECT 1564.160 2499.270 1566.210 2499.410 ;
        RECT 1565.930 2496.000 1566.210 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.580 365.170 3502.640 ;
        RECT 1580.630 3502.580 1580.950 3502.640 ;
        RECT 364.850 3502.440 1580.950 3502.580 ;
        RECT 364.850 3502.380 365.170 3502.440 ;
        RECT 1580.630 3502.380 1580.950 3502.440 ;
      LAYER via ;
        RECT 364.880 3502.380 365.140 3502.640 ;
        RECT 1580.660 3502.380 1580.920 3502.640 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 364.730 3519.700 365.290 3524.800 ;
=======
        RECT 364.730 3517.600 365.290 3524.800 ;
<<<<<<< HEAD
        RECT 364.940 3502.330 365.080 3517.600 ;
        RECT 364.880 3502.010 365.140 3502.330 ;
        RECT 1576.520 3502.010 1576.780 3502.330 ;
        RECT 1576.580 2518.030 1576.720 3502.010 ;
        RECT 1576.520 2517.710 1576.780 2518.030 ;
        RECT 1595.840 2517.710 1596.100 2518.030 ;
        RECT 1595.900 2500.000 1596.040 2517.710 ;
        RECT 1595.830 2496.000 1596.110 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 364.940 3502.670 365.080 3517.600 ;
        RECT 364.880 3502.350 365.140 3502.670 ;
        RECT 1580.660 3502.350 1580.920 3502.670 ;
        RECT 1580.720 2500.770 1580.860 3502.350 ;
        RECT 1580.720 2500.630 1583.160 2500.770 ;
        RECT 1583.020 2499.410 1583.160 2500.630 ;
        RECT 1585.250 2499.410 1585.530 2500.000 ;
        RECT 1583.020 2499.270 1585.530 2499.410 ;
        RECT 1585.250 2496.000 1585.530 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 40.430 3519.700 40.990 3524.800 ;
=======
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
        RECT 1600.890 3501.475 1601.170 3501.845 ;
        RECT 1600.960 2500.770 1601.100 3501.475 ;
        RECT 1600.960 2500.630 1602.480 2500.770 ;
        RECT 1602.340 2499.410 1602.480 2500.630 ;
        RECT 1604.570 2499.410 1604.850 2500.000 ;
        RECT 1602.340 2499.270 1604.850 2499.410 ;
        RECT 1604.570 2496.000 1604.850 2499.270 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
        RECT 1600.890 3501.520 1601.170 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 1600.865 3501.810 1601.195 3501.825 ;
        RECT 40.545 3501.510 1601.195 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
<<<<<<< HEAD
        RECT 1597.185 3501.495 1597.515 3501.510 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1600.865 3501.495 1601.195 3501.510 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 1621.570 3263.900 1621.890 3263.960 ;
        RECT 15.250 3263.760 1621.890 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 1621.570 3263.700 1621.890 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 1621.600 3263.700 1621.860 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 1621.600 3263.670 1621.860 3263.990 ;
        RECT 1621.660 2499.410 1621.800 3263.670 ;
        RECT 1623.890 2499.410 1624.170 2500.000 ;
        RECT 1621.660 2499.270 1624.170 2499.410 ;
        RECT 1623.890 2496.000 1624.170 2499.270 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3267.140 0.300 3268.340 ;
=======
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2974.220 17.870 2974.280 ;
        RECT 1642.270 2974.220 1642.590 2974.280 ;
        RECT 17.550 2974.080 1642.590 2974.220 ;
        RECT 17.550 2974.020 17.870 2974.080 ;
        RECT 1642.270 2974.020 1642.590 2974.080 ;
      LAYER via ;
        RECT 17.580 2974.020 17.840 2974.280 ;
        RECT 1642.300 2974.020 1642.560 2974.280 ;
      LAYER met2 ;
        RECT 17.570 2979.915 17.850 2980.285 ;
        RECT 17.640 2974.310 17.780 2979.915 ;
        RECT 17.580 2973.990 17.840 2974.310 ;
        RECT 1642.300 2973.990 1642.560 2974.310 ;
        RECT 1642.360 2499.410 1642.500 2973.990 ;
        RECT 1643.210 2499.410 1643.490 2500.000 ;
        RECT 1642.360 2499.270 1643.490 2499.410 ;
        RECT 1643.210 2496.000 1643.490 2499.270 ;
      LAYER via2 ;
        RECT 17.570 2979.960 17.850 2980.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2979.500 0.300 2980.700 ;
=======
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 17.545 2980.250 17.875 2980.265 ;
        RECT -4.800 2979.950 17.875 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
<<<<<<< HEAD
        RECT 16.165 2979.935 16.495 2979.950 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 17.545 2979.935 17.875 2979.950 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 2691.340 16.490 2691.400 ;
        RECT 1656.530 2691.340 1656.850 2691.400 ;
        RECT 16.170 2691.200 1656.850 2691.340 ;
        RECT 16.170 2691.140 16.490 2691.200 ;
        RECT 1656.530 2691.140 1656.850 2691.200 ;
      LAYER via ;
        RECT 16.200 2691.140 16.460 2691.400 ;
        RECT 1656.560 2691.140 1656.820 2691.400 ;
      LAYER met2 ;
        RECT 16.190 2692.955 16.470 2693.325 ;
        RECT 16.260 2691.430 16.400 2692.955 ;
        RECT 16.200 2691.110 16.460 2691.430 ;
        RECT 1656.560 2691.110 1656.820 2691.430 ;
        RECT 1656.620 2500.090 1656.760 2691.110 ;
        RECT 1656.620 2499.950 1660.900 2500.090 ;
        RECT 1660.760 2499.410 1660.900 2499.950 ;
        RECT 1662.530 2499.410 1662.810 2500.000 ;
        RECT 1660.760 2499.270 1662.810 2499.410 ;
        RECT 1662.530 2496.000 1662.810 2499.270 ;
      LAYER via2 ;
        RECT 16.190 2693.000 16.470 2693.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2692.540 0.300 2693.740 ;
=======
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 16.165 2693.290 16.495 2693.305 ;
        RECT -4.800 2692.990 16.495 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
<<<<<<< HEAD
        RECT 17.085 2692.975 17.415 2692.990 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.165 2692.975 16.495 2692.990 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1135.350 2502.640 1135.670 2502.700 ;
        RECT 1681.830 2502.640 1682.150 2502.700 ;
        RECT 1135.350 2502.500 1682.150 2502.640 ;
        RECT 1135.350 2502.440 1135.670 2502.500 ;
        RECT 1681.830 2502.440 1682.150 2502.500 ;
        RECT 16.170 2408.120 16.490 2408.180 ;
        RECT 1135.350 2408.120 1135.670 2408.180 ;
        RECT 16.170 2407.980 1135.670 2408.120 ;
        RECT 16.170 2407.920 16.490 2407.980 ;
        RECT 1135.350 2407.920 1135.670 2407.980 ;
      LAYER via ;
        RECT 1135.380 2502.440 1135.640 2502.700 ;
        RECT 1681.860 2502.440 1682.120 2502.700 ;
        RECT 16.200 2407.920 16.460 2408.180 ;
        RECT 1135.380 2407.920 1135.640 2408.180 ;
      LAYER met2 ;
        RECT 1135.380 2502.410 1135.640 2502.730 ;
        RECT 1681.860 2502.410 1682.120 2502.730 ;
        RECT 1135.440 2408.210 1135.580 2502.410 ;
        RECT 1681.920 2500.000 1682.060 2502.410 ;
        RECT 1681.850 2496.000 1682.130 2500.000 ;
        RECT 16.200 2407.890 16.460 2408.210 ;
        RECT 1135.380 2407.890 1135.640 2408.210 ;
        RECT 16.260 2405.685 16.400 2407.890 ;
        RECT 16.190 2405.315 16.470 2405.685 ;
      LAYER via2 ;
        RECT 16.190 2405.360 16.470 2405.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2404.900 0.300 2406.100 ;
=======
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 16.165 2405.650 16.495 2405.665 ;
        RECT -4.800 2405.350 16.495 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
<<<<<<< HEAD
        RECT 13.865 2405.335 14.195 2405.350 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.165 2405.335 16.495 2405.350 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1173.605 2495.855 1173.775 2496.195 ;
        RECT 1207.645 2496.025 1207.815 2496.875 ;
        RECT 1172.685 2495.685 1173.775 2495.855 ;
        RECT 1255.485 2495.685 1255.655 2496.875 ;
        RECT 1304.245 2496.025 1304.415 2497.215 ;
        RECT 1352.085 2495.685 1352.255 2497.215 ;
        RECT 1390.725 2495.345 1390.895 2496.535 ;
        RECT 1401.305 2495.515 1401.475 2497.215 ;
        RECT 1448.685 2495.685 1448.855 2497.215 ;
        RECT 1400.845 2495.345 1401.475 2495.515 ;
        RECT 1497.445 2495.345 1497.615 2496.195 ;
        RECT 1521.365 2495.345 1521.535 2496.195 ;
      LAYER mcon ;
        RECT 1304.245 2497.045 1304.415 2497.215 ;
        RECT 1207.645 2496.705 1207.815 2496.875 ;
        RECT 1173.605 2496.025 1173.775 2496.195 ;
        RECT 1255.485 2496.705 1255.655 2496.875 ;
        RECT 1352.085 2497.045 1352.255 2497.215 ;
        RECT 1401.305 2497.045 1401.475 2497.215 ;
        RECT 1390.725 2496.365 1390.895 2496.535 ;
        RECT 1448.685 2497.045 1448.855 2497.215 ;
        RECT 1497.445 2496.025 1497.615 2496.195 ;
        RECT 1521.365 2496.025 1521.535 2496.195 ;
      LAYER met1 ;
        RECT 1304.185 2497.200 1304.475 2497.245 ;
        RECT 1352.025 2497.200 1352.315 2497.245 ;
        RECT 1304.185 2497.060 1352.315 2497.200 ;
        RECT 1304.185 2497.015 1304.475 2497.060 ;
        RECT 1352.025 2497.015 1352.315 2497.060 ;
        RECT 1401.245 2497.200 1401.535 2497.245 ;
        RECT 1448.625 2497.200 1448.915 2497.245 ;
        RECT 1401.245 2497.060 1448.915 2497.200 ;
        RECT 1401.245 2497.015 1401.535 2497.060 ;
        RECT 1448.625 2497.015 1448.915 2497.060 ;
        RECT 1207.585 2496.860 1207.875 2496.905 ;
        RECT 1255.425 2496.860 1255.715 2496.905 ;
        RECT 1207.585 2496.720 1255.715 2496.860 ;
        RECT 1207.585 2496.675 1207.875 2496.720 ;
        RECT 1255.425 2496.675 1255.715 2496.720 ;
        RECT 1390.665 2496.520 1390.955 2496.565 ;
        RECT 1700.230 2496.520 1700.550 2496.580 ;
        RECT 1366.820 2496.380 1390.955 2496.520 ;
        RECT 1173.545 2496.180 1173.835 2496.225 ;
        RECT 1207.585 2496.180 1207.875 2496.225 ;
        RECT 1304.185 2496.180 1304.475 2496.225 ;
        RECT 1366.820 2496.180 1366.960 2496.380 ;
        RECT 1390.665 2496.335 1390.955 2496.380 ;
        RECT 1546.220 2496.380 1561.540 2496.520 ;
        RECT 1497.385 2496.180 1497.675 2496.225 ;
        RECT 1173.545 2496.040 1207.875 2496.180 ;
        RECT 1173.545 2495.995 1173.835 2496.040 ;
        RECT 1207.585 2495.995 1207.875 2496.040 ;
        RECT 1269.760 2496.040 1304.475 2496.180 ;
        RECT 1134.890 2495.840 1135.210 2495.900 ;
        RECT 1172.625 2495.840 1172.915 2495.885 ;
        RECT 1134.890 2495.700 1172.915 2495.840 ;
        RECT 1134.890 2495.640 1135.210 2495.700 ;
        RECT 1172.625 2495.655 1172.915 2495.700 ;
        RECT 1255.425 2495.840 1255.715 2495.885 ;
        RECT 1269.760 2495.840 1269.900 2496.040 ;
        RECT 1304.185 2495.995 1304.475 2496.040 ;
        RECT 1366.360 2496.040 1366.960 2496.180 ;
        RECT 1462.960 2496.040 1497.675 2496.180 ;
        RECT 1255.425 2495.700 1269.900 2495.840 ;
        RECT 1352.025 2495.840 1352.315 2495.885 ;
        RECT 1366.360 2495.840 1366.500 2496.040 ;
        RECT 1352.025 2495.700 1366.500 2495.840 ;
        RECT 1448.625 2495.840 1448.915 2495.885 ;
        RECT 1462.960 2495.840 1463.100 2496.040 ;
        RECT 1497.385 2495.995 1497.675 2496.040 ;
        RECT 1521.305 2496.180 1521.595 2496.225 ;
        RECT 1546.220 2496.180 1546.360 2496.380 ;
        RECT 1521.305 2496.040 1546.360 2496.180 ;
        RECT 1561.400 2496.180 1561.540 2496.380 ;
        RECT 1608.780 2496.380 1700.550 2496.520 ;
        RECT 1608.780 2496.180 1608.920 2496.380 ;
        RECT 1700.230 2496.320 1700.550 2496.380 ;
        RECT 1561.400 2496.040 1608.920 2496.180 ;
        RECT 1521.305 2495.995 1521.595 2496.040 ;
        RECT 1448.625 2495.700 1463.100 2495.840 ;
        RECT 1255.425 2495.655 1255.715 2495.700 ;
        RECT 1352.025 2495.655 1352.315 2495.700 ;
        RECT 1448.625 2495.655 1448.915 2495.700 ;
        RECT 1390.665 2495.500 1390.955 2495.545 ;
        RECT 1400.785 2495.500 1401.075 2495.545 ;
        RECT 1390.665 2495.360 1401.075 2495.500 ;
        RECT 1390.665 2495.315 1390.955 2495.360 ;
        RECT 1400.785 2495.315 1401.075 2495.360 ;
        RECT 1497.385 2495.500 1497.675 2495.545 ;
        RECT 1521.305 2495.500 1521.595 2495.545 ;
        RECT 1497.385 2495.360 1521.595 2495.500 ;
        RECT 1497.385 2495.315 1497.675 2495.360 ;
        RECT 1521.305 2495.315 1521.595 2495.360 ;
        RECT 16.630 2125.240 16.950 2125.300 ;
        RECT 1134.890 2125.240 1135.210 2125.300 ;
        RECT 16.630 2125.100 1135.210 2125.240 ;
        RECT 16.630 2125.040 16.950 2125.100 ;
        RECT 1134.890 2125.040 1135.210 2125.100 ;
      LAYER via ;
        RECT 1134.920 2495.640 1135.180 2495.900 ;
        RECT 1700.260 2496.320 1700.520 2496.580 ;
        RECT 16.660 2125.040 16.920 2125.300 ;
        RECT 1134.920 2125.040 1135.180 2125.300 ;
      LAYER met2 ;
        RECT 1701.630 2496.690 1701.910 2500.000 ;
        RECT 1700.320 2496.610 1701.910 2496.690 ;
        RECT 1700.260 2496.550 1701.910 2496.610 ;
        RECT 1700.260 2496.290 1700.520 2496.550 ;
        RECT 1701.630 2496.000 1701.910 2496.550 ;
        RECT 1134.920 2495.610 1135.180 2495.930 ;
        RECT 1134.980 2125.330 1135.120 2495.610 ;
        RECT 16.660 2125.010 16.920 2125.330 ;
        RECT 1134.920 2125.010 1135.180 2125.330 ;
        RECT 16.720 2118.725 16.860 2125.010 ;
        RECT 16.650 2118.355 16.930 2118.725 ;
      LAYER via2 ;
        RECT 16.650 2118.400 16.930 2118.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2117.940 0.300 2119.140 ;
=======
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.625 2118.690 16.955 2118.705 ;
        RECT -4.800 2118.390 16.955 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
<<<<<<< HEAD
        RECT 13.865 2118.375 14.195 2118.390 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 2118.375 16.955 2118.390 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1080.150 2509.780 1080.470 2509.840 ;
        RECT 1720.930 2509.780 1721.250 2509.840 ;
        RECT 1080.150 2509.640 1721.250 2509.780 ;
        RECT 1080.150 2509.580 1080.470 2509.640 ;
        RECT 1720.930 2509.580 1721.250 2509.640 ;
        RECT 15.710 1835.220 16.030 1835.280 ;
        RECT 1080.150 1835.220 1080.470 1835.280 ;
        RECT 15.710 1835.080 1080.470 1835.220 ;
        RECT 15.710 1835.020 16.030 1835.080 ;
        RECT 1080.150 1835.020 1080.470 1835.080 ;
      LAYER via ;
        RECT 1080.180 2509.580 1080.440 2509.840 ;
        RECT 1720.960 2509.580 1721.220 2509.840 ;
        RECT 15.740 1835.020 16.000 1835.280 ;
        RECT 1080.180 1835.020 1080.440 1835.280 ;
      LAYER met2 ;
        RECT 1080.180 2509.550 1080.440 2509.870 ;
        RECT 1720.960 2509.550 1721.220 2509.870 ;
        RECT 1080.240 1835.310 1080.380 2509.550 ;
        RECT 1721.020 2500.000 1721.160 2509.550 ;
        RECT 1720.950 2496.000 1721.230 2500.000 ;
        RECT 15.740 1834.990 16.000 1835.310 ;
        RECT 1080.180 1834.990 1080.440 1835.310 ;
        RECT 15.800 1831.085 15.940 1834.990 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1830.300 0.300 1831.500 ;
=======
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1200.210 2498.560 1200.530 2498.620 ;
        RECT 1997.390 2498.560 1997.710 2498.620 ;
        RECT 1200.210 2498.420 1997.710 2498.560 ;
        RECT 1200.210 2498.360 1200.530 2498.420 ;
        RECT 1997.390 2498.360 1997.710 2498.420 ;
        RECT 1997.390 676.160 1997.710 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 1997.390 676.020 2901.150 676.160 ;
        RECT 1997.390 675.960 1997.710 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 1200.240 2498.360 1200.500 2498.620 ;
        RECT 1997.420 2498.360 1997.680 2498.620 ;
        RECT 1997.420 675.960 1997.680 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 1198.390 2498.730 1198.670 2500.000 ;
        RECT 1198.390 2498.650 1200.440 2498.730 ;
        RECT 1198.390 2498.590 1200.500 2498.650 ;
        RECT 1198.390 2496.000 1198.670 2498.590 ;
        RECT 1200.240 2498.330 1200.500 2498.590 ;
        RECT 1997.420 2498.330 1997.680 2498.650 ;
        RECT 1997.480 676.250 1997.620 2498.330 ;
        RECT 1997.420 675.930 1997.680 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 673.620 2924.800 674.820 ;
=======
        RECT 1199.745 2498.140 1200.075 2498.145 ;
        RECT 1199.745 2498.130 1200.330 2498.140 ;
        RECT 1199.745 2497.830 1200.530 2498.130 ;
        RECT 1199.745 2497.820 1200.330 2497.830 ;
        RECT 1199.745 2497.815 1200.075 2497.820 ;
=======
        RECT 2900.825 674.370 2901.155 674.385 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
<<<<<<< HEAD
        RECT 2835.750 669.990 2883.890 670.290 ;
        RECT 2786.990 669.310 2788.210 669.610 ;
        RECT 2883.590 669.610 2883.890 669.990 ;
        RECT 2884.510 669.990 2917.010 670.290 ;
        RECT 2884.510 669.610 2884.810 669.990 ;
        RECT 2883.590 669.310 2884.810 669.610 ;
        RECT 2052.585 669.295 2052.915 669.310 ;
        RECT 1895.265 667.950 1931.690 668.250 ;
        RECT 1895.265 667.935 1895.595 667.950 ;
      LAYER via3 ;
        RECT 1199.980 2497.820 1200.300 2498.140 ;
        RECT 1980.140 672.020 1980.460 672.340 ;
        RECT 1199.980 670.660 1200.300 670.980 ;
        RECT 1980.140 670.660 1980.460 670.980 ;
      LAYER met4 ;
        RECT 1199.975 2497.815 1200.305 2498.145 ;
        RECT 1199.990 670.985 1200.290 2497.815 ;
        RECT 1980.135 672.015 1980.465 672.345 ;
        RECT 1980.150 670.985 1980.450 672.015 ;
        RECT 1199.975 670.655 1200.305 670.985 ;
        RECT 1980.135 670.655 1980.465 670.985 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1400.845 2497.385 1401.935 2497.555 ;
        RECT 1197.065 2494.325 1197.235 2495.515 ;
        RECT 1245.365 2494.325 1245.535 2495.515 ;
        RECT 1292.285 2495.345 1292.455 2496.875 ;
        RECT 1341.965 2495.345 1342.135 2496.875 ;
        RECT 1390.265 2495.345 1390.435 2496.875 ;
        RECT 1400.845 2496.705 1401.015 2497.385 ;
        RECT 1401.765 2495.685 1401.935 2497.385 ;
        RECT 1414.185 2495.515 1414.355 2495.855 ;
        RECT 1414.185 2495.345 1414.815 2495.515 ;
        RECT 1473.985 2495.345 1474.155 2496.535 ;
        RECT 1535.165 2495.345 1535.335 2496.535 ;
        RECT 1631.765 2495.685 1631.935 2496.875 ;
        RECT 1656.145 2495.685 1656.315 2496.875 ;
      LAYER mcon ;
        RECT 1292.285 2496.705 1292.455 2496.875 ;
        RECT 1197.065 2495.345 1197.235 2495.515 ;
        RECT 1245.365 2495.345 1245.535 2495.515 ;
        RECT 1341.965 2496.705 1342.135 2496.875 ;
        RECT 1390.265 2496.705 1390.435 2496.875 ;
        RECT 1631.765 2496.705 1631.935 2496.875 ;
        RECT 1473.985 2496.365 1474.155 2496.535 ;
        RECT 1414.185 2495.685 1414.355 2495.855 ;
        RECT 1414.645 2495.345 1414.815 2495.515 ;
        RECT 1535.165 2496.365 1535.335 2496.535 ;
        RECT 1656.145 2496.705 1656.315 2496.875 ;
      LAYER met1 ;
        RECT 1292.225 2496.860 1292.515 2496.905 ;
        RECT 1341.905 2496.860 1342.195 2496.905 ;
        RECT 1292.225 2496.720 1342.195 2496.860 ;
        RECT 1292.225 2496.675 1292.515 2496.720 ;
        RECT 1341.905 2496.675 1342.195 2496.720 ;
        RECT 1390.205 2496.860 1390.495 2496.905 ;
        RECT 1400.785 2496.860 1401.075 2496.905 ;
        RECT 1390.205 2496.720 1401.075 2496.860 ;
        RECT 1390.205 2496.675 1390.495 2496.720 ;
        RECT 1400.785 2496.675 1401.075 2496.720 ;
        RECT 1631.705 2496.860 1631.995 2496.905 ;
        RECT 1656.085 2496.860 1656.375 2496.905 ;
        RECT 1631.705 2496.720 1656.375 2496.860 ;
        RECT 1631.705 2496.675 1631.995 2496.720 ;
        RECT 1656.085 2496.675 1656.375 2496.720 ;
        RECT 1473.925 2496.520 1474.215 2496.565 ;
        RECT 1535.105 2496.520 1535.395 2496.565 ;
        RECT 1473.925 2496.380 1535.395 2496.520 ;
        RECT 1473.925 2496.335 1474.215 2496.380 ;
        RECT 1535.105 2496.335 1535.395 2496.380 ;
        RECT 1739.330 2496.320 1739.650 2496.580 ;
        RECT 1112.900 2496.040 1134.660 2496.180 ;
        RECT 1066.350 2495.840 1066.670 2495.900 ;
        RECT 1112.900 2495.840 1113.040 2496.040 ;
        RECT 1066.350 2495.700 1113.040 2495.840 ;
        RECT 1066.350 2495.640 1066.670 2495.700 ;
        RECT 1134.520 2495.500 1134.660 2496.040 ;
        RECT 1401.705 2495.840 1401.995 2495.885 ;
        RECT 1414.125 2495.840 1414.415 2495.885 ;
        RECT 1631.705 2495.840 1631.995 2495.885 ;
        RECT 1401.705 2495.700 1414.415 2495.840 ;
        RECT 1401.705 2495.655 1401.995 2495.700 ;
        RECT 1414.125 2495.655 1414.415 2495.700 ;
        RECT 1569.680 2495.700 1631.995 2495.840 ;
        RECT 1197.005 2495.500 1197.295 2495.545 ;
        RECT 1134.520 2495.360 1197.295 2495.500 ;
        RECT 1197.005 2495.315 1197.295 2495.360 ;
        RECT 1245.305 2495.500 1245.595 2495.545 ;
        RECT 1292.225 2495.500 1292.515 2495.545 ;
        RECT 1245.305 2495.360 1292.515 2495.500 ;
        RECT 1245.305 2495.315 1245.595 2495.360 ;
        RECT 1292.225 2495.315 1292.515 2495.360 ;
        RECT 1341.905 2495.500 1342.195 2495.545 ;
        RECT 1390.205 2495.500 1390.495 2495.545 ;
        RECT 1341.905 2495.360 1390.495 2495.500 ;
        RECT 1341.905 2495.315 1342.195 2495.360 ;
        RECT 1390.205 2495.315 1390.495 2495.360 ;
        RECT 1414.585 2495.500 1414.875 2495.545 ;
        RECT 1473.925 2495.500 1474.215 2495.545 ;
        RECT 1414.585 2495.360 1474.215 2495.500 ;
        RECT 1414.585 2495.315 1414.875 2495.360 ;
        RECT 1473.925 2495.315 1474.215 2495.360 ;
        RECT 1535.105 2495.500 1535.395 2495.545 ;
        RECT 1569.680 2495.500 1569.820 2495.700 ;
        RECT 1631.705 2495.655 1631.995 2495.700 ;
        RECT 1656.085 2495.840 1656.375 2495.885 ;
        RECT 1739.420 2495.840 1739.560 2496.320 ;
        RECT 1656.085 2495.700 1680.680 2495.840 ;
        RECT 1656.085 2495.655 1656.375 2495.700 ;
        RECT 1535.105 2495.360 1569.820 2495.500 ;
        RECT 1680.540 2495.500 1680.680 2495.700 ;
        RECT 1724.700 2495.700 1739.560 2495.840 ;
        RECT 1724.700 2495.500 1724.840 2495.700 ;
        RECT 1680.540 2495.360 1724.840 2495.500 ;
        RECT 1535.105 2495.315 1535.395 2495.360 ;
        RECT 1197.005 2494.480 1197.295 2494.525 ;
        RECT 1245.305 2494.480 1245.595 2494.525 ;
        RECT 1197.005 2494.340 1245.595 2494.480 ;
        RECT 1197.005 2494.295 1197.295 2494.340 ;
        RECT 1245.305 2494.295 1245.595 2494.340 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 1066.350 1545.540 1066.670 1545.600 ;
        RECT 16.630 1545.400 1066.670 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 1066.350 1545.340 1066.670 1545.400 ;
      LAYER via ;
        RECT 1739.360 2496.320 1739.620 2496.580 ;
        RECT 1066.380 2495.640 1066.640 2495.900 ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 1066.380 1545.340 1066.640 1545.600 ;
      LAYER met2 ;
        RECT 1740.270 2496.690 1740.550 2500.000 ;
        RECT 1739.420 2496.610 1740.550 2496.690 ;
        RECT 1739.360 2496.550 1740.550 2496.610 ;
        RECT 1739.360 2496.290 1739.620 2496.550 ;
        RECT 1740.270 2496.000 1740.550 2496.550 ;
        RECT 1066.380 2495.610 1066.640 2495.930 ;
        RECT 1066.440 1545.630 1066.580 2495.610 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 1066.380 1545.310 1066.640 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1543.340 0.300 1544.540 ;
=======
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1045.650 2509.100 1045.970 2509.160 ;
        RECT 1759.570 2509.100 1759.890 2509.160 ;
        RECT 1045.650 2508.960 1759.890 2509.100 ;
        RECT 1045.650 2508.900 1045.970 2508.960 ;
        RECT 1759.570 2508.900 1759.890 2508.960 ;
        RECT 15.710 1331.680 16.030 1331.740 ;
        RECT 1045.650 1331.680 1045.970 1331.740 ;
        RECT 15.710 1331.540 1045.970 1331.680 ;
        RECT 15.710 1331.480 16.030 1331.540 ;
        RECT 1045.650 1331.480 1045.970 1331.540 ;
      LAYER via ;
        RECT 1045.680 2508.900 1045.940 2509.160 ;
        RECT 1759.600 2508.900 1759.860 2509.160 ;
        RECT 15.740 1331.480 16.000 1331.740 ;
        RECT 1045.680 1331.480 1045.940 1331.740 ;
      LAYER met2 ;
        RECT 1045.680 2508.870 1045.940 2509.190 ;
        RECT 1759.600 2508.870 1759.860 2509.190 ;
        RECT 1045.740 1331.770 1045.880 2508.870 ;
        RECT 1759.660 2500.000 1759.800 2508.870 ;
        RECT 1759.590 2496.000 1759.870 2500.000 ;
        RECT 15.740 1331.450 16.000 1331.770 ;
        RECT 1045.680 1331.450 1045.940 1331.770 ;
        RECT 15.800 1328.565 15.940 1331.450 ;
        RECT 15.730 1328.195 16.010 1328.565 ;
      LAYER via2 ;
        RECT 15.730 1328.240 16.010 1328.520 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1327.780 0.300 1328.980 ;
=======
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 15.705 1328.530 16.035 1328.545 ;
        RECT -4.800 1328.230 16.035 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
<<<<<<< HEAD
        RECT 13.865 1328.215 14.195 1328.230 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 15.705 1328.215 16.035 1328.230 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1058.990 2500.940 1059.310 2501.000 ;
        RECT 1778.890 2500.940 1779.210 2501.000 ;
        RECT 1058.990 2500.800 1779.210 2500.940 ;
        RECT 1058.990 2500.740 1059.310 2500.800 ;
        RECT 1778.890 2500.740 1779.210 2500.800 ;
        RECT 16.630 1117.820 16.950 1117.880 ;
        RECT 1058.990 1117.820 1059.310 1117.880 ;
        RECT 16.630 1117.680 1059.310 1117.820 ;
        RECT 16.630 1117.620 16.950 1117.680 ;
        RECT 1058.990 1117.620 1059.310 1117.680 ;
      LAYER via ;
        RECT 1059.020 2500.740 1059.280 2501.000 ;
        RECT 1778.920 2500.740 1779.180 2501.000 ;
        RECT 16.660 1117.620 16.920 1117.880 ;
        RECT 1059.020 1117.620 1059.280 1117.880 ;
      LAYER met2 ;
        RECT 1059.020 2500.710 1059.280 2501.030 ;
        RECT 1778.920 2500.710 1779.180 2501.030 ;
        RECT 1059.080 1117.910 1059.220 2500.710 ;
        RECT 1778.980 2500.000 1779.120 2500.710 ;
        RECT 1778.910 2496.000 1779.190 2500.000 ;
        RECT 16.660 1117.590 16.920 1117.910 ;
        RECT 1059.020 1117.590 1059.280 1117.910 ;
        RECT 16.720 1113.005 16.860 1117.590 ;
        RECT 16.650 1112.635 16.930 1113.005 ;
      LAYER via2 ;
        RECT 16.650 1112.680 16.930 1112.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1112.220 0.300 1113.420 ;
=======
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 16.625 1112.970 16.955 1112.985 ;
        RECT -4.800 1112.670 16.955 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
<<<<<<< HEAD
        RECT 13.865 1112.655 14.195 1112.670 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 1112.655 16.955 1112.670 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1796.905 2494.665 1797.075 2496.875 ;
      LAYER mcon ;
        RECT 1796.905 2496.705 1797.075 2496.875 ;
      LAYER met1 ;
        RECT 1796.830 2496.860 1797.150 2496.920 ;
        RECT 1796.635 2496.720 1797.150 2496.860 ;
        RECT 1796.830 2496.660 1797.150 2496.720 ;
        RECT 1079.690 2494.820 1080.010 2494.880 ;
        RECT 1796.845 2494.820 1797.135 2494.865 ;
        RECT 1079.690 2494.680 1797.135 2494.820 ;
        RECT 1079.690 2494.620 1080.010 2494.680 ;
        RECT 1796.845 2494.635 1797.135 2494.680 ;
        RECT 16.630 903.960 16.950 904.020 ;
        RECT 1079.690 903.960 1080.010 904.020 ;
        RECT 16.630 903.820 1080.010 903.960 ;
        RECT 16.630 903.760 16.950 903.820 ;
        RECT 1079.690 903.760 1080.010 903.820 ;
      LAYER via ;
        RECT 1796.860 2496.660 1797.120 2496.920 ;
        RECT 1079.720 2494.620 1079.980 2494.880 ;
        RECT 16.660 903.760 16.920 904.020 ;
        RECT 1079.720 903.760 1079.980 904.020 ;
      LAYER met2 ;
        RECT 1796.860 2496.690 1797.120 2496.950 ;
        RECT 1798.230 2496.690 1798.510 2500.000 ;
        RECT 1796.860 2496.630 1798.510 2496.690 ;
        RECT 1796.920 2496.550 1798.510 2496.630 ;
        RECT 1798.230 2496.000 1798.510 2496.550 ;
        RECT 1079.720 2494.590 1079.980 2494.910 ;
        RECT 1079.780 904.050 1079.920 2494.590 ;
        RECT 16.660 903.730 16.920 904.050 ;
        RECT 1079.720 903.730 1079.980 904.050 ;
        RECT 16.720 897.445 16.860 903.730 ;
        RECT 16.650 897.075 16.930 897.445 ;
      LAYER via2 ;
        RECT 16.650 897.120 16.930 897.400 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 896.660 0.300 897.860 ;
=======
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.625 897.410 16.955 897.425 ;
        RECT -4.800 897.110 16.955 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
<<<<<<< HEAD
        RECT 13.865 897.095 14.195 897.110 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 897.095 16.955 897.110 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1065.890 2508.420 1066.210 2508.480 ;
        RECT 1817.530 2508.420 1817.850 2508.480 ;
        RECT 1065.890 2508.280 1817.850 2508.420 ;
        RECT 1065.890 2508.220 1066.210 2508.280 ;
        RECT 1817.530 2508.220 1817.850 2508.280 ;
        RECT 17.550 682.960 17.870 683.020 ;
        RECT 1065.890 682.960 1066.210 683.020 ;
        RECT 17.550 682.820 1066.210 682.960 ;
        RECT 17.550 682.760 17.870 682.820 ;
        RECT 1065.890 682.760 1066.210 682.820 ;
      LAYER via ;
        RECT 1065.920 2508.220 1066.180 2508.480 ;
        RECT 1817.560 2508.220 1817.820 2508.480 ;
        RECT 17.580 682.760 17.840 683.020 ;
        RECT 1065.920 682.760 1066.180 683.020 ;
      LAYER met2 ;
        RECT 1065.920 2508.190 1066.180 2508.510 ;
        RECT 1817.560 2508.190 1817.820 2508.510 ;
        RECT 1065.980 683.050 1066.120 2508.190 ;
        RECT 1817.620 2500.000 1817.760 2508.190 ;
        RECT 1817.550 2496.000 1817.830 2500.000 ;
        RECT 17.580 682.730 17.840 683.050 ;
        RECT 1065.920 682.730 1066.180 683.050 ;
        RECT 17.640 681.885 17.780 682.730 ;
        RECT 17.570 681.515 17.850 681.885 ;
      LAYER via2 ;
        RECT 17.570 681.560 17.850 681.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 681.100 0.300 682.300 ;
=======
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 17.545 681.850 17.875 681.865 ;
        RECT -4.800 681.550 17.875 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
<<<<<<< HEAD
        RECT 18.465 681.535 18.795 681.550 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 17.545 681.535 17.875 681.550 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1017.590 2497.880 1017.910 2497.940 ;
        RECT 1835.470 2497.880 1835.790 2497.940 ;
        RECT 1017.590 2497.740 1835.790 2497.880 ;
        RECT 1017.590 2497.680 1017.910 2497.740 ;
        RECT 1835.470 2497.680 1835.790 2497.740 ;
        RECT 17.550 469.100 17.870 469.160 ;
        RECT 1017.590 469.100 1017.910 469.160 ;
        RECT 17.550 468.960 1017.910 469.100 ;
        RECT 17.550 468.900 17.870 468.960 ;
        RECT 1017.590 468.900 1017.910 468.960 ;
      LAYER via ;
        RECT 1017.620 2497.680 1017.880 2497.940 ;
        RECT 1835.500 2497.680 1835.760 2497.940 ;
        RECT 17.580 468.900 17.840 469.160 ;
        RECT 1017.620 468.900 1017.880 469.160 ;
      LAYER met2 ;
        RECT 1836.870 2498.050 1837.150 2500.000 ;
        RECT 1835.560 2497.970 1837.150 2498.050 ;
        RECT 1017.620 2497.650 1017.880 2497.970 ;
        RECT 1835.500 2497.910 1837.150 2497.970 ;
        RECT 1835.500 2497.650 1835.760 2497.910 ;
        RECT 1017.680 469.190 1017.820 2497.650 ;
        RECT 1836.870 2496.000 1837.150 2497.910 ;
        RECT 17.580 468.870 17.840 469.190 ;
        RECT 1017.620 468.870 1017.880 469.190 ;
        RECT 17.640 466.325 17.780 468.870 ;
        RECT 17.570 465.955 17.850 466.325 ;
      LAYER via2 ;
        RECT 17.570 466.000 17.850 466.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 465.540 0.300 466.740 ;
=======
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.545 466.290 17.875 466.305 ;
        RECT -4.800 465.990 17.875 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
<<<<<<< HEAD
        RECT 13.865 465.975 14.195 465.990 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 17.545 465.975 17.875 465.990 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1855.785 2492.965 1855.955 2496.535 ;
      LAYER mcon ;
        RECT 1855.785 2496.365 1855.955 2496.535 ;
      LAYER met1 ;
        RECT 1855.710 2496.520 1856.030 2496.580 ;
        RECT 1855.515 2496.380 1856.030 2496.520 ;
        RECT 1855.710 2496.320 1856.030 2496.380 ;
        RECT 1045.190 2493.120 1045.510 2493.180 ;
        RECT 1855.725 2493.120 1856.015 2493.165 ;
        RECT 1045.190 2492.980 1856.015 2493.120 ;
        RECT 1045.190 2492.920 1045.510 2492.980 ;
        RECT 1855.725 2492.935 1856.015 2492.980 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 1045.190 255.240 1045.510 255.300 ;
        RECT 17.090 255.100 1045.510 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 1045.190 255.040 1045.510 255.100 ;
      LAYER via ;
        RECT 1855.740 2496.320 1856.000 2496.580 ;
        RECT 1045.220 2492.920 1045.480 2493.180 ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 1045.220 255.040 1045.480 255.300 ;
      LAYER met2 ;
        RECT 1856.190 2496.690 1856.470 2500.000 ;
        RECT 1855.800 2496.610 1856.470 2496.690 ;
        RECT 1855.740 2496.550 1856.470 2496.610 ;
        RECT 1855.740 2496.290 1856.000 2496.550 ;
        RECT 1856.190 2496.000 1856.470 2496.550 ;
        RECT 1045.220 2492.890 1045.480 2493.210 ;
        RECT 1045.280 255.330 1045.420 2492.890 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 1045.220 255.010 1045.480 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 249.980 0.300 251.180 ;
=======
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
<<<<<<< HEAD
        RECT 13.865 250.415 14.195 250.430 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 17.085 250.415 17.415 250.430 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 65.390 2505.360 65.710 2505.420 ;
        RECT 1875.490 2505.360 1875.810 2505.420 ;
        RECT 65.390 2505.220 1875.810 2505.360 ;
        RECT 65.390 2505.160 65.710 2505.220 ;
        RECT 1875.490 2505.160 1875.810 2505.220 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 65.390 41.380 65.710 41.440 ;
        RECT 17.090 41.240 65.710 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 65.390 41.180 65.710 41.240 ;
      LAYER via ;
        RECT 65.420 2505.160 65.680 2505.420 ;
        RECT 1875.520 2505.160 1875.780 2505.420 ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 65.420 41.180 65.680 41.440 ;
      LAYER met2 ;
        RECT 65.420 2505.130 65.680 2505.450 ;
        RECT 1875.520 2505.130 1875.780 2505.450 ;
        RECT 65.480 41.470 65.620 2505.130 ;
        RECT 1875.580 2500.000 1875.720 2505.130 ;
        RECT 1875.510 2496.000 1875.790 2500.000 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 65.420 41.150 65.680 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT -4.800 35.100 0.300 36.300 ;
=======
        RECT 17.085 2515.130 17.415 2515.145 ;
        RECT 1893.425 2515.130 1893.755 2515.145 ;
        RECT 17.085 2514.830 1893.755 2515.130 ;
        RECT 17.085 2514.815 17.415 2514.830 ;
        RECT 1893.425 2514.815 1893.755 2514.830 ;
=======
>>>>>>> re-updated local openlane
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1883.770 905.660 1884.090 905.720 ;
        RECT 1898.490 905.660 1898.810 905.720 ;
        RECT 1883.770 905.520 1898.810 905.660 ;
        RECT 1883.770 905.460 1884.090 905.520 ;
        RECT 1898.490 905.460 1898.810 905.520 ;
        RECT 1932.070 905.320 1932.390 905.380 ;
        RECT 1970.250 905.320 1970.570 905.380 ;
        RECT 1932.070 905.180 1970.570 905.320 ;
        RECT 1932.070 905.120 1932.390 905.180 ;
        RECT 1970.250 905.120 1970.570 905.180 ;
        RECT 2283.510 905.320 2283.830 905.380 ;
        RECT 2318.010 905.320 2318.330 905.380 ;
        RECT 2283.510 905.180 2318.330 905.320 ;
        RECT 2283.510 905.120 2283.830 905.180 ;
        RECT 2318.010 905.120 2318.330 905.180 ;
        RECT 1799.130 904.980 1799.450 905.040 ;
        RECT 1801.890 904.980 1802.210 905.040 ;
        RECT 1799.130 904.840 1802.210 904.980 ;
        RECT 1799.130 904.780 1799.450 904.840 ;
        RECT 1801.890 904.780 1802.210 904.840 ;
        RECT 2476.710 904.640 2477.030 904.700 ;
        RECT 2504.310 904.640 2504.630 904.700 ;
        RECT 2476.710 904.500 2504.630 904.640 ;
        RECT 2476.710 904.440 2477.030 904.500 ;
        RECT 2504.310 904.440 2504.630 904.500 ;
        RECT 1642.270 904.300 1642.590 904.360 ;
        RECT 1690.110 904.300 1690.430 904.360 ;
        RECT 1642.270 904.160 1690.430 904.300 ;
        RECT 1642.270 904.100 1642.590 904.160 ;
        RECT 1690.110 904.100 1690.430 904.160 ;
      LAYER via ;
        RECT 1883.800 905.460 1884.060 905.720 ;
        RECT 1898.520 905.460 1898.780 905.720 ;
        RECT 1932.100 905.120 1932.360 905.380 ;
        RECT 1970.280 905.120 1970.540 905.380 ;
        RECT 2283.540 905.120 2283.800 905.380 ;
        RECT 2318.040 905.120 2318.300 905.380 ;
        RECT 1799.160 904.780 1799.420 905.040 ;
        RECT 1801.920 904.780 1802.180 905.040 ;
        RECT 2476.740 904.440 2477.000 904.700 ;
        RECT 2504.340 904.440 2504.600 904.700 ;
        RECT 1642.300 904.100 1642.560 904.360 ;
        RECT 1690.140 904.100 1690.400 904.360 ;
      LAYER met2 ;
        RECT 1217.710 2498.050 1217.990 2500.000 ;
        RECT 1219.550 2498.050 1219.830 2498.165 ;
        RECT 1217.710 2497.910 1219.830 2498.050 ;
        RECT 1217.710 2496.000 1217.990 2497.910 ;
        RECT 1219.550 2497.795 1219.830 2497.910 ;
        RECT 1970.270 905.915 1970.550 906.285 ;
        RECT 1883.800 905.605 1884.060 905.750 ;
        RECT 1898.520 905.605 1898.780 905.750 ;
        RECT 1690.130 905.235 1690.410 905.605 ;
        RECT 1883.790 905.235 1884.070 905.605 ;
        RECT 1898.510 905.235 1898.790 905.605 ;
        RECT 1970.340 905.410 1970.480 905.915 ;
        RECT 1606.410 904.555 1606.690 904.925 ;
        RECT 1606.480 902.885 1606.620 904.555 ;
        RECT 1690.200 904.390 1690.340 905.235 ;
        RECT 1932.100 905.090 1932.360 905.410 ;
        RECT 1970.280 905.090 1970.540 905.410 ;
        RECT 2283.530 905.235 2283.810 905.605 ;
        RECT 2318.030 905.235 2318.310 905.605 ;
        RECT 2573.330 905.235 2573.610 905.605 ;
        RECT 2283.540 905.090 2283.800 905.235 ;
        RECT 2318.040 905.090 2318.300 905.235 ;
        RECT 1799.160 904.925 1799.420 905.070 ;
        RECT 1801.920 904.925 1802.180 905.070 ;
        RECT 1932.160 904.925 1932.300 905.090 ;
        RECT 1799.150 904.555 1799.430 904.925 ;
        RECT 1801.910 904.555 1802.190 904.925 ;
        RECT 1932.090 904.555 1932.370 904.925 ;
        RECT 1993.730 904.810 1994.010 904.925 ;
        RECT 1994.650 904.810 1994.930 904.925 ;
        RECT 1993.730 904.670 1994.930 904.810 ;
        RECT 1993.730 904.555 1994.010 904.670 ;
        RECT 1994.650 904.555 1994.930 904.670 ;
        RECT 2476.730 904.555 2477.010 904.925 ;
        RECT 2573.400 904.810 2573.540 905.235 ;
        RECT 2574.250 904.810 2574.530 904.925 ;
        RECT 2476.740 904.410 2477.000 904.555 ;
        RECT 2504.340 904.410 2504.600 904.730 ;
        RECT 2573.400 904.670 2574.530 904.810 ;
        RECT 2574.250 904.555 2574.530 904.670 ;
        RECT 1642.300 904.245 1642.560 904.390 ;
        RECT 1642.290 903.875 1642.570 904.245 ;
        RECT 1690.140 904.070 1690.400 904.390 ;
        RECT 2504.400 904.245 2504.540 904.410 ;
        RECT 2504.330 903.875 2504.610 904.245 ;
        RECT 1606.410 902.515 1606.690 902.885 ;
      LAYER via2 ;
        RECT 1219.550 2497.840 1219.830 2498.120 ;
        RECT 1970.270 905.960 1970.550 906.240 ;
        RECT 1690.130 905.280 1690.410 905.560 ;
        RECT 1883.790 905.280 1884.070 905.560 ;
        RECT 1898.510 905.280 1898.790 905.560 ;
        RECT 1606.410 904.600 1606.690 904.880 ;
        RECT 2283.530 905.280 2283.810 905.560 ;
        RECT 2318.030 905.280 2318.310 905.560 ;
        RECT 2573.330 905.280 2573.610 905.560 ;
        RECT 1799.150 904.600 1799.430 904.880 ;
        RECT 1801.910 904.600 1802.190 904.880 ;
        RECT 1932.090 904.600 1932.370 904.880 ;
        RECT 1993.730 904.600 1994.010 904.880 ;
        RECT 1994.650 904.600 1994.930 904.880 ;
        RECT 2476.730 904.600 2477.010 904.880 ;
        RECT 2574.250 904.600 2574.530 904.880 ;
        RECT 1642.290 903.920 1642.570 904.200 ;
        RECT 2504.330 903.920 2504.610 904.200 ;
        RECT 1606.410 902.560 1606.690 902.840 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 908.900 2924.800 910.100 ;
=======
        RECT 1219.985 2498.140 1220.315 2498.145 ;
        RECT 1219.985 2498.130 1220.570 2498.140 ;
        RECT 1219.985 2497.830 1220.770 2498.130 ;
        RECT 1219.985 2497.820 1220.570 2497.830 ;
        RECT 1219.985 2497.815 1220.315 2497.820 ;
=======
        RECT 1219.525 2498.130 1219.855 2498.145 ;
        RECT 1220.190 2498.130 1220.570 2498.140 ;
        RECT 1219.525 2497.830 1220.570 2498.130 ;
        RECT 1219.525 2497.815 1219.855 2497.830 ;
        RECT 1220.190 2497.820 1220.570 2497.830 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2916.710 909.350 2924.800 909.650 ;
        RECT 1441.910 906.930 1442.290 906.940 ;
        RECT 1441.910 906.630 1490.090 906.930 ;
        RECT 1441.910 906.620 1442.290 906.630 ;
        RECT 1345.310 906.250 1345.690 906.260 ;
        RECT 1489.790 906.250 1490.090 906.630 ;
        RECT 1970.245 906.250 1970.575 906.265 ;
        RECT 1980.110 906.250 1980.490 906.260 ;
        RECT 1268.990 905.950 1318.970 906.250 ;
        RECT 1220.190 904.890 1220.570 904.900 ;
        RECT 1268.990 904.890 1269.290 905.950 ;
        RECT 1220.190 904.590 1269.290 904.890 ;
        RECT 1318.670 904.890 1318.970 905.950 ;
        RECT 1345.310 905.950 1370.490 906.250 ;
        RECT 1489.790 905.950 1509.410 906.250 ;
        RECT 1345.310 905.940 1345.690 905.950 ;
        RECT 1370.190 905.570 1370.490 905.950 ;
        RECT 1440.990 905.570 1441.370 905.580 ;
        RECT 1370.190 905.270 1441.370 905.570 ;
        RECT 1440.990 905.260 1441.370 905.270 ;
        RECT 1345.310 904.890 1345.690 904.900 ;
        RECT 1318.670 904.590 1345.690 904.890 ;
        RECT 1220.190 904.580 1220.570 904.590 ;
        RECT 1345.310 904.580 1345.690 904.590 ;
        RECT 1509.110 904.210 1509.410 905.950 ;
        RECT 1970.245 905.950 1980.490 906.250 ;
        RECT 1970.245 905.935 1970.575 905.950 ;
        RECT 1980.110 905.940 1980.490 905.950 ;
        RECT 1690.105 905.570 1690.435 905.585 ;
        RECT 1883.765 905.570 1884.095 905.585 ;
        RECT 1690.105 905.270 1704.450 905.570 ;
        RECT 1690.105 905.255 1690.435 905.270 ;
        RECT 1606.385 904.890 1606.715 904.905 ;
        RECT 1559.710 904.590 1606.715 904.890 ;
        RECT 1559.710 904.210 1560.010 904.590 ;
        RECT 1606.385 904.575 1606.715 904.590 ;
        RECT 1642.265 904.210 1642.595 904.225 ;
        RECT 1509.110 903.910 1560.010 904.210 ;
        RECT 1641.590 903.910 1642.595 904.210 ;
        RECT 1704.150 904.210 1704.450 905.270 ;
        RECT 1849.510 905.270 1884.095 905.570 ;
        RECT 1799.125 904.890 1799.455 904.905 ;
        RECT 1752.910 904.590 1799.455 904.890 ;
        RECT 1752.910 904.210 1753.210 904.590 ;
        RECT 1799.125 904.575 1799.455 904.590 ;
        RECT 1801.885 904.890 1802.215 904.905 ;
        RECT 1801.885 904.590 1835.090 904.890 ;
        RECT 1801.885 904.575 1802.215 904.590 ;
        RECT 1704.150 903.910 1753.210 904.210 ;
        RECT 1834.790 904.210 1835.090 904.590 ;
        RECT 1849.510 904.210 1849.810 905.270 ;
        RECT 1883.765 905.255 1884.095 905.270 ;
        RECT 1898.485 905.570 1898.815 905.585 ;
        RECT 2283.505 905.570 2283.835 905.585 ;
        RECT 1898.485 905.270 1931.690 905.570 ;
        RECT 1898.485 905.255 1898.815 905.270 ;
        RECT 1931.390 904.890 1931.690 905.270 ;
        RECT 2062.950 905.270 2090.850 905.570 ;
        RECT 1932.065 904.890 1932.395 904.905 ;
        RECT 1931.390 904.590 1932.395 904.890 ;
        RECT 1932.065 904.575 1932.395 904.590 ;
        RECT 1980.110 904.890 1980.490 904.900 ;
        RECT 1993.705 904.890 1994.035 904.905 ;
        RECT 1980.110 904.590 1994.035 904.890 ;
        RECT 1980.110 904.580 1980.490 904.590 ;
        RECT 1993.705 904.575 1994.035 904.590 ;
        RECT 1994.625 904.890 1994.955 904.905 ;
        RECT 1994.625 904.590 2042.090 904.890 ;
        RECT 1994.625 904.575 1994.955 904.590 ;
        RECT 1834.790 903.910 1849.810 904.210 ;
        RECT 2041.790 904.210 2042.090 904.590 ;
        RECT 2062.950 904.210 2063.250 905.270 ;
        RECT 2090.550 904.890 2090.850 905.270 ;
        RECT 2159.550 905.270 2283.835 905.570 ;
        RECT 2090.550 904.590 2138.690 904.890 ;
        RECT 2041.790 903.910 2063.250 904.210 ;
        RECT 2138.390 904.210 2138.690 904.590 ;
        RECT 2159.550 904.210 2159.850 905.270 ;
        RECT 2283.505 905.255 2283.835 905.270 ;
        RECT 2318.005 905.570 2318.335 905.585 ;
        RECT 2573.305 905.570 2573.635 905.585 ;
        RECT 2318.005 905.270 2331.890 905.570 ;
        RECT 2318.005 905.255 2318.335 905.270 ;
        RECT 2138.390 903.910 2159.850 904.210 ;
        RECT 2331.590 904.210 2331.890 905.270 ;
        RECT 2380.350 905.270 2428.490 905.570 ;
        RECT 2380.350 904.210 2380.650 905.270 ;
        RECT 2331.590 903.910 2380.650 904.210 ;
        RECT 2428.190 904.210 2428.490 905.270 ;
        RECT 2553.310 905.270 2573.635 905.570 ;
        RECT 2476.705 904.890 2477.035 904.905 ;
        RECT 2553.310 904.890 2553.610 905.270 ;
        RECT 2573.305 905.255 2573.635 905.270 ;
        RECT 2739.150 905.270 2787.290 905.570 ;
        RECT 2429.110 904.590 2477.035 904.890 ;
        RECT 2429.110 904.210 2429.410 904.590 ;
        RECT 2476.705 904.575 2477.035 904.590 ;
        RECT 2525.710 904.590 2553.610 904.890 ;
        RECT 2574.225 904.890 2574.555 904.905 ;
        RECT 2574.225 904.590 2621.690 904.890 ;
        RECT 2428.190 903.910 2429.410 904.210 ;
        RECT 2504.305 904.210 2504.635 904.225 ;
        RECT 2525.710 904.210 2526.010 904.590 ;
        RECT 2574.225 904.575 2574.555 904.590 ;
        RECT 2504.305 903.910 2526.010 904.210 ;
        RECT 2621.390 904.210 2621.690 904.590 ;
        RECT 2739.150 904.210 2739.450 905.270 ;
        RECT 2621.390 903.910 2739.450 904.210 ;
        RECT 2786.990 904.210 2787.290 905.270 ;
        RECT 2787.910 905.270 2836.050 905.570 ;
        RECT 2787.910 904.210 2788.210 905.270 ;
        RECT 2835.750 904.890 2836.050 905.270 ;
        RECT 2916.710 904.890 2917.010 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
        RECT 2835.750 904.590 2883.890 904.890 ;
        RECT 2786.990 903.910 2788.210 904.210 ;
        RECT 2883.590 904.210 2883.890 904.590 ;
        RECT 2884.510 904.590 2917.010 904.890 ;
        RECT 2884.510 904.210 2884.810 904.590 ;
        RECT 2883.590 903.910 2884.810 904.210 ;
        RECT 1606.385 902.850 1606.715 902.865 ;
        RECT 1641.590 902.850 1641.890 903.910 ;
        RECT 1642.265 903.895 1642.595 903.910 ;
        RECT 2504.305 903.895 2504.635 903.910 ;
        RECT 1606.385 902.550 1641.890 902.850 ;
        RECT 1606.385 902.535 1606.715 902.550 ;
      LAYER via3 ;
        RECT 1220.220 2497.820 1220.540 2498.140 ;
        RECT 1441.940 906.620 1442.260 906.940 ;
        RECT 1220.220 904.580 1220.540 904.900 ;
        RECT 1345.340 905.940 1345.660 906.260 ;
        RECT 1441.020 905.260 1441.340 905.580 ;
        RECT 1345.340 904.580 1345.660 904.900 ;
        RECT 1980.140 905.940 1980.460 906.260 ;
        RECT 1980.140 904.580 1980.460 904.900 ;
      LAYER met4 ;
        RECT 1220.215 2497.815 1220.545 2498.145 ;
        RECT 1220.230 904.905 1220.530 2497.815 ;
        RECT 1441.935 906.615 1442.265 906.945 ;
        RECT 1345.335 905.935 1345.665 906.265 ;
        RECT 1441.950 906.250 1442.250 906.615 ;
        RECT 1441.030 905.950 1442.250 906.250 ;
        RECT 1345.350 904.905 1345.650 905.935 ;
        RECT 1441.030 905.585 1441.330 905.950 ;
        RECT 1980.135 905.935 1980.465 906.265 ;
        RECT 1441.015 905.255 1441.345 905.585 ;
        RECT 1980.150 904.905 1980.450 905.935 ;
        RECT 1220.215 904.575 1220.545 904.905 ;
        RECT 1345.335 904.575 1345.665 904.905 ;
<<<<<<< HEAD
        RECT 1346.255 904.575 1346.585 904.905 ;
        RECT 1345.350 902.850 1345.650 904.575 ;
        RECT 1346.270 902.850 1346.570 904.575 ;
        RECT 1345.350 902.550 1346.570 902.850 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1980.135 904.575 1980.465 904.905 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1973.470 1140.600 1973.790 1140.660 ;
        RECT 1997.850 1140.600 1998.170 1140.660 ;
        RECT 1973.470 1140.460 1998.170 1140.600 ;
        RECT 1973.470 1140.400 1973.790 1140.460 ;
        RECT 1997.850 1140.400 1998.170 1140.460 ;
        RECT 1390.190 1139.920 1390.510 1139.980 ;
        RECT 1421.010 1139.920 1421.330 1139.980 ;
        RECT 1390.190 1139.780 1421.330 1139.920 ;
        RECT 1390.190 1139.720 1390.510 1139.780 ;
        RECT 1421.010 1139.720 1421.330 1139.780 ;
        RECT 2607.810 1139.920 2608.130 1139.980 ;
        RECT 2625.750 1139.920 2626.070 1139.980 ;
        RECT 2607.810 1139.780 2626.070 1139.920 ;
        RECT 2607.810 1139.720 2608.130 1139.780 ;
        RECT 2625.750 1139.720 2626.070 1139.780 ;
        RECT 1435.270 1139.580 1435.590 1139.640 ;
        RECT 1483.110 1139.580 1483.430 1139.640 ;
        RECT 1435.270 1139.440 1483.430 1139.580 ;
        RECT 1435.270 1139.380 1435.590 1139.440 ;
        RECT 1483.110 1139.380 1483.430 1139.440 ;
        RECT 1799.130 1139.580 1799.450 1139.640 ;
        RECT 1801.890 1139.580 1802.210 1139.640 ;
        RECT 1799.130 1139.440 1802.210 1139.580 ;
        RECT 1799.130 1139.380 1799.450 1139.440 ;
        RECT 1801.890 1139.380 1802.210 1139.440 ;
        RECT 2476.710 1139.580 2477.030 1139.640 ;
        RECT 2511.210 1139.580 2511.530 1139.640 ;
        RECT 2476.710 1139.440 2511.530 1139.580 ;
        RECT 2476.710 1139.380 2477.030 1139.440 ;
        RECT 2511.210 1139.380 2511.530 1139.440 ;
        RECT 1642.270 1138.900 1642.590 1138.960 ;
        RECT 1690.110 1138.900 1690.430 1138.960 ;
        RECT 1642.270 1138.760 1690.430 1138.900 ;
        RECT 1642.270 1138.700 1642.590 1138.760 ;
        RECT 1690.110 1138.700 1690.430 1138.760 ;
        RECT 2649.670 1138.900 2649.990 1138.960 ;
        RECT 2697.510 1138.900 2697.830 1138.960 ;
        RECT 2649.670 1138.760 2697.830 1138.900 ;
        RECT 2649.670 1138.700 2649.990 1138.760 ;
        RECT 2697.510 1138.700 2697.830 1138.760 ;
      LAYER via ;
        RECT 1973.500 1140.400 1973.760 1140.660 ;
        RECT 1997.880 1140.400 1998.140 1140.660 ;
        RECT 1390.220 1139.720 1390.480 1139.980 ;
        RECT 1421.040 1139.720 1421.300 1139.980 ;
        RECT 2607.840 1139.720 2608.100 1139.980 ;
        RECT 2625.780 1139.720 2626.040 1139.980 ;
        RECT 1435.300 1139.380 1435.560 1139.640 ;
        RECT 1483.140 1139.380 1483.400 1139.640 ;
        RECT 1799.160 1139.380 1799.420 1139.640 ;
        RECT 1801.920 1139.380 1802.180 1139.640 ;
        RECT 2476.740 1139.380 2477.000 1139.640 ;
        RECT 2511.240 1139.380 2511.500 1139.640 ;
        RECT 1642.300 1138.700 1642.560 1138.960 ;
        RECT 1690.140 1138.700 1690.400 1138.960 ;
        RECT 2649.700 1138.700 2649.960 1138.960 ;
        RECT 2697.540 1138.700 2697.800 1138.960 ;
      LAYER met2 ;
        RECT 1237.030 2498.050 1237.310 2500.000 ;
        RECT 1238.870 2498.050 1239.150 2498.165 ;
        RECT 1237.030 2497.910 1239.150 2498.050 ;
        RECT 1237.030 2496.000 1237.310 2497.910 ;
        RECT 1238.870 2497.795 1239.150 2497.910 ;
        RECT 1390.210 1140.515 1390.490 1140.885 ;
        RECT 1973.490 1140.515 1973.770 1140.885 ;
        RECT 1390.280 1140.010 1390.420 1140.515 ;
        RECT 1973.500 1140.370 1973.760 1140.515 ;
        RECT 1997.880 1140.370 1998.140 1140.690 ;
        RECT 2221.890 1140.515 2222.170 1140.885 ;
        RECT 1390.220 1139.690 1390.480 1140.010 ;
        RECT 1421.040 1139.690 1421.300 1140.010 ;
        RECT 1490.030 1139.835 1490.310 1140.205 ;
        RECT 1690.130 1139.835 1690.410 1140.205 ;
        RECT 1876.890 1139.835 1877.170 1140.205 ;
        RECT 1421.100 1139.525 1421.240 1139.690 ;
        RECT 1435.300 1139.525 1435.560 1139.670 ;
        RECT 1483.140 1139.525 1483.400 1139.670 ;
        RECT 1490.100 1139.525 1490.240 1139.835 ;
        RECT 1421.030 1139.155 1421.310 1139.525 ;
        RECT 1435.290 1139.155 1435.570 1139.525 ;
        RECT 1483.130 1139.155 1483.410 1139.525 ;
        RECT 1490.030 1139.155 1490.310 1139.525 ;
        RECT 1538.330 1139.155 1538.610 1139.525 ;
        RECT 1606.410 1139.155 1606.690 1139.525 ;
        RECT 1538.400 1138.845 1538.540 1139.155 ;
        RECT 1538.330 1138.475 1538.610 1138.845 ;
        RECT 1606.480 1137.485 1606.620 1139.155 ;
        RECT 1690.200 1138.990 1690.340 1139.835 ;
        RECT 1799.160 1139.525 1799.420 1139.670 ;
        RECT 1801.920 1139.525 1802.180 1139.670 ;
        RECT 1876.960 1139.525 1877.100 1139.835 ;
        RECT 1997.940 1139.525 1998.080 1140.370 ;
        RECT 1799.150 1139.155 1799.430 1139.525 ;
        RECT 1801.910 1139.155 1802.190 1139.525 ;
        RECT 1876.890 1139.155 1877.170 1139.525 ;
        RECT 1997.870 1139.155 1998.150 1139.525 ;
        RECT 1642.300 1138.845 1642.560 1138.990 ;
        RECT 1642.290 1138.475 1642.570 1138.845 ;
        RECT 1690.140 1138.670 1690.400 1138.990 ;
        RECT 2221.960 1138.845 2222.100 1140.515 ;
        RECT 2283.990 1140.090 2284.270 1140.205 ;
        RECT 2283.600 1139.950 2284.270 1140.090 ;
        RECT 2283.600 1139.525 2283.740 1139.950 ;
        RECT 2283.990 1139.835 2284.270 1139.950 ;
        RECT 2511.230 1139.835 2511.510 1140.205 ;
        RECT 2607.830 1139.835 2608.110 1140.205 ;
        RECT 2511.300 1139.670 2511.440 1139.835 ;
        RECT 2607.840 1139.690 2608.100 1139.835 ;
        RECT 2625.780 1139.690 2626.040 1140.010 ;
        RECT 2697.530 1139.835 2697.810 1140.205 ;
        RECT 2476.740 1139.525 2477.000 1139.670 ;
        RECT 2283.530 1139.155 2283.810 1139.525 ;
        RECT 2476.730 1139.155 2477.010 1139.525 ;
        RECT 2511.240 1139.350 2511.500 1139.670 ;
        RECT 2625.840 1138.845 2625.980 1139.690 ;
        RECT 2697.600 1138.990 2697.740 1139.835 ;
        RECT 2649.700 1138.845 2649.960 1138.990 ;
        RECT 2221.890 1138.475 2222.170 1138.845 ;
        RECT 2625.770 1138.475 2626.050 1138.845 ;
        RECT 2649.690 1138.475 2649.970 1138.845 ;
        RECT 2697.540 1138.670 2697.800 1138.990 ;
        RECT 1606.410 1137.115 1606.690 1137.485 ;
      LAYER via2 ;
        RECT 1238.870 2497.840 1239.150 2498.120 ;
        RECT 1390.210 1140.560 1390.490 1140.840 ;
        RECT 1973.490 1140.560 1973.770 1140.840 ;
        RECT 2221.890 1140.560 2222.170 1140.840 ;
        RECT 1490.030 1139.880 1490.310 1140.160 ;
        RECT 1690.130 1139.880 1690.410 1140.160 ;
        RECT 1876.890 1139.880 1877.170 1140.160 ;
        RECT 1421.030 1139.200 1421.310 1139.480 ;
        RECT 1435.290 1139.200 1435.570 1139.480 ;
        RECT 1483.130 1139.200 1483.410 1139.480 ;
        RECT 1490.030 1139.200 1490.310 1139.480 ;
        RECT 1538.330 1139.200 1538.610 1139.480 ;
        RECT 1606.410 1139.200 1606.690 1139.480 ;
        RECT 1538.330 1138.520 1538.610 1138.800 ;
        RECT 1799.150 1139.200 1799.430 1139.480 ;
        RECT 1801.910 1139.200 1802.190 1139.480 ;
        RECT 1876.890 1139.200 1877.170 1139.480 ;
        RECT 1997.870 1139.200 1998.150 1139.480 ;
        RECT 1642.290 1138.520 1642.570 1138.800 ;
        RECT 2283.990 1139.880 2284.270 1140.160 ;
        RECT 2511.230 1139.880 2511.510 1140.160 ;
        RECT 2607.830 1139.880 2608.110 1140.160 ;
        RECT 2697.530 1139.880 2697.810 1140.160 ;
        RECT 2283.530 1139.200 2283.810 1139.480 ;
        RECT 2476.730 1139.200 2477.010 1139.480 ;
        RECT 2221.890 1138.520 2222.170 1138.800 ;
        RECT 2625.770 1138.520 2626.050 1138.800 ;
        RECT 2649.690 1138.520 2649.970 1138.800 ;
        RECT 1606.410 1137.160 1606.690 1137.440 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1143.500 2924.800 1144.700 ;
=======
        RECT 1240.685 2498.130 1241.015 2498.145 ;
=======
        RECT 1238.845 2498.130 1239.175 2498.145 ;
>>>>>>> re-updated local openlane
        RECT 1241.350 2498.130 1241.730 2498.140 ;
        RECT 1238.845 2497.830 1241.730 2498.130 ;
        RECT 1238.845 2497.815 1239.175 2497.830 ;
        RECT 1241.350 2497.820 1241.730 2497.830 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2916.710 1143.950 2924.800 1144.250 ;
        RECT 1390.185 1140.850 1390.515 1140.865 ;
        RECT 1280.030 1140.550 1390.515 1140.850 ;
        RECT 1241.350 1140.170 1241.730 1140.180 ;
        RECT 1241.350 1139.870 1269.290 1140.170 ;
        RECT 1241.350 1139.860 1241.730 1139.870 ;
        RECT 1268.990 1139.490 1269.290 1139.870 ;
        RECT 1280.030 1139.490 1280.330 1140.550 ;
        RECT 1390.185 1140.535 1390.515 1140.550 ;
        RECT 1924.910 1140.850 1925.290 1140.860 ;
        RECT 1973.465 1140.850 1973.795 1140.865 ;
        RECT 2221.865 1140.850 2222.195 1140.865 ;
        RECT 1924.910 1140.550 1973.795 1140.850 ;
        RECT 1924.910 1140.540 1925.290 1140.550 ;
        RECT 1973.465 1140.535 1973.795 1140.550 ;
        RECT 2197.270 1140.550 2222.195 1140.850 ;
        RECT 1490.005 1140.170 1490.335 1140.185 ;
        RECT 1690.105 1140.170 1690.435 1140.185 ;
        RECT 1876.865 1140.170 1877.195 1140.185 ;
        RECT 1490.005 1139.870 1491.010 1140.170 ;
        RECT 1490.005 1139.855 1490.335 1139.870 ;
        RECT 1268.990 1139.190 1280.330 1139.490 ;
        RECT 1421.005 1139.490 1421.335 1139.505 ;
        RECT 1435.265 1139.490 1435.595 1139.505 ;
        RECT 1421.005 1139.190 1435.595 1139.490 ;
        RECT 1421.005 1139.175 1421.335 1139.190 ;
        RECT 1435.265 1139.175 1435.595 1139.190 ;
        RECT 1483.105 1139.490 1483.435 1139.505 ;
        RECT 1490.005 1139.490 1490.335 1139.505 ;
        RECT 1483.105 1139.190 1490.335 1139.490 ;
        RECT 1490.710 1139.490 1491.010 1139.870 ;
        RECT 1690.105 1139.870 1704.450 1140.170 ;
        RECT 1690.105 1139.855 1690.435 1139.870 ;
        RECT 1538.305 1139.490 1538.635 1139.505 ;
        RECT 1606.385 1139.490 1606.715 1139.505 ;
        RECT 1490.710 1139.190 1538.635 1139.490 ;
        RECT 1483.105 1139.175 1483.435 1139.190 ;
        RECT 1490.005 1139.175 1490.335 1139.190 ;
        RECT 1538.305 1139.175 1538.635 1139.190 ;
        RECT 1559.710 1139.190 1606.715 1139.490 ;
        RECT 1538.305 1138.810 1538.635 1138.825 ;
        RECT 1559.710 1138.810 1560.010 1139.190 ;
        RECT 1606.385 1139.175 1606.715 1139.190 ;
        RECT 1642.265 1138.810 1642.595 1138.825 ;
        RECT 1538.305 1138.510 1560.010 1138.810 ;
        RECT 1641.590 1138.510 1642.595 1138.810 ;
        RECT 1704.150 1138.810 1704.450 1139.870 ;
        RECT 1849.510 1139.870 1877.195 1140.170 ;
        RECT 1799.125 1139.490 1799.455 1139.505 ;
        RECT 1752.910 1139.190 1799.455 1139.490 ;
        RECT 1752.910 1138.810 1753.210 1139.190 ;
        RECT 1799.125 1139.175 1799.455 1139.190 ;
        RECT 1801.885 1139.490 1802.215 1139.505 ;
        RECT 1801.885 1139.190 1835.090 1139.490 ;
        RECT 1801.885 1139.175 1802.215 1139.190 ;
        RECT 1704.150 1138.510 1753.210 1138.810 ;
        RECT 1834.790 1138.810 1835.090 1139.190 ;
        RECT 1849.510 1138.810 1849.810 1139.870 ;
        RECT 1876.865 1139.855 1877.195 1139.870 ;
        RECT 2062.950 1139.870 2111.090 1140.170 ;
        RECT 1876.865 1139.490 1877.195 1139.505 ;
        RECT 1923.990 1139.490 1924.370 1139.500 ;
        RECT 1876.865 1139.190 1924.370 1139.490 ;
        RECT 1876.865 1139.175 1877.195 1139.190 ;
        RECT 1923.990 1139.180 1924.370 1139.190 ;
        RECT 1997.845 1139.490 1998.175 1139.505 ;
        RECT 1997.845 1139.190 2042.090 1139.490 ;
        RECT 1997.845 1139.175 1998.175 1139.190 ;
        RECT 1834.790 1138.510 1849.810 1138.810 ;
        RECT 2041.790 1138.810 2042.090 1139.190 ;
        RECT 2062.950 1138.810 2063.250 1139.870 ;
        RECT 2041.790 1138.510 2063.250 1138.810 ;
        RECT 2110.790 1138.810 2111.090 1139.870 ;
        RECT 2111.710 1139.870 2163.530 1140.170 ;
        RECT 2111.710 1138.810 2112.010 1139.870 ;
        RECT 2110.790 1138.510 2112.010 1138.810 ;
        RECT 2163.230 1138.810 2163.530 1139.870 ;
        RECT 2197.270 1138.810 2197.570 1140.550 ;
        RECT 2221.865 1140.535 2222.195 1140.550 ;
        RECT 2283.965 1140.170 2284.295 1140.185 ;
        RECT 2511.205 1140.170 2511.535 1140.185 ;
        RECT 2607.805 1140.170 2608.135 1140.185 ;
        RECT 2283.965 1139.870 2353.050 1140.170 ;
        RECT 2283.965 1139.855 2284.295 1139.870 ;
        RECT 2283.505 1139.490 2283.835 1139.505 ;
        RECT 2269.950 1139.190 2283.835 1139.490 ;
        RECT 2352.750 1139.490 2353.050 1139.870 ;
        RECT 2401.510 1139.870 2429.410 1140.170 ;
        RECT 2352.750 1139.190 2400.890 1139.490 ;
        RECT 2163.230 1138.510 2197.570 1138.810 ;
        RECT 2221.865 1138.810 2222.195 1138.825 ;
        RECT 2269.950 1138.810 2270.250 1139.190 ;
        RECT 2283.505 1139.175 2283.835 1139.190 ;
        RECT 2221.865 1138.510 2270.250 1138.810 ;
        RECT 2400.590 1138.810 2400.890 1139.190 ;
        RECT 2401.510 1138.810 2401.810 1139.870 ;
        RECT 2429.110 1139.490 2429.410 1139.870 ;
        RECT 2511.205 1139.870 2526.010 1140.170 ;
        RECT 2511.205 1139.855 2511.535 1139.870 ;
        RECT 2476.705 1139.490 2477.035 1139.505 ;
        RECT 2429.110 1139.190 2477.035 1139.490 ;
        RECT 2476.705 1139.175 2477.035 1139.190 ;
        RECT 2400.590 1138.510 2401.810 1138.810 ;
        RECT 2525.710 1138.810 2526.010 1139.870 ;
        RECT 2572.630 1139.870 2608.135 1140.170 ;
        RECT 2572.630 1138.810 2572.930 1139.870 ;
        RECT 2607.805 1139.855 2608.135 1139.870 ;
        RECT 2697.505 1140.170 2697.835 1140.185 ;
        RECT 2697.505 1139.870 2739.450 1140.170 ;
        RECT 2697.505 1139.855 2697.835 1139.870 ;
        RECT 2739.150 1139.490 2739.450 1139.870 ;
        RECT 2787.910 1139.870 2836.050 1140.170 ;
        RECT 2739.150 1139.190 2787.290 1139.490 ;
        RECT 2525.710 1138.510 2572.930 1138.810 ;
        RECT 2625.745 1138.810 2626.075 1138.825 ;
        RECT 2649.665 1138.810 2649.995 1138.825 ;
        RECT 2625.745 1138.510 2649.995 1138.810 ;
        RECT 2786.990 1138.810 2787.290 1139.190 ;
        RECT 2787.910 1138.810 2788.210 1139.870 ;
        RECT 2835.750 1139.490 2836.050 1139.870 ;
        RECT 2916.710 1139.490 2917.010 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT 2835.750 1139.190 2883.890 1139.490 ;
        RECT 2786.990 1138.510 2788.210 1138.810 ;
        RECT 2883.590 1138.810 2883.890 1139.190 ;
        RECT 2884.510 1139.190 2917.010 1139.490 ;
        RECT 2884.510 1138.810 2884.810 1139.190 ;
        RECT 2883.590 1138.510 2884.810 1138.810 ;
        RECT 1538.305 1138.495 1538.635 1138.510 ;
        RECT 1606.385 1137.450 1606.715 1137.465 ;
        RECT 1641.590 1137.450 1641.890 1138.510 ;
        RECT 1642.265 1138.495 1642.595 1138.510 ;
        RECT 2221.865 1138.495 2222.195 1138.510 ;
        RECT 2625.745 1138.495 2626.075 1138.510 ;
        RECT 2649.665 1138.495 2649.995 1138.510 ;
        RECT 1923.990 1138.130 1924.370 1138.140 ;
        RECT 1924.910 1138.130 1925.290 1138.140 ;
        RECT 1923.990 1137.830 1925.290 1138.130 ;
        RECT 1923.990 1137.820 1924.370 1137.830 ;
        RECT 1924.910 1137.820 1925.290 1137.830 ;
        RECT 1606.385 1137.150 1641.890 1137.450 ;
        RECT 1606.385 1137.135 1606.715 1137.150 ;
      LAYER via3 ;
        RECT 1241.380 2497.820 1241.700 2498.140 ;
        RECT 1241.380 1139.860 1241.700 1140.180 ;
        RECT 1924.940 1140.540 1925.260 1140.860 ;
        RECT 1924.020 1139.180 1924.340 1139.500 ;
        RECT 1924.020 1137.820 1924.340 1138.140 ;
        RECT 1924.940 1137.820 1925.260 1138.140 ;
      LAYER met4 ;
        RECT 1241.375 2497.815 1241.705 2498.145 ;
        RECT 1241.390 1140.185 1241.690 2497.815 ;
        RECT 1924.935 1140.535 1925.265 1140.865 ;
        RECT 1241.375 1139.855 1241.705 1140.185 ;
<<<<<<< HEAD
        RECT 1980.135 1139.855 1980.465 1140.185 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1924.015 1139.175 1924.345 1139.505 ;
        RECT 1924.030 1138.145 1924.330 1139.175 ;
        RECT 1924.950 1138.145 1925.250 1140.535 ;
        RECT 1924.015 1137.815 1924.345 1138.145 ;
        RECT 1924.935 1137.815 1925.265 1138.145 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2186.910 1374.520 2187.230 1374.580 ;
        RECT 2221.410 1374.520 2221.730 1374.580 ;
        RECT 2186.910 1374.380 2221.730 1374.520 ;
        RECT 2186.910 1374.320 2187.230 1374.380 ;
        RECT 2221.410 1374.320 2221.730 1374.380 ;
        RECT 1799.130 1374.180 1799.450 1374.240 ;
        RECT 1801.890 1374.180 1802.210 1374.240 ;
        RECT 1799.130 1374.040 1802.210 1374.180 ;
        RECT 1799.130 1373.980 1799.450 1374.040 ;
        RECT 1801.890 1373.980 1802.210 1374.040 ;
        RECT 1932.070 1374.180 1932.390 1374.240 ;
        RECT 1970.250 1374.180 1970.570 1374.240 ;
        RECT 1932.070 1374.040 1970.570 1374.180 ;
        RECT 1932.070 1373.980 1932.390 1374.040 ;
        RECT 1970.250 1373.980 1970.570 1374.040 ;
        RECT 2456.470 1374.180 2456.790 1374.240 ;
        RECT 2504.310 1374.180 2504.630 1374.240 ;
        RECT 2456.470 1374.040 2504.630 1374.180 ;
        RECT 2456.470 1373.980 2456.790 1374.040 ;
        RECT 2504.310 1373.980 2504.630 1374.040 ;
        RECT 2621.610 1373.840 2621.930 1373.900 ;
        RECT 2622.530 1373.840 2622.850 1373.900 ;
        RECT 2621.610 1373.700 2622.850 1373.840 ;
        RECT 2621.610 1373.640 2621.930 1373.700 ;
        RECT 2622.530 1373.640 2622.850 1373.700 ;
        RECT 1642.270 1373.500 1642.590 1373.560 ;
        RECT 1690.110 1373.500 1690.430 1373.560 ;
        RECT 1642.270 1373.360 1690.430 1373.500 ;
        RECT 1642.270 1373.300 1642.590 1373.360 ;
        RECT 1690.110 1373.300 1690.430 1373.360 ;
        RECT 2649.670 1373.500 2649.990 1373.560 ;
        RECT 2697.510 1373.500 2697.830 1373.560 ;
        RECT 2649.670 1373.360 2697.830 1373.500 ;
        RECT 2649.670 1373.300 2649.990 1373.360 ;
        RECT 2697.510 1373.300 2697.830 1373.360 ;
      LAYER via ;
        RECT 2186.940 1374.320 2187.200 1374.580 ;
        RECT 2221.440 1374.320 2221.700 1374.580 ;
        RECT 1799.160 1373.980 1799.420 1374.240 ;
        RECT 1801.920 1373.980 1802.180 1374.240 ;
        RECT 1932.100 1373.980 1932.360 1374.240 ;
        RECT 1970.280 1373.980 1970.540 1374.240 ;
        RECT 2456.500 1373.980 2456.760 1374.240 ;
        RECT 2504.340 1373.980 2504.600 1374.240 ;
        RECT 2621.640 1373.640 2621.900 1373.900 ;
        RECT 2622.560 1373.640 2622.820 1373.900 ;
        RECT 1642.300 1373.300 1642.560 1373.560 ;
        RECT 1690.140 1373.300 1690.400 1373.560 ;
        RECT 2649.700 1373.300 2649.960 1373.560 ;
        RECT 2697.540 1373.300 2697.800 1373.560 ;
      LAYER met2 ;
        RECT 1256.350 2498.050 1256.630 2500.000 ;
        RECT 1258.190 2498.050 1258.470 2498.165 ;
        RECT 1256.350 2497.910 1258.470 2498.050 ;
        RECT 1256.350 2496.000 1256.630 2497.910 ;
        RECT 1258.190 2497.795 1258.470 2497.910 ;
        RECT 1562.710 1375.795 1562.990 1376.165 ;
        RECT 1562.780 1374.805 1562.920 1375.795 ;
        RECT 1970.270 1375.115 1970.550 1375.485 ;
        RECT 1562.710 1374.435 1562.990 1374.805 ;
        RECT 1690.130 1374.435 1690.410 1374.805 ;
        RECT 1424.710 1373.755 1424.990 1374.125 ;
        RECT 1606.410 1373.755 1606.690 1374.125 ;
        RECT 1424.780 1372.765 1424.920 1373.755 ;
        RECT 1424.710 1372.395 1424.990 1372.765 ;
        RECT 1606.480 1372.085 1606.620 1373.755 ;
        RECT 1690.200 1373.590 1690.340 1374.435 ;
        RECT 1970.340 1374.270 1970.480 1375.115 ;
        RECT 2186.930 1374.435 2187.210 1374.805 ;
        RECT 2221.430 1374.435 2221.710 1374.805 ;
        RECT 2304.230 1374.435 2304.510 1374.805 ;
        RECT 2504.330 1374.435 2504.610 1374.805 ;
        RECT 2697.530 1374.435 2697.810 1374.805 ;
        RECT 2186.940 1374.290 2187.200 1374.435 ;
        RECT 2221.440 1374.290 2221.700 1374.435 ;
        RECT 1799.160 1374.125 1799.420 1374.270 ;
        RECT 1801.920 1374.125 1802.180 1374.270 ;
        RECT 1932.100 1374.125 1932.360 1374.270 ;
        RECT 1799.150 1373.755 1799.430 1374.125 ;
        RECT 1801.910 1373.755 1802.190 1374.125 ;
        RECT 1932.090 1373.755 1932.370 1374.125 ;
        RECT 1970.280 1373.950 1970.540 1374.270 ;
        RECT 1993.730 1374.010 1994.010 1374.125 ;
        RECT 1994.650 1374.010 1994.930 1374.125 ;
        RECT 1993.730 1373.870 1994.930 1374.010 ;
        RECT 1993.730 1373.755 1994.010 1373.870 ;
        RECT 1994.650 1373.755 1994.930 1373.870 ;
        RECT 1642.300 1373.445 1642.560 1373.590 ;
        RECT 1642.290 1373.075 1642.570 1373.445 ;
        RECT 1690.140 1373.270 1690.400 1373.590 ;
        RECT 2304.300 1372.765 2304.440 1374.435 ;
        RECT 2504.400 1374.270 2504.540 1374.435 ;
        RECT 2456.500 1374.125 2456.760 1374.270 ;
        RECT 2456.490 1373.755 2456.770 1374.125 ;
        RECT 2504.340 1373.950 2504.600 1374.270 ;
        RECT 2574.250 1374.010 2574.530 1374.125 ;
        RECT 2573.400 1373.870 2574.530 1374.010 ;
        RECT 2573.400 1373.445 2573.540 1373.870 ;
        RECT 2574.250 1373.755 2574.530 1373.870 ;
        RECT 2621.630 1373.755 2621.910 1374.125 ;
        RECT 2621.640 1373.610 2621.900 1373.755 ;
        RECT 2622.560 1373.610 2622.820 1373.930 ;
        RECT 2622.620 1373.445 2622.760 1373.610 ;
        RECT 2697.600 1373.590 2697.740 1374.435 ;
        RECT 2649.700 1373.445 2649.960 1373.590 ;
        RECT 2573.330 1373.075 2573.610 1373.445 ;
        RECT 2622.550 1373.075 2622.830 1373.445 ;
        RECT 2649.690 1373.075 2649.970 1373.445 ;
        RECT 2697.540 1373.270 2697.800 1373.590 ;
        RECT 2304.230 1372.395 2304.510 1372.765 ;
        RECT 1606.410 1371.715 1606.690 1372.085 ;
      LAYER via2 ;
        RECT 1258.190 2497.840 1258.470 2498.120 ;
        RECT 1562.710 1375.840 1562.990 1376.120 ;
        RECT 1970.270 1375.160 1970.550 1375.440 ;
        RECT 1562.710 1374.480 1562.990 1374.760 ;
        RECT 1690.130 1374.480 1690.410 1374.760 ;
        RECT 1424.710 1373.800 1424.990 1374.080 ;
        RECT 1606.410 1373.800 1606.690 1374.080 ;
        RECT 1424.710 1372.440 1424.990 1372.720 ;
        RECT 2186.930 1374.480 2187.210 1374.760 ;
        RECT 2221.430 1374.480 2221.710 1374.760 ;
        RECT 2304.230 1374.480 2304.510 1374.760 ;
        RECT 2504.330 1374.480 2504.610 1374.760 ;
        RECT 2697.530 1374.480 2697.810 1374.760 ;
        RECT 1799.150 1373.800 1799.430 1374.080 ;
        RECT 1801.910 1373.800 1802.190 1374.080 ;
        RECT 1932.090 1373.800 1932.370 1374.080 ;
        RECT 1993.730 1373.800 1994.010 1374.080 ;
        RECT 1994.650 1373.800 1994.930 1374.080 ;
        RECT 1642.290 1373.120 1642.570 1373.400 ;
        RECT 2456.490 1373.800 2456.770 1374.080 ;
        RECT 2574.250 1373.800 2574.530 1374.080 ;
        RECT 2621.630 1373.800 2621.910 1374.080 ;
        RECT 2573.330 1373.120 2573.610 1373.400 ;
        RECT 2622.550 1373.120 2622.830 1373.400 ;
        RECT 2649.690 1373.120 2649.970 1373.400 ;
        RECT 2304.230 1372.440 2304.510 1372.720 ;
        RECT 1606.410 1371.760 1606.690 1372.040 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1378.100 2924.800 1379.300 ;
=======
        RECT 1260.005 2498.130 1260.335 2498.145 ;
=======
        RECT 1258.165 2498.130 1258.495 2498.145 ;
>>>>>>> re-updated local openlane
        RECT 1261.590 2498.130 1261.970 2498.140 ;
        RECT 1258.165 2497.830 1261.970 2498.130 ;
        RECT 1258.165 2497.815 1258.495 2497.830 ;
        RECT 1261.590 2497.820 1261.970 2497.830 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2916.710 1378.550 2924.800 1378.850 ;
        RECT 1538.510 1376.130 1538.890 1376.140 ;
        RECT 1562.685 1376.130 1563.015 1376.145 ;
        RECT 1538.510 1375.830 1563.015 1376.130 ;
        RECT 1538.510 1375.820 1538.890 1375.830 ;
        RECT 1562.685 1375.815 1563.015 1375.830 ;
        RECT 1261.590 1375.450 1261.970 1375.460 ;
        RECT 1970.245 1375.450 1970.575 1375.465 ;
        RECT 1980.110 1375.450 1980.490 1375.460 ;
        RECT 1261.590 1375.150 1270.210 1375.450 ;
        RECT 1261.590 1375.140 1261.970 1375.150 ;
        RECT 1269.910 1374.770 1270.210 1375.150 ;
        RECT 1970.245 1375.150 1980.490 1375.450 ;
        RECT 1970.245 1375.135 1970.575 1375.150 ;
        RECT 1980.110 1375.140 1980.490 1375.150 ;
        RECT 1303.910 1374.770 1304.290 1374.780 ;
        RECT 1441.910 1374.770 1442.290 1374.780 ;
        RECT 1538.510 1374.770 1538.890 1374.780 ;
        RECT 1269.910 1374.470 1304.290 1374.770 ;
        RECT 1303.910 1374.460 1304.290 1374.470 ;
        RECT 1352.710 1374.470 1377.850 1374.770 ;
        RECT 1352.710 1374.090 1353.010 1374.470 ;
        RECT 1304.870 1373.790 1353.010 1374.090 ;
        RECT 1377.550 1374.090 1377.850 1374.470 ;
        RECT 1441.910 1374.470 1538.890 1374.770 ;
        RECT 1441.910 1374.460 1442.290 1374.470 ;
        RECT 1538.510 1374.460 1538.890 1374.470 ;
        RECT 1562.685 1374.770 1563.015 1374.785 ;
        RECT 1690.105 1374.770 1690.435 1374.785 ;
        RECT 1883.510 1374.770 1883.890 1374.780 ;
        RECT 2186.905 1374.770 2187.235 1374.785 ;
        RECT 1562.685 1374.470 1586.690 1374.770 ;
        RECT 1562.685 1374.455 1563.015 1374.470 ;
        RECT 1424.685 1374.090 1425.015 1374.105 ;
        RECT 1377.550 1373.790 1425.015 1374.090 ;
        RECT 1586.390 1374.090 1586.690 1374.470 ;
        RECT 1690.105 1374.470 1704.450 1374.770 ;
        RECT 1690.105 1374.455 1690.435 1374.470 ;
        RECT 1606.385 1374.090 1606.715 1374.105 ;
        RECT 1586.390 1373.790 1606.715 1374.090 ;
        RECT 1303.910 1373.410 1304.290 1373.420 ;
        RECT 1304.870 1373.410 1305.170 1373.790 ;
        RECT 1424.685 1373.775 1425.015 1373.790 ;
        RECT 1606.385 1373.775 1606.715 1373.790 ;
        RECT 1642.265 1373.410 1642.595 1373.425 ;
        RECT 1303.910 1373.110 1305.170 1373.410 ;
        RECT 1641.590 1373.110 1642.595 1373.410 ;
        RECT 1704.150 1373.410 1704.450 1374.470 ;
        RECT 1849.510 1374.470 1883.890 1374.770 ;
        RECT 1799.125 1374.090 1799.455 1374.105 ;
        RECT 1752.910 1373.790 1799.455 1374.090 ;
        RECT 1752.910 1373.410 1753.210 1373.790 ;
        RECT 1799.125 1373.775 1799.455 1373.790 ;
        RECT 1801.885 1374.090 1802.215 1374.105 ;
        RECT 1801.885 1373.790 1835.090 1374.090 ;
        RECT 1801.885 1373.775 1802.215 1373.790 ;
        RECT 1704.150 1373.110 1753.210 1373.410 ;
        RECT 1834.790 1373.410 1835.090 1373.790 ;
        RECT 1849.510 1373.410 1849.810 1374.470 ;
        RECT 1883.510 1374.460 1883.890 1374.470 ;
        RECT 2062.950 1374.470 2111.090 1374.770 ;
        RECT 1932.065 1374.090 1932.395 1374.105 ;
        RECT 1834.790 1373.110 1849.810 1373.410 ;
        RECT 1931.390 1373.790 1932.395 1374.090 ;
        RECT 1303.910 1373.100 1304.290 1373.110 ;
        RECT 1424.685 1372.730 1425.015 1372.745 ;
        RECT 1441.910 1372.730 1442.290 1372.740 ;
        RECT 1424.685 1372.430 1442.290 1372.730 ;
        RECT 1424.685 1372.415 1425.015 1372.430 ;
        RECT 1441.910 1372.420 1442.290 1372.430 ;
        RECT 1606.385 1372.050 1606.715 1372.065 ;
        RECT 1641.590 1372.050 1641.890 1373.110 ;
        RECT 1642.265 1373.095 1642.595 1373.110 ;
        RECT 1883.510 1372.730 1883.890 1372.740 ;
        RECT 1931.390 1372.730 1931.690 1373.790 ;
        RECT 1932.065 1373.775 1932.395 1373.790 ;
        RECT 1980.110 1374.090 1980.490 1374.100 ;
        RECT 1993.705 1374.090 1994.035 1374.105 ;
        RECT 1980.110 1373.790 1994.035 1374.090 ;
        RECT 1980.110 1373.780 1980.490 1373.790 ;
        RECT 1993.705 1373.775 1994.035 1373.790 ;
        RECT 1994.625 1374.090 1994.955 1374.105 ;
        RECT 1994.625 1373.790 2042.090 1374.090 ;
        RECT 1994.625 1373.775 1994.955 1373.790 ;
        RECT 2041.790 1373.410 2042.090 1373.790 ;
        RECT 2062.950 1373.410 2063.250 1374.470 ;
        RECT 2041.790 1373.110 2063.250 1373.410 ;
        RECT 2110.790 1373.410 2111.090 1374.470 ;
        RECT 2111.710 1374.470 2187.235 1374.770 ;
        RECT 2111.710 1373.410 2112.010 1374.470 ;
        RECT 2186.905 1374.455 2187.235 1374.470 ;
        RECT 2221.405 1374.770 2221.735 1374.785 ;
        RECT 2304.205 1374.770 2304.535 1374.785 ;
        RECT 2504.305 1374.770 2504.635 1374.785 ;
        RECT 2697.505 1374.770 2697.835 1374.785 ;
        RECT 2221.405 1374.470 2235.290 1374.770 ;
        RECT 2221.405 1374.455 2221.735 1374.470 ;
        RECT 2110.790 1373.110 2112.010 1373.410 ;
        RECT 2234.990 1373.410 2235.290 1374.470 ;
        RECT 2304.205 1374.470 2353.050 1374.770 ;
        RECT 2304.205 1374.455 2304.535 1374.470 ;
        RECT 2269.910 1374.090 2270.290 1374.100 ;
        RECT 2235.910 1373.790 2270.290 1374.090 ;
        RECT 2352.750 1374.090 2353.050 1374.470 ;
        RECT 2401.510 1374.470 2429.410 1374.770 ;
        RECT 2352.750 1373.790 2400.890 1374.090 ;
        RECT 2235.910 1373.410 2236.210 1373.790 ;
        RECT 2269.910 1373.780 2270.290 1373.790 ;
        RECT 2234.990 1373.110 2236.210 1373.410 ;
        RECT 2400.590 1373.410 2400.890 1373.790 ;
        RECT 2401.510 1373.410 2401.810 1374.470 ;
        RECT 2429.110 1374.090 2429.410 1374.470 ;
        RECT 2504.305 1374.470 2526.010 1374.770 ;
        RECT 2504.305 1374.455 2504.635 1374.470 ;
        RECT 2456.465 1374.090 2456.795 1374.105 ;
        RECT 2429.110 1373.790 2456.795 1374.090 ;
        RECT 2456.465 1373.775 2456.795 1373.790 ;
        RECT 2400.590 1373.110 2401.810 1373.410 ;
        RECT 2525.710 1373.410 2526.010 1374.470 ;
        RECT 2697.505 1374.470 2739.450 1374.770 ;
        RECT 2697.505 1374.455 2697.835 1374.470 ;
        RECT 2574.225 1374.090 2574.555 1374.105 ;
        RECT 2621.605 1374.090 2621.935 1374.105 ;
        RECT 2574.225 1373.790 2621.935 1374.090 ;
        RECT 2739.150 1374.090 2739.450 1374.470 ;
        RECT 2787.910 1374.470 2836.050 1374.770 ;
        RECT 2739.150 1373.790 2787.290 1374.090 ;
        RECT 2574.225 1373.775 2574.555 1373.790 ;
        RECT 2621.605 1373.775 2621.935 1373.790 ;
        RECT 2573.305 1373.410 2573.635 1373.425 ;
        RECT 2525.710 1373.110 2573.635 1373.410 ;
        RECT 2573.305 1373.095 2573.635 1373.110 ;
        RECT 2622.525 1373.410 2622.855 1373.425 ;
        RECT 2649.665 1373.410 2649.995 1373.425 ;
        RECT 2622.525 1373.110 2649.995 1373.410 ;
        RECT 2786.990 1373.410 2787.290 1373.790 ;
        RECT 2787.910 1373.410 2788.210 1374.470 ;
        RECT 2835.750 1374.090 2836.050 1374.470 ;
        RECT 2916.710 1374.090 2917.010 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 2835.750 1373.790 2883.890 1374.090 ;
        RECT 2786.990 1373.110 2788.210 1373.410 ;
        RECT 2883.590 1373.410 2883.890 1373.790 ;
        RECT 2884.510 1373.790 2917.010 1374.090 ;
        RECT 2884.510 1373.410 2884.810 1373.790 ;
        RECT 2883.590 1373.110 2884.810 1373.410 ;
        RECT 2622.525 1373.095 2622.855 1373.110 ;
        RECT 2649.665 1373.095 2649.995 1373.110 ;
        RECT 1883.510 1372.430 1931.690 1372.730 ;
        RECT 2269.910 1372.730 2270.290 1372.740 ;
        RECT 2304.205 1372.730 2304.535 1372.745 ;
        RECT 2269.910 1372.430 2304.535 1372.730 ;
        RECT 1883.510 1372.420 1883.890 1372.430 ;
        RECT 2269.910 1372.420 2270.290 1372.430 ;
        RECT 2304.205 1372.415 2304.535 1372.430 ;
        RECT 1606.385 1371.750 1641.890 1372.050 ;
        RECT 1606.385 1371.735 1606.715 1371.750 ;
      LAYER via3 ;
        RECT 1261.620 2497.820 1261.940 2498.140 ;
        RECT 1538.540 1375.820 1538.860 1376.140 ;
        RECT 1261.620 1375.140 1261.940 1375.460 ;
        RECT 1980.140 1375.140 1980.460 1375.460 ;
        RECT 1303.940 1374.460 1304.260 1374.780 ;
        RECT 1441.940 1374.460 1442.260 1374.780 ;
        RECT 1538.540 1374.460 1538.860 1374.780 ;
        RECT 1303.940 1373.100 1304.260 1373.420 ;
        RECT 1883.540 1374.460 1883.860 1374.780 ;
        RECT 1441.940 1372.420 1442.260 1372.740 ;
        RECT 1883.540 1372.420 1883.860 1372.740 ;
        RECT 1980.140 1373.780 1980.460 1374.100 ;
        RECT 2269.940 1373.780 2270.260 1374.100 ;
        RECT 2269.940 1372.420 2270.260 1372.740 ;
      LAYER met4 ;
        RECT 1261.615 2497.815 1261.945 2498.145 ;
        RECT 1261.630 1375.465 1261.930 2497.815 ;
        RECT 1538.535 1375.815 1538.865 1376.145 ;
        RECT 1261.615 1375.135 1261.945 1375.465 ;
        RECT 1538.550 1374.785 1538.850 1375.815 ;
        RECT 1980.135 1375.135 1980.465 1375.465 ;
        RECT 1303.935 1374.455 1304.265 1374.785 ;
        RECT 1441.935 1374.455 1442.265 1374.785 ;
<<<<<<< HEAD
        RECT 1980.135 1374.455 1980.465 1374.785 ;
        RECT 1386.735 1373.775 1387.065 1374.105 ;
        RECT 1441.950 1373.425 1442.250 1374.455 ;
        RECT 1331.535 1373.095 1331.865 1373.425 ;
        RECT 1441.935 1373.095 1442.265 1373.425 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1538.535 1374.455 1538.865 1374.785 ;
        RECT 1883.535 1374.455 1883.865 1374.785 ;
        RECT 1303.950 1373.425 1304.250 1374.455 ;
        RECT 1303.935 1373.095 1304.265 1373.425 ;
        RECT 1441.950 1372.745 1442.250 1374.455 ;
        RECT 1883.550 1372.745 1883.850 1374.455 ;
        RECT 1980.150 1374.105 1980.450 1375.135 ;
        RECT 1980.135 1373.775 1980.465 1374.105 ;
        RECT 2269.935 1373.775 2270.265 1374.105 ;
        RECT 2269.950 1372.745 2270.250 1373.775 ;
        RECT 1441.935 1372.415 1442.265 1372.745 ;
        RECT 1883.535 1372.415 1883.865 1372.745 ;
        RECT 2269.935 1372.415 2270.265 1372.745 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1497.370 1609.120 1497.690 1609.180 ;
        RECT 1562.690 1609.120 1563.010 1609.180 ;
        RECT 1497.370 1608.980 1563.010 1609.120 ;
        RECT 1497.370 1608.920 1497.690 1608.980 ;
        RECT 1562.690 1608.920 1563.010 1608.980 ;
        RECT 1642.270 1608.100 1642.590 1608.160 ;
        RECT 1690.110 1608.100 1690.430 1608.160 ;
        RECT 1642.270 1607.960 1690.430 1608.100 ;
        RECT 1642.270 1607.900 1642.590 1607.960 ;
        RECT 1690.110 1607.900 1690.430 1607.960 ;
        RECT 1738.870 1608.100 1739.190 1608.160 ;
        RECT 1753.590 1608.100 1753.910 1608.160 ;
        RECT 1738.870 1607.960 1753.910 1608.100 ;
        RECT 1738.870 1607.900 1739.190 1607.960 ;
        RECT 1753.590 1607.900 1753.910 1607.960 ;
      LAYER via ;
        RECT 1497.400 1608.920 1497.660 1609.180 ;
        RECT 1562.720 1608.920 1562.980 1609.180 ;
        RECT 1642.300 1607.900 1642.560 1608.160 ;
        RECT 1690.140 1607.900 1690.400 1608.160 ;
        RECT 1738.900 1607.900 1739.160 1608.160 ;
        RECT 1753.620 1607.900 1753.880 1608.160 ;
      LAYER met2 ;
        RECT 1275.210 2496.690 1275.490 2496.805 ;
        RECT 1275.670 2496.690 1275.950 2500.000 ;
        RECT 1275.210 2496.550 1275.950 2496.690 ;
        RECT 1275.210 2496.435 1275.490 2496.550 ;
        RECT 1275.670 2496.000 1275.950 2496.550 ;
        RECT 1328.110 1610.395 1328.390 1610.765 ;
        RECT 1328.180 1608.725 1328.320 1610.395 ;
        RECT 1483.130 1609.035 1483.410 1609.405 ;
        RECT 1497.390 1609.035 1497.670 1609.405 ;
        RECT 1483.200 1608.725 1483.340 1609.035 ;
        RECT 1497.400 1608.890 1497.660 1609.035 ;
        RECT 1562.720 1608.890 1562.980 1609.210 ;
        RECT 1690.130 1609.035 1690.410 1609.405 ;
        RECT 1994.650 1609.035 1994.930 1609.405 ;
        RECT 2091.250 1609.035 2091.530 1609.405 ;
        RECT 2186.930 1609.290 2187.210 1609.405 ;
        RECT 2187.850 1609.290 2188.130 1609.405 ;
        RECT 2186.930 1609.150 2188.130 1609.290 ;
        RECT 2186.930 1609.035 2187.210 1609.150 ;
        RECT 2187.850 1609.035 2188.130 1609.150 ;
        RECT 2283.530 1609.290 2283.810 1609.405 ;
        RECT 2284.450 1609.290 2284.730 1609.405 ;
        RECT 2283.530 1609.150 2284.730 1609.290 ;
        RECT 2283.530 1609.035 2283.810 1609.150 ;
        RECT 2284.450 1609.035 2284.730 1609.150 ;
        RECT 2380.130 1609.290 2380.410 1609.405 ;
        RECT 2381.050 1609.290 2381.330 1609.405 ;
        RECT 2380.130 1609.150 2381.330 1609.290 ;
        RECT 2380.130 1609.035 2380.410 1609.150 ;
        RECT 2381.050 1609.035 2381.330 1609.150 ;
        RECT 2573.330 1609.035 2573.610 1609.405 ;
        RECT 1562.780 1608.725 1562.920 1608.890 ;
        RECT 1328.110 1608.355 1328.390 1608.725 ;
        RECT 1483.130 1608.355 1483.410 1608.725 ;
        RECT 1562.710 1608.355 1562.990 1608.725 ;
        RECT 1606.410 1608.355 1606.690 1608.725 ;
        RECT 1606.480 1606.685 1606.620 1608.355 ;
        RECT 1690.200 1608.190 1690.340 1609.035 ;
        RECT 1753.610 1608.355 1753.890 1608.725 ;
        RECT 1835.490 1608.355 1835.770 1608.725 ;
        RECT 1993.730 1608.610 1994.010 1608.725 ;
        RECT 1994.720 1608.610 1994.860 1609.035 ;
        RECT 1993.730 1608.470 1994.860 1608.610 ;
        RECT 2090.330 1608.610 2090.610 1608.725 ;
        RECT 2091.320 1608.610 2091.460 1609.035 ;
        RECT 2090.330 1608.470 2091.460 1608.610 ;
        RECT 2524.570 1608.610 2524.850 1608.725 ;
        RECT 2525.950 1608.610 2526.230 1608.725 ;
        RECT 2524.570 1608.470 2526.230 1608.610 ;
        RECT 2573.400 1608.610 2573.540 1609.035 ;
        RECT 2573.790 1608.610 2574.070 1608.725 ;
        RECT 2573.400 1608.470 2574.070 1608.610 ;
        RECT 1993.730 1608.355 1994.010 1608.470 ;
        RECT 2090.330 1608.355 2090.610 1608.470 ;
        RECT 2524.570 1608.355 2524.850 1608.470 ;
        RECT 2525.950 1608.355 2526.230 1608.470 ;
        RECT 2573.790 1608.355 2574.070 1608.470 ;
        RECT 1753.680 1608.190 1753.820 1608.355 ;
        RECT 1642.300 1608.045 1642.560 1608.190 ;
        RECT 1642.290 1607.675 1642.570 1608.045 ;
        RECT 1690.140 1607.870 1690.400 1608.190 ;
        RECT 1738.900 1608.045 1739.160 1608.190 ;
        RECT 1738.890 1607.675 1739.170 1608.045 ;
        RECT 1753.620 1607.870 1753.880 1608.190 ;
        RECT 1835.560 1606.685 1835.700 1608.355 ;
        RECT 1606.410 1606.315 1606.690 1606.685 ;
        RECT 1835.490 1606.315 1835.770 1606.685 ;
      LAYER via2 ;
        RECT 1275.210 2496.480 1275.490 2496.760 ;
        RECT 1328.110 1610.440 1328.390 1610.720 ;
        RECT 1483.130 1609.080 1483.410 1609.360 ;
        RECT 1497.390 1609.080 1497.670 1609.360 ;
        RECT 1690.130 1609.080 1690.410 1609.360 ;
        RECT 1994.650 1609.080 1994.930 1609.360 ;
        RECT 2091.250 1609.080 2091.530 1609.360 ;
        RECT 2186.930 1609.080 2187.210 1609.360 ;
        RECT 2187.850 1609.080 2188.130 1609.360 ;
        RECT 2283.530 1609.080 2283.810 1609.360 ;
        RECT 2284.450 1609.080 2284.730 1609.360 ;
        RECT 2380.130 1609.080 2380.410 1609.360 ;
        RECT 2381.050 1609.080 2381.330 1609.360 ;
        RECT 2573.330 1609.080 2573.610 1609.360 ;
        RECT 1328.110 1608.400 1328.390 1608.680 ;
        RECT 1483.130 1608.400 1483.410 1608.680 ;
        RECT 1562.710 1608.400 1562.990 1608.680 ;
        RECT 1606.410 1608.400 1606.690 1608.680 ;
        RECT 1753.610 1608.400 1753.890 1608.680 ;
        RECT 1835.490 1608.400 1835.770 1608.680 ;
        RECT 1993.730 1608.400 1994.010 1608.680 ;
        RECT 2090.330 1608.400 2090.610 1608.680 ;
        RECT 2524.570 1608.400 2524.850 1608.680 ;
        RECT 2525.950 1608.400 2526.230 1608.680 ;
        RECT 2573.790 1608.400 2574.070 1608.680 ;
        RECT 1642.290 1607.720 1642.570 1608.000 ;
        RECT 1738.890 1607.720 1739.170 1608.000 ;
        RECT 1606.410 1606.360 1606.690 1606.640 ;
        RECT 1835.490 1606.360 1835.770 1606.640 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1612.700 2924.800 1613.900 ;
=======
        RECT 1280.245 2498.130 1280.575 2498.145 ;
        RECT 1280.910 2498.130 1281.290 2498.140 ;
        RECT 1280.245 2497.830 1281.290 2498.130 ;
        RECT 1280.245 2497.815 1280.575 2497.830 ;
        RECT 1280.910 2497.820 1281.290 2497.830 ;
=======
        RECT 1275.185 2496.780 1275.515 2496.785 ;
        RECT 1275.185 2496.770 1275.770 2496.780 ;
        RECT 1275.185 2496.470 1275.970 2496.770 ;
        RECT 1275.185 2496.460 1275.770 2496.470 ;
        RECT 1275.185 2496.455 1275.515 2496.460 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2916.710 1613.150 2924.800 1613.450 ;
        RECT 1275.390 1610.730 1275.770 1610.740 ;
        RECT 1328.085 1610.730 1328.415 1610.745 ;
        RECT 1275.390 1610.430 1328.415 1610.730 ;
        RECT 1275.390 1610.420 1275.770 1610.430 ;
        RECT 1328.085 1610.415 1328.415 1610.430 ;
        RECT 1483.105 1609.370 1483.435 1609.385 ;
        RECT 1497.365 1609.370 1497.695 1609.385 ;
        RECT 1483.105 1609.070 1497.695 1609.370 ;
        RECT 1483.105 1609.055 1483.435 1609.070 ;
        RECT 1497.365 1609.055 1497.695 1609.070 ;
        RECT 1690.105 1609.370 1690.435 1609.385 ;
        RECT 1994.625 1609.370 1994.955 1609.385 ;
        RECT 2091.225 1609.370 2091.555 1609.385 ;
        RECT 2186.905 1609.370 2187.235 1609.385 ;
        RECT 1690.105 1609.070 1704.450 1609.370 ;
        RECT 1690.105 1609.055 1690.435 1609.070 ;
        RECT 1328.085 1608.690 1328.415 1608.705 ;
        RECT 1338.870 1608.690 1339.250 1608.700 ;
        RECT 1483.105 1608.690 1483.435 1608.705 ;
        RECT 1328.085 1608.390 1339.250 1608.690 ;
        RECT 1328.085 1608.375 1328.415 1608.390 ;
        RECT 1338.870 1608.380 1339.250 1608.390 ;
        RECT 1441.030 1608.390 1483.435 1608.690 ;
        RECT 1441.030 1608.010 1441.330 1608.390 ;
        RECT 1483.105 1608.375 1483.435 1608.390 ;
        RECT 1562.685 1608.690 1563.015 1608.705 ;
        RECT 1606.385 1608.690 1606.715 1608.705 ;
        RECT 1562.685 1608.390 1606.715 1608.690 ;
        RECT 1562.685 1608.375 1563.015 1608.390 ;
        RECT 1606.385 1608.375 1606.715 1608.390 ;
        RECT 1642.265 1608.010 1642.595 1608.025 ;
        RECT 1394.110 1607.710 1441.330 1608.010 ;
        RECT 1641.590 1607.710 1642.595 1608.010 ;
        RECT 1704.150 1608.010 1704.450 1609.070 ;
        RECT 1994.625 1609.070 2043.010 1609.370 ;
        RECT 1994.625 1609.055 1994.955 1609.070 ;
        RECT 1753.585 1608.690 1753.915 1608.705 ;
        RECT 1835.465 1608.690 1835.795 1608.705 ;
        RECT 1753.585 1608.390 1835.795 1608.690 ;
        RECT 1753.585 1608.375 1753.915 1608.390 ;
        RECT 1835.465 1608.375 1835.795 1608.390 ;
        RECT 1882.590 1608.690 1882.970 1608.700 ;
        RECT 1993.705 1608.690 1994.035 1608.705 ;
        RECT 1882.590 1608.390 1896.730 1608.690 ;
        RECT 1882.590 1608.380 1882.970 1608.390 ;
        RECT 1738.865 1608.010 1739.195 1608.025 ;
        RECT 1704.150 1607.710 1739.195 1608.010 ;
        RECT 1394.110 1606.650 1394.410 1607.710 ;
        RECT 1386.750 1606.350 1394.410 1606.650 ;
        RECT 1606.385 1606.650 1606.715 1606.665 ;
        RECT 1641.590 1606.650 1641.890 1607.710 ;
        RECT 1642.265 1607.695 1642.595 1607.710 ;
        RECT 1738.865 1607.695 1739.195 1607.710 ;
        RECT 1896.430 1607.330 1896.730 1608.390 ;
        RECT 1898.270 1608.390 1994.035 1608.690 ;
        RECT 2042.710 1608.690 2043.010 1609.070 ;
        RECT 2091.225 1609.070 2139.610 1609.370 ;
        RECT 2091.225 1609.055 2091.555 1609.070 ;
        RECT 2090.305 1608.690 2090.635 1608.705 ;
        RECT 2042.710 1608.390 2090.635 1608.690 ;
        RECT 2139.310 1608.690 2139.610 1609.070 ;
        RECT 2185.310 1609.070 2187.235 1609.370 ;
        RECT 2185.310 1608.690 2185.610 1609.070 ;
        RECT 2186.905 1609.055 2187.235 1609.070 ;
        RECT 2187.825 1609.370 2188.155 1609.385 ;
        RECT 2283.505 1609.370 2283.835 1609.385 ;
        RECT 2187.825 1609.070 2236.210 1609.370 ;
        RECT 2187.825 1609.055 2188.155 1609.070 ;
        RECT 2139.310 1608.390 2185.610 1608.690 ;
        RECT 2235.910 1608.690 2236.210 1609.070 ;
        RECT 2281.910 1609.070 2283.835 1609.370 ;
        RECT 2281.910 1608.690 2282.210 1609.070 ;
        RECT 2283.505 1609.055 2283.835 1609.070 ;
        RECT 2284.425 1609.370 2284.755 1609.385 ;
        RECT 2380.105 1609.370 2380.435 1609.385 ;
        RECT 2284.425 1609.070 2332.810 1609.370 ;
        RECT 2284.425 1609.055 2284.755 1609.070 ;
        RECT 2235.910 1608.390 2282.210 1608.690 ;
        RECT 2332.510 1608.690 2332.810 1609.070 ;
        RECT 2378.510 1609.070 2380.435 1609.370 ;
        RECT 2378.510 1608.690 2378.810 1609.070 ;
        RECT 2380.105 1609.055 2380.435 1609.070 ;
        RECT 2381.025 1609.370 2381.355 1609.385 ;
        RECT 2573.305 1609.370 2573.635 1609.385 ;
        RECT 2381.025 1609.070 2477.250 1609.370 ;
        RECT 2381.025 1609.055 2381.355 1609.070 ;
        RECT 2332.510 1608.390 2378.810 1608.690 ;
        RECT 2476.950 1608.690 2477.250 1609.070 ;
        RECT 2559.750 1609.070 2573.635 1609.370 ;
        RECT 2524.545 1608.690 2524.875 1608.705 ;
        RECT 2476.950 1608.390 2524.875 1608.690 ;
        RECT 1898.270 1607.330 1898.570 1608.390 ;
        RECT 1993.705 1608.375 1994.035 1608.390 ;
        RECT 2090.305 1608.375 2090.635 1608.390 ;
        RECT 2524.545 1608.375 2524.875 1608.390 ;
        RECT 2525.925 1608.690 2526.255 1608.705 ;
        RECT 2559.750 1608.690 2560.050 1609.070 ;
        RECT 2573.305 1609.055 2573.635 1609.070 ;
        RECT 2594.710 1609.070 2642.850 1609.370 ;
        RECT 2525.925 1608.390 2560.050 1608.690 ;
        RECT 2573.765 1608.690 2574.095 1608.705 ;
        RECT 2594.710 1608.690 2595.010 1609.070 ;
        RECT 2573.765 1608.390 2595.010 1608.690 ;
        RECT 2642.550 1608.690 2642.850 1609.070 ;
        RECT 2691.310 1609.070 2739.450 1609.370 ;
        RECT 2642.550 1608.390 2690.690 1608.690 ;
        RECT 2525.925 1608.375 2526.255 1608.390 ;
        RECT 2573.765 1608.375 2574.095 1608.390 ;
        RECT 2690.390 1608.010 2690.690 1608.390 ;
        RECT 2691.310 1608.010 2691.610 1609.070 ;
        RECT 2739.150 1608.690 2739.450 1609.070 ;
        RECT 2787.910 1609.070 2836.050 1609.370 ;
        RECT 2739.150 1608.390 2787.290 1608.690 ;
        RECT 2690.390 1607.710 2691.610 1608.010 ;
        RECT 2786.990 1608.010 2787.290 1608.390 ;
        RECT 2787.910 1608.010 2788.210 1609.070 ;
        RECT 2835.750 1608.690 2836.050 1609.070 ;
        RECT 2916.710 1608.690 2917.010 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 2835.750 1608.390 2883.890 1608.690 ;
        RECT 2786.990 1607.710 2788.210 1608.010 ;
        RECT 2883.590 1608.010 2883.890 1608.390 ;
        RECT 2884.510 1608.390 2917.010 1608.690 ;
        RECT 2884.510 1608.010 2884.810 1608.390 ;
        RECT 2883.590 1607.710 2884.810 1608.010 ;
        RECT 1896.430 1607.030 1898.570 1607.330 ;
        RECT 1606.385 1606.350 1641.890 1606.650 ;
        RECT 1835.465 1606.650 1835.795 1606.665 ;
        RECT 1882.590 1606.650 1882.970 1606.660 ;
        RECT 1835.465 1606.350 1882.970 1606.650 ;
        RECT 1339.790 1605.970 1340.170 1605.980 ;
        RECT 1386.750 1605.970 1387.050 1606.350 ;
        RECT 1606.385 1606.335 1606.715 1606.350 ;
        RECT 1835.465 1606.335 1835.795 1606.350 ;
        RECT 1882.590 1606.340 1882.970 1606.350 ;
        RECT 1339.790 1605.670 1387.050 1605.970 ;
        RECT 1339.790 1605.660 1340.170 1605.670 ;
      LAYER via3 ;
        RECT 1275.420 2496.460 1275.740 2496.780 ;
        RECT 1275.420 1610.420 1275.740 1610.740 ;
        RECT 1338.900 1608.380 1339.220 1608.700 ;
        RECT 1882.620 1608.380 1882.940 1608.700 ;
        RECT 1339.820 1605.660 1340.140 1605.980 ;
        RECT 1882.620 1606.340 1882.940 1606.660 ;
      LAYER met4 ;
<<<<<<< HEAD
        RECT 1280.935 2497.815 1281.265 2498.145 ;
        RECT 1280.950 1609.385 1281.250 2497.815 ;
        RECT 1280.935 1609.055 1281.265 1609.385 ;
        RECT 1400.535 1609.055 1400.865 1609.385 ;
        RECT 1441.935 1609.055 1442.265 1609.385 ;
        RECT 1400.550 1608.025 1400.850 1609.055 ;
        RECT 1441.950 1608.025 1442.250 1609.055 ;
        RECT 1400.535 1607.695 1400.865 1608.025 ;
        RECT 1441.935 1607.695 1442.265 1608.025 ;
        RECT 1730.815 1607.695 1731.145 1608.025 ;
        RECT 1730.830 1605.305 1731.130 1607.695 ;
        RECT 1730.815 1604.975 1731.145 1605.305 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1275.415 2496.455 1275.745 2496.785 ;
        RECT 1275.430 1610.745 1275.730 2496.455 ;
        RECT 1275.415 1610.415 1275.745 1610.745 ;
        RECT 1338.895 1608.690 1339.225 1608.705 ;
        RECT 1338.895 1608.390 1340.130 1608.690 ;
        RECT 1338.895 1608.375 1339.225 1608.390 ;
        RECT 1339.830 1605.985 1340.130 1608.390 ;
        RECT 1882.615 1608.375 1882.945 1608.705 ;
        RECT 1882.630 1606.665 1882.930 1608.375 ;
        RECT 1882.615 1606.335 1882.945 1606.665 ;
        RECT 1339.815 1605.655 1340.145 1605.985 ;
>>>>>>> re-updated local openlane
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1296.885 2493.985 1297.055 2496.535 ;
      LAYER mcon ;
        RECT 1296.885 2496.365 1297.055 2496.535 ;
      LAYER met1 ;
        RECT 1296.810 2496.520 1297.130 2496.580 ;
        RECT 1296.615 2496.380 1297.130 2496.520 ;
        RECT 1296.810 2496.320 1297.130 2496.380 ;
        RECT 1296.825 2494.140 1297.115 2494.185 ;
        RECT 2059.490 2494.140 2059.810 2494.200 ;
        RECT 1296.825 2494.000 2059.810 2494.140 ;
        RECT 1296.825 2493.955 1297.115 2494.000 ;
        RECT 2059.490 2493.940 2059.810 2494.000 ;
        RECT 2059.490 1849.160 2059.810 1849.220 ;
        RECT 2900.830 1849.160 2901.150 1849.220 ;
        RECT 2059.490 1849.020 2901.150 1849.160 ;
        RECT 2059.490 1848.960 2059.810 1849.020 ;
        RECT 2900.830 1848.960 2901.150 1849.020 ;
      LAYER via ;
        RECT 1296.840 2496.320 1297.100 2496.580 ;
        RECT 2059.520 2493.940 2059.780 2494.200 ;
        RECT 2059.520 1848.960 2059.780 1849.220 ;
        RECT 2900.860 1848.960 2901.120 1849.220 ;
      LAYER met2 ;
        RECT 1294.990 2496.690 1295.270 2500.000 ;
        RECT 1294.990 2496.610 1297.040 2496.690 ;
        RECT 1294.990 2496.550 1297.100 2496.610 ;
        RECT 1294.990 2496.000 1295.270 2496.550 ;
        RECT 1296.840 2496.290 1297.100 2496.550 ;
        RECT 2059.520 2493.910 2059.780 2494.230 ;
        RECT 2059.580 1849.250 2059.720 2493.910 ;
        RECT 2059.520 1848.930 2059.780 1849.250 ;
        RECT 2900.860 1848.930 2901.120 1849.250 ;
        RECT 2900.920 1848.085 2901.060 1848.930 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1847.300 2924.800 1848.500 ;
=======
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1316.130 2499.920 1316.450 2499.980 ;
        RECT 2066.390 2499.920 2066.710 2499.980 ;
        RECT 1316.130 2499.780 2066.710 2499.920 ;
        RECT 1316.130 2499.720 1316.450 2499.780 ;
        RECT 2066.390 2499.720 2066.710 2499.780 ;
        RECT 2066.390 2083.760 2066.710 2083.820 ;
        RECT 2900.830 2083.760 2901.150 2083.820 ;
        RECT 2066.390 2083.620 2901.150 2083.760 ;
        RECT 2066.390 2083.560 2066.710 2083.620 ;
        RECT 2900.830 2083.560 2901.150 2083.620 ;
      LAYER via ;
        RECT 1316.160 2499.720 1316.420 2499.980 ;
        RECT 2066.420 2499.720 2066.680 2499.980 ;
        RECT 2066.420 2083.560 2066.680 2083.820 ;
        RECT 2900.860 2083.560 2901.120 2083.820 ;
      LAYER met2 ;
        RECT 1314.310 2499.410 1314.590 2500.000 ;
        RECT 1316.160 2499.690 1316.420 2500.010 ;
        RECT 2066.420 2499.690 2066.680 2500.010 ;
        RECT 1316.220 2499.410 1316.360 2499.690 ;
        RECT 1314.310 2499.270 1316.360 2499.410 ;
        RECT 1314.310 2496.000 1314.590 2499.270 ;
        RECT 2066.480 2083.850 2066.620 2499.690 ;
        RECT 2066.420 2083.530 2066.680 2083.850 ;
        RECT 2900.860 2083.530 2901.120 2083.850 ;
        RECT 2900.920 2082.685 2901.060 2083.530 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2081.900 2924.800 2083.100 ;
=======
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1333.610 2514.540 1333.930 2514.600 ;
        RECT 1943.570 2514.540 1943.890 2514.600 ;
        RECT 1333.610 2514.400 1943.890 2514.540 ;
        RECT 1333.610 2514.340 1333.930 2514.400 ;
        RECT 1943.570 2514.340 1943.890 2514.400 ;
        RECT 1945.410 2318.360 1945.730 2318.420 ;
        RECT 2900.830 2318.360 2901.150 2318.420 ;
        RECT 1945.410 2318.220 2901.150 2318.360 ;
        RECT 1945.410 2318.160 1945.730 2318.220 ;
        RECT 2900.830 2318.160 2901.150 2318.220 ;
      LAYER via ;
        RECT 1333.640 2514.340 1333.900 2514.600 ;
        RECT 1943.600 2514.340 1943.860 2514.600 ;
        RECT 1945.440 2318.160 1945.700 2318.420 ;
        RECT 2900.860 2318.160 2901.120 2318.420 ;
      LAYER met2 ;
        RECT 1333.640 2514.310 1333.900 2514.630 ;
        RECT 1943.600 2514.310 1943.860 2514.630 ;
        RECT 1333.700 2500.000 1333.840 2514.310 ;
        RECT 1333.630 2496.000 1333.910 2500.000 ;
        RECT 1943.660 2317.850 1943.800 2514.310 ;
        RECT 1945.440 2318.130 1945.700 2318.450 ;
        RECT 2900.860 2318.130 2901.120 2318.450 ;
        RECT 1945.500 2317.850 1945.640 2318.130 ;
        RECT 1943.660 2317.710 1945.640 2317.850 ;
        RECT 2900.920 2317.285 2901.060 2318.130 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2316.500 2924.800 2317.700 ;
=======
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1166.170 2506.040 1166.490 2506.100 ;
        RECT 2011.190 2506.040 2011.510 2506.100 ;
        RECT 1166.170 2505.900 2011.510 2506.040 ;
        RECT 1166.170 2505.840 1166.490 2505.900 ;
        RECT 2011.190 2505.840 2011.510 2505.900 ;
        RECT 2011.190 151.540 2011.510 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 2011.190 151.400 2901.150 151.540 ;
        RECT 2011.190 151.340 2011.510 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 1166.200 2505.840 1166.460 2506.100 ;
        RECT 2011.220 2505.840 2011.480 2506.100 ;
        RECT 2011.220 151.340 2011.480 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 1166.200 2505.810 1166.460 2506.130 ;
        RECT 2011.220 2505.810 2011.480 2506.130 ;
        RECT 1166.260 2500.000 1166.400 2505.810 ;
        RECT 1166.190 2496.000 1166.470 2500.000 ;
        RECT 2011.280 151.630 2011.420 2505.810 ;
        RECT 2011.220 151.310 2011.480 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 145.940 2924.800 147.140 ;
=======
        RECT 1168.005 2498.130 1168.335 2498.145 ;
        RECT 1169.590 2498.130 1169.970 2498.140 ;
        RECT 1168.005 2497.830 1169.970 2498.130 ;
        RECT 1168.005 2497.815 1168.335 2497.830 ;
        RECT 1169.590 2497.820 1169.970 2497.830 ;
        RECT 1290.110 149.410 1290.490 149.420 ;
        RECT 1318.885 149.410 1319.215 149.425 ;
        RECT 1290.110 149.110 1319.215 149.410 ;
        RECT 1290.110 149.100 1290.490 149.110 ;
        RECT 1318.885 149.095 1319.215 149.110 ;
        RECT 1447.470 148.430 1483.650 148.730 ;
        RECT 1169.590 148.050 1169.970 148.060 ;
        RECT 1265.985 148.050 1266.315 148.065 ;
        RECT 1290.110 148.050 1290.490 148.060 ;
        RECT 1169.590 147.750 1200.290 148.050 ;
        RECT 1169.590 147.740 1169.970 147.750 ;
        RECT 1199.990 146.690 1200.290 147.750 ;
        RECT 1265.985 147.750 1290.490 148.050 ;
        RECT 1265.985 147.735 1266.315 147.750 ;
        RECT 1290.110 147.740 1290.490 147.750 ;
        RECT 1200.665 146.690 1200.995 146.705 ;
        RECT 1199.990 146.390 1200.995 146.690 ;
        RECT 1200.665 146.375 1200.995 146.390 ;
        RECT 1318.885 146.690 1319.215 146.705 ;
        RECT 1344.645 146.690 1344.975 146.705 ;
        RECT 1447.470 146.690 1447.770 148.430 ;
        RECT 1483.350 148.050 1483.650 148.430 ;
        RECT 1483.350 147.750 1531.490 148.050 ;
        RECT 1531.190 147.370 1531.490 147.750 ;
        RECT 1702.310 147.750 1738.490 148.050 ;
        RECT 1531.190 147.070 1545.290 147.370 ;
        RECT 1318.885 146.390 1344.975 146.690 ;
        RECT 1318.885 146.375 1319.215 146.390 ;
        RECT 1344.645 146.375 1344.975 146.390 ;
        RECT 1394.110 146.390 1447.770 146.690 ;
        RECT 1394.110 146.010 1394.410 146.390 ;
        RECT 1393.190 145.710 1394.410 146.010 ;
        RECT 1544.990 146.010 1545.290 147.070 ;
        RECT 1617.670 146.390 1641.890 146.690 ;
        RECT 1617.670 146.010 1617.970 146.390 ;
        RECT 1544.990 145.710 1617.970 146.010 ;
        RECT 1386.505 145.330 1386.835 145.345 ;
        RECT 1393.190 145.330 1393.490 145.710 ;
        RECT 1386.505 145.030 1393.490 145.330 ;
        RECT 1641.590 145.330 1641.890 146.390 ;
        RECT 1702.310 146.010 1702.610 147.750 ;
        RECT 1738.190 147.380 1738.490 147.750 ;
        RECT 1798.910 147.750 1835.090 148.050 ;
        RECT 1738.150 147.060 1738.530 147.380 ;
        RECT 1798.910 146.010 1799.210 147.750 ;
        RECT 1834.790 147.380 1835.090 147.750 ;
        RECT 1834.750 147.060 1835.130 147.380 ;
        RECT 1956.445 146.690 1956.775 146.705 ;
        RECT 1993.705 146.690 1994.035 146.705 ;
        RECT 1956.445 146.390 1994.035 146.690 ;
        RECT 1956.445 146.375 1956.775 146.390 ;
        RECT 1993.705 146.375 1994.035 146.390 ;
        RECT 2124.805 146.690 2125.135 146.705 ;
=======
        RECT 2900.825 146.690 2901.155 146.705 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
<<<<<<< HEAD
        RECT 2884.510 145.330 2884.810 145.710 ;
        RECT 2883.590 145.030 2884.810 145.330 ;
        RECT 2069.605 145.015 2069.935 145.030 ;
      LAYER via3 ;
        RECT 1169.620 2497.820 1169.940 2498.140 ;
        RECT 1290.140 149.100 1290.460 149.420 ;
        RECT 1169.620 147.740 1169.940 148.060 ;
        RECT 1290.140 147.740 1290.460 148.060 ;
        RECT 1738.180 147.060 1738.500 147.380 ;
        RECT 1834.780 147.060 1835.100 147.380 ;
        RECT 1738.180 145.020 1738.500 145.340 ;
        RECT 1834.780 145.020 1835.100 145.340 ;
      LAYER met4 ;
        RECT 1169.615 2497.815 1169.945 2498.145 ;
        RECT 1169.630 148.065 1169.930 2497.815 ;
        RECT 1290.135 149.095 1290.465 149.425 ;
        RECT 1290.150 148.065 1290.450 149.095 ;
        RECT 1169.615 147.735 1169.945 148.065 ;
        RECT 1290.135 147.735 1290.465 148.065 ;
        RECT 1738.175 147.055 1738.505 147.385 ;
        RECT 1834.775 147.055 1835.105 147.385 ;
        RECT 1738.190 145.345 1738.490 147.055 ;
        RECT 1834.790 145.345 1835.090 147.055 ;
        RECT 1738.175 145.015 1738.505 145.345 ;
        RECT 1834.775 145.015 1835.105 145.345 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1361.285 2492.285 1361.455 2496.535 ;
      LAYER mcon ;
        RECT 1361.285 2496.365 1361.455 2496.535 ;
      LAYER met1 ;
        RECT 1361.210 2496.520 1361.530 2496.580 ;
        RECT 1361.015 2496.380 1361.530 2496.520 ;
        RECT 1361.210 2496.320 1361.530 2496.380 ;
        RECT 1361.225 2492.440 1361.515 2492.485 ;
        RECT 2899.910 2492.440 2900.230 2492.500 ;
        RECT 1361.225 2492.300 2900.230 2492.440 ;
        RECT 1361.225 2492.255 1361.515 2492.300 ;
        RECT 2899.910 2492.240 2900.230 2492.300 ;
      LAYER via ;
        RECT 1361.240 2496.320 1361.500 2496.580 ;
        RECT 2899.940 2492.240 2900.200 2492.500 ;
      LAYER met2 ;
        RECT 1359.390 2496.690 1359.670 2500.000 ;
        RECT 1359.390 2496.610 1361.440 2496.690 ;
        RECT 1359.390 2496.550 1361.500 2496.610 ;
        RECT 1359.390 2496.000 1359.670 2496.550 ;
        RECT 1361.240 2496.290 1361.500 2496.550 ;
        RECT 2899.930 2493.035 2900.210 2493.405 ;
        RECT 2900.000 2492.530 2900.140 2493.035 ;
        RECT 2899.940 2492.210 2900.200 2492.530 ;
      LAYER via2 ;
        RECT 2899.930 2493.080 2900.210 2493.360 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 2492.620 2924.800 2493.820 ;
=======
        RECT 2900.825 2493.370 2901.155 2493.385 ;
=======
        RECT 2899.905 2493.370 2900.235 2493.385 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2899.905 2493.070 2924.800 2493.370 ;
        RECT 2899.905 2493.055 2900.235 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1379.610 2725.680 1379.930 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 1379.610 2725.540 2901.150 2725.680 ;
        RECT 1379.610 2725.480 1379.930 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
      LAYER via ;
        RECT 1379.640 2725.480 1379.900 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 1379.640 2725.450 1379.900 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 1378.710 2499.410 1378.990 2500.000 ;
        RECT 1379.700 2499.410 1379.840 2725.450 ;
        RECT 1378.710 2499.270 1379.840 2499.410 ;
        RECT 1378.710 2496.000 1378.990 2499.270 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2727.220 2924.800 2728.420 ;
=======
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1400.310 2960.280 1400.630 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 1400.310 2960.140 2901.150 2960.280 ;
        RECT 1400.310 2960.080 1400.630 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 1400.340 2960.080 1400.600 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 1400.340 2960.050 1400.600 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 1398.030 2499.410 1398.310 2500.000 ;
        RECT 1400.400 2499.410 1400.540 2960.050 ;
        RECT 1398.030 2499.270 1400.540 2499.410 ;
        RECT 1398.030 2496.000 1398.310 2499.270 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2961.820 2924.800 2963.020 ;
=======
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 3194.880 1421.330 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 1421.010 3194.740 2901.150 3194.880 ;
        RECT 1421.010 3194.680 1421.330 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 1421.040 3194.680 1421.300 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 1421.040 3194.650 1421.300 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 1417.350 2499.410 1417.630 2500.000 ;
        RECT 1421.100 2499.410 1421.240 3194.650 ;
        RECT 1417.350 2499.270 1421.240 2499.410 ;
        RECT 1417.350 2496.000 1417.630 2499.270 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3196.420 2924.800 3197.620 ;
=======
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2146.060 3429.680 2149.880 3429.820 ;
        RECT 1441.710 3429.480 1442.030 3429.540 ;
        RECT 2146.060 3429.480 2146.200 3429.680 ;
        RECT 1441.710 3429.340 2146.200 3429.480 ;
        RECT 2149.740 3429.480 2149.880 3429.680 ;
        RECT 2228.860 3429.680 2231.300 3429.820 ;
        RECT 2228.860 3429.480 2229.000 3429.680 ;
        RECT 2149.740 3429.340 2229.000 3429.480 ;
        RECT 2231.160 3429.480 2231.300 3429.680 ;
        RECT 2762.920 3429.680 2798.940 3429.820 ;
        RECT 2762.920 3429.480 2763.060 3429.680 ;
        RECT 2231.160 3429.340 2763.060 3429.480 ;
        RECT 2798.800 3429.480 2798.940 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2798.800 3429.340 2901.150 3429.480 ;
        RECT 1441.710 3429.280 1442.030 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
        RECT 1437.110 2515.900 1437.430 2515.960 ;
        RECT 1441.710 2515.900 1442.030 2515.960 ;
        RECT 1437.110 2515.760 1442.030 2515.900 ;
        RECT 1437.110 2515.700 1437.430 2515.760 ;
        RECT 1441.710 2515.700 1442.030 2515.760 ;
      LAYER via ;
        RECT 1441.740 3429.280 1442.000 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
        RECT 1437.140 2515.700 1437.400 2515.960 ;
        RECT 1441.740 2515.700 1442.000 2515.960 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1441.740 3429.250 1442.000 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1441.800 2515.990 1441.940 3429.250 ;
        RECT 1437.140 2515.670 1437.400 2515.990 ;
        RECT 1441.740 2515.670 1442.000 2515.990 ;
        RECT 1437.200 2500.000 1437.340 2515.670 ;
        RECT 1437.130 2496.000 1437.410 2500.000 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 3431.020 2924.800 3432.220 ;
=======
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1462.410 3502.240 1462.730 3502.300 ;
        RECT 2717.290 3502.240 2717.610 3502.300 ;
        RECT 1462.410 3502.100 2717.610 3502.240 ;
        RECT 1462.410 3502.040 1462.730 3502.100 ;
        RECT 2717.290 3502.040 2717.610 3502.100 ;
        RECT 1456.430 2516.240 1456.750 2516.300 ;
        RECT 1462.410 2516.240 1462.730 2516.300 ;
        RECT 1456.430 2516.100 1462.730 2516.240 ;
        RECT 1456.430 2516.040 1456.750 2516.100 ;
        RECT 1462.410 2516.040 1462.730 2516.100 ;
      LAYER via ;
        RECT 1462.440 3502.040 1462.700 3502.300 ;
        RECT 2717.320 3502.040 2717.580 3502.300 ;
        RECT 1456.460 2516.040 1456.720 2516.300 ;
        RECT 1462.440 2516.040 1462.700 2516.300 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2717.170 3519.700 2717.730 3524.800 ;
=======
        RECT 2717.170 3517.600 2717.730 3524.800 ;
<<<<<<< HEAD
        RECT 2717.380 3517.370 2717.520 3517.600 ;
        RECT 2717.380 3517.230 2717.980 3517.370 ;
        RECT 2717.840 3491.450 2717.980 3517.230 ;
        RECT 2713.640 3491.130 2713.900 3491.450 ;
        RECT 2717.780 3491.130 2718.040 3491.450 ;
        RECT 2713.700 3443.510 2713.840 3491.130 ;
        RECT 2713.640 3443.190 2713.900 3443.510 ;
        RECT 2712.720 3442.850 2712.980 3443.170 ;
        RECT 2712.780 3429.650 2712.920 3442.850 ;
        RECT 2712.320 3429.510 2712.920 3429.650 ;
        RECT 2712.320 3422.430 2712.460 3429.510 ;
        RECT 2712.260 3422.110 2712.520 3422.430 ;
        RECT 2714.100 3332.690 2714.360 3333.010 ;
        RECT 2714.160 3298.410 2714.300 3332.690 ;
        RECT 2713.240 3298.270 2714.300 3298.410 ;
        RECT 2713.240 3236.450 2713.380 3298.270 ;
        RECT 2712.720 3236.130 2712.980 3236.450 ;
        RECT 2713.180 3236.130 2713.440 3236.450 ;
        RECT 2712.780 3201.850 2712.920 3236.130 ;
        RECT 2712.780 3201.710 2713.380 3201.850 ;
        RECT 2713.240 3187.830 2713.380 3201.710 ;
        RECT 2713.180 3187.510 2713.440 3187.830 ;
        RECT 2713.640 3139.570 2713.900 3139.890 ;
        RECT 2713.700 3132.750 2713.840 3139.570 ;
        RECT 2713.640 3132.430 2713.900 3132.750 ;
        RECT 2712.720 3088.570 2712.980 3088.890 ;
        RECT 2712.780 3084.325 2712.920 3088.570 ;
        RECT 2712.710 3083.955 2712.990 3084.325 ;
        RECT 2713.630 3083.955 2713.910 3084.325 ;
        RECT 2713.700 3036.530 2713.840 3083.955 ;
        RECT 2713.180 3036.210 2713.440 3036.530 ;
        RECT 2713.640 3036.210 2713.900 3036.530 ;
        RECT 2713.240 3035.930 2713.380 3036.210 ;
        RECT 2713.240 3035.850 2713.840 3035.930 ;
        RECT 2713.240 3035.790 2713.900 3035.850 ;
        RECT 2713.640 3035.530 2713.900 3035.790 ;
        RECT 2714.100 2946.450 2714.360 2946.770 ;
        RECT 2714.160 2912.430 2714.300 2946.450 ;
        RECT 2714.100 2912.110 2714.360 2912.430 ;
        RECT 2713.640 2911.430 2713.900 2911.750 ;
        RECT 2713.700 2863.210 2713.840 2911.430 ;
        RECT 2712.780 2863.070 2713.840 2863.210 ;
        RECT 2712.780 2849.610 2712.920 2863.070 ;
        RECT 2712.320 2849.470 2712.920 2849.610 ;
        RECT 2712.320 2815.870 2712.460 2849.470 ;
        RECT 2712.260 2815.550 2712.520 2815.870 ;
        RECT 2712.260 2814.870 2712.520 2815.190 ;
        RECT 2712.320 2801.250 2712.460 2814.870 ;
        RECT 2712.260 2800.930 2712.520 2801.250 ;
        RECT 2713.180 2752.990 2713.440 2753.310 ;
        RECT 2713.240 2718.290 2713.380 2752.990 ;
        RECT 2712.260 2717.970 2712.520 2718.290 ;
        RECT 2713.180 2717.970 2713.440 2718.290 ;
        RECT 2712.320 2670.350 2712.460 2717.970 ;
        RECT 2712.260 2670.030 2712.520 2670.350 ;
        RECT 2713.180 2670.030 2713.440 2670.350 ;
        RECT 2713.240 2622.410 2713.380 2670.030 ;
        RECT 2713.180 2622.090 2713.440 2622.410 ;
        RECT 2713.640 2621.750 2713.900 2622.070 ;
        RECT 2713.700 2608.325 2713.840 2621.750 ;
        RECT 2712.710 2607.955 2712.990 2608.325 ;
        RECT 2713.630 2607.955 2713.910 2608.325 ;
        RECT 2712.780 2560.190 2712.920 2607.955 ;
        RECT 2712.720 2559.870 2712.980 2560.190 ;
        RECT 2714.100 2559.870 2714.360 2560.190 ;
        RECT 1463.820 2514.990 1464.080 2515.310 ;
        RECT 1463.880 2500.000 1464.020 2514.990 ;
        RECT 2714.160 2514.970 2714.300 2559.870 ;
        RECT 2714.100 2514.650 2714.360 2514.970 ;
        RECT 1463.810 2496.000 1464.090 2500.000 ;
      LAYER via2 ;
        RECT 2712.710 3084.000 2712.990 3084.280 ;
        RECT 2713.630 3084.000 2713.910 3084.280 ;
        RECT 2712.710 2608.000 2712.990 2608.280 ;
        RECT 2713.630 2608.000 2713.910 2608.280 ;
      LAYER met3 ;
        RECT 2712.685 3084.290 2713.015 3084.305 ;
        RECT 2713.605 3084.290 2713.935 3084.305 ;
        RECT 2712.685 3083.990 2713.935 3084.290 ;
        RECT 2712.685 3083.975 2713.015 3083.990 ;
        RECT 2713.605 3083.975 2713.935 3083.990 ;
        RECT 2712.685 2608.290 2713.015 2608.305 ;
        RECT 2713.605 2608.290 2713.935 2608.305 ;
        RECT 2712.685 2607.990 2713.935 2608.290 ;
        RECT 2712.685 2607.975 2713.015 2607.990 ;
        RECT 2713.605 2607.975 2713.935 2607.990 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2717.380 3502.330 2717.520 3517.600 ;
        RECT 1462.440 3502.010 1462.700 3502.330 ;
        RECT 2717.320 3502.010 2717.580 3502.330 ;
        RECT 1462.500 2516.330 1462.640 3502.010 ;
        RECT 1456.460 2516.010 1456.720 2516.330 ;
        RECT 1462.440 2516.010 1462.700 2516.330 ;
        RECT 1456.520 2500.000 1456.660 2516.010 ;
        RECT 1456.450 2496.000 1456.730 2500.000 ;
>>>>>>> re-updated local openlane
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1476.210 3503.940 1476.530 3504.000 ;
        RECT 2392.530 3503.940 2392.850 3504.000 ;
        RECT 1476.210 3503.800 2392.850 3503.940 ;
        RECT 1476.210 3503.740 1476.530 3503.800 ;
        RECT 2392.530 3503.740 2392.850 3503.800 ;
      LAYER via ;
        RECT 1476.240 3503.740 1476.500 3504.000 ;
        RECT 2392.560 3503.740 2392.820 3504.000 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2392.410 3519.700 2392.970 3524.800 ;
=======
        RECT 2392.410 3517.600 2392.970 3524.800 ;
<<<<<<< HEAD
        RECT 2392.620 3517.370 2392.760 3517.600 ;
        RECT 2392.620 3517.230 2393.220 3517.370 ;
        RECT 2393.080 3430.445 2393.220 3517.230 ;
        RECT 2393.010 3430.075 2393.290 3430.445 ;
        RECT 2388.410 3429.395 2388.690 3429.765 ;
        RECT 2388.480 3394.970 2388.620 3429.395 ;
        RECT 2387.560 3394.830 2388.620 3394.970 ;
        RECT 2387.560 3380.950 2387.700 3394.830 ;
        RECT 2387.500 3380.630 2387.760 3380.950 ;
        RECT 2387.960 3332.690 2388.220 3333.010 ;
        RECT 2388.020 3298.410 2388.160 3332.690 ;
        RECT 2388.020 3298.270 2388.620 3298.410 ;
        RECT 2388.480 3270.790 2388.620 3298.270 ;
        RECT 2387.500 3270.470 2387.760 3270.790 ;
        RECT 2388.420 3270.470 2388.680 3270.790 ;
        RECT 2387.560 3222.250 2387.700 3270.470 ;
        RECT 2387.560 3222.110 2388.620 3222.250 ;
        RECT 2388.480 3174.230 2388.620 3222.110 ;
        RECT 2387.500 3173.910 2387.760 3174.230 ;
        RECT 2388.420 3173.910 2388.680 3174.230 ;
        RECT 2387.560 3125.690 2387.700 3173.910 ;
        RECT 2387.560 3125.550 2388.620 3125.690 ;
        RECT 2388.480 3077.670 2388.620 3125.550 ;
        RECT 2387.500 3077.350 2387.760 3077.670 ;
        RECT 2388.420 3077.350 2388.680 3077.670 ;
        RECT 2387.560 3029.130 2387.700 3077.350 ;
        RECT 2387.560 3028.990 2388.620 3029.130 ;
        RECT 2388.480 2981.110 2388.620 3028.990 ;
        RECT 2387.500 2980.850 2387.760 2981.110 ;
        RECT 2387.500 2980.790 2388.160 2980.850 ;
        RECT 2388.420 2980.790 2388.680 2981.110 ;
        RECT 2387.560 2980.710 2388.160 2980.790 ;
        RECT 2388.020 2980.170 2388.160 2980.710 ;
        RECT 2388.020 2980.030 2388.620 2980.170 ;
        RECT 2388.480 2959.770 2388.620 2980.030 ;
        RECT 2388.020 2959.630 2388.620 2959.770 ;
        RECT 2388.020 2946.430 2388.160 2959.630 ;
        RECT 2386.580 2946.110 2386.840 2946.430 ;
        RECT 2387.960 2946.110 2388.220 2946.430 ;
        RECT 2386.640 2898.685 2386.780 2946.110 ;
        RECT 2386.570 2898.315 2386.850 2898.685 ;
        RECT 2387.490 2898.315 2387.770 2898.685 ;
        RECT 2387.560 2863.210 2387.700 2898.315 ;
        RECT 2387.560 2863.070 2388.160 2863.210 ;
        RECT 2388.020 2849.530 2388.160 2863.070 ;
        RECT 2387.960 2849.210 2388.220 2849.530 ;
        RECT 2388.880 2815.210 2389.140 2815.530 ;
        RECT 2388.940 2801.445 2389.080 2815.210 ;
        RECT 2387.950 2801.075 2388.230 2801.445 ;
        RECT 2388.870 2801.075 2389.150 2801.445 ;
        RECT 2388.020 2753.310 2388.160 2801.075 ;
        RECT 2387.960 2752.990 2388.220 2753.310 ;
        RECT 2389.340 2752.990 2389.600 2753.310 ;
        RECT 2389.400 2719.310 2389.540 2752.990 ;
        RECT 2389.340 2718.990 2389.600 2719.310 ;
        RECT 2388.880 2718.310 2389.140 2718.630 ;
        RECT 2388.940 2670.690 2389.080 2718.310 ;
        RECT 2388.880 2670.370 2389.140 2670.690 ;
        RECT 2389.340 2669.690 2389.600 2670.010 ;
        RECT 2389.400 2649.610 2389.540 2669.690 ;
        RECT 2389.340 2649.290 2389.600 2649.610 ;
        RECT 2390.260 2649.290 2390.520 2649.610 ;
        RECT 2390.320 2573.450 2390.460 2649.290 ;
        RECT 2389.340 2573.130 2389.600 2573.450 ;
        RECT 2390.260 2573.130 2390.520 2573.450 ;
        RECT 2389.400 2515.310 2389.540 2573.130 ;
        RECT 1485.440 2514.990 1485.700 2515.310 ;
        RECT 2389.340 2514.990 2389.600 2515.310 ;
        RECT 1483.590 2499.410 1483.870 2500.000 ;
        RECT 1485.500 2499.410 1485.640 2514.990 ;
        RECT 1483.590 2499.270 1485.640 2499.410 ;
        RECT 1483.590 2496.000 1483.870 2499.270 ;
      LAYER via2 ;
        RECT 2393.010 3430.120 2393.290 3430.400 ;
        RECT 2388.410 3429.440 2388.690 3429.720 ;
        RECT 2386.570 2898.360 2386.850 2898.640 ;
        RECT 2387.490 2898.360 2387.770 2898.640 ;
        RECT 2387.950 2801.120 2388.230 2801.400 ;
        RECT 2388.870 2801.120 2389.150 2801.400 ;
      LAYER met3 ;
        RECT 2392.985 3430.410 2393.315 3430.425 ;
        RECT 2387.710 3430.110 2393.315 3430.410 ;
        RECT 2387.710 3429.730 2388.010 3430.110 ;
        RECT 2392.985 3430.095 2393.315 3430.110 ;
        RECT 2388.385 3429.730 2388.715 3429.745 ;
        RECT 2387.710 3429.430 2388.715 3429.730 ;
        RECT 2388.385 3429.415 2388.715 3429.430 ;
        RECT 2386.545 2898.650 2386.875 2898.665 ;
        RECT 2387.465 2898.650 2387.795 2898.665 ;
        RECT 2386.545 2898.350 2387.795 2898.650 ;
        RECT 2386.545 2898.335 2386.875 2898.350 ;
        RECT 2387.465 2898.335 2387.795 2898.350 ;
        RECT 2387.925 2801.410 2388.255 2801.425 ;
        RECT 2388.845 2801.410 2389.175 2801.425 ;
        RECT 2387.925 2801.110 2389.175 2801.410 ;
        RECT 2387.925 2801.095 2388.255 2801.110 ;
        RECT 2388.845 2801.095 2389.175 2801.110 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2392.620 3504.030 2392.760 3517.600 ;
        RECT 1476.240 3503.710 1476.500 3504.030 ;
        RECT 2392.560 3503.710 2392.820 3504.030 ;
        RECT 1475.770 2499.410 1476.050 2500.000 ;
        RECT 1476.300 2499.410 1476.440 3503.710 ;
        RECT 1475.770 2499.270 1476.440 2499.410 ;
        RECT 1475.770 2496.000 1476.050 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1496.910 3500.880 1497.230 3500.940 ;
        RECT 2068.230 3500.880 2068.550 3500.940 ;
        RECT 1496.910 3500.740 2068.550 3500.880 ;
        RECT 1496.910 3500.680 1497.230 3500.740 ;
        RECT 2068.230 3500.680 2068.550 3500.740 ;
      LAYER via ;
        RECT 1496.940 3500.680 1497.200 3500.940 ;
        RECT 2068.260 3500.680 2068.520 3500.940 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2068.110 3519.700 2068.670 3524.800 ;
=======
        RECT 2068.110 3517.600 2068.670 3524.800 ;
<<<<<<< HEAD
        RECT 2068.320 3517.370 2068.460 3517.600 ;
        RECT 2068.320 3517.230 2068.920 3517.370 ;
        RECT 2068.780 3491.450 2068.920 3517.230 ;
        RECT 2065.040 3491.130 2065.300 3491.450 ;
        RECT 2068.720 3491.130 2068.980 3491.450 ;
        RECT 2065.100 3443.510 2065.240 3491.130 ;
        RECT 2065.040 3443.190 2065.300 3443.510 ;
        RECT 2064.120 3442.850 2064.380 3443.170 ;
        RECT 2064.180 3429.650 2064.320 3442.850 ;
        RECT 2063.720 3429.510 2064.320 3429.650 ;
        RECT 2063.720 3422.430 2063.860 3429.510 ;
        RECT 2063.660 3422.110 2063.920 3422.430 ;
        RECT 2065.500 3332.690 2065.760 3333.010 ;
        RECT 2065.560 3298.410 2065.700 3332.690 ;
        RECT 2064.640 3298.270 2065.700 3298.410 ;
        RECT 2064.640 3236.450 2064.780 3298.270 ;
        RECT 2064.120 3236.130 2064.380 3236.450 ;
        RECT 2064.580 3236.130 2064.840 3236.450 ;
        RECT 2064.180 3202.110 2064.320 3236.130 ;
        RECT 2064.120 3201.790 2064.380 3202.110 ;
        RECT 2064.580 3201.790 2064.840 3202.110 ;
        RECT 2064.640 3153.490 2064.780 3201.790 ;
        RECT 2063.660 3153.170 2063.920 3153.490 ;
        RECT 2064.580 3153.170 2064.840 3153.490 ;
        RECT 2063.720 3152.890 2063.860 3153.170 ;
        RECT 2063.720 3152.750 2064.320 3152.890 ;
        RECT 2064.180 3105.290 2064.320 3152.750 ;
        RECT 2064.180 3105.150 2064.780 3105.290 ;
        RECT 2064.640 3056.930 2064.780 3105.150 ;
        RECT 2063.660 3056.610 2063.920 3056.930 ;
        RECT 2064.580 3056.610 2064.840 3056.930 ;
        RECT 2063.720 3056.330 2063.860 3056.610 ;
        RECT 2063.720 3056.190 2064.320 3056.330 ;
        RECT 2064.180 3042.990 2064.320 3056.190 ;
        RECT 2064.120 3042.670 2064.380 3042.990 ;
        RECT 2065.040 3008.330 2065.300 3008.650 ;
        RECT 2065.100 2994.710 2065.240 3008.330 ;
        RECT 2065.040 2994.390 2065.300 2994.710 ;
        RECT 2065.500 2946.450 2065.760 2946.770 ;
        RECT 2065.560 2912.430 2065.700 2946.450 ;
        RECT 2065.500 2912.110 2065.760 2912.430 ;
        RECT 2065.040 2911.430 2065.300 2911.750 ;
        RECT 2065.100 2863.210 2065.240 2911.430 ;
        RECT 2064.180 2863.070 2065.240 2863.210 ;
        RECT 2064.180 2849.610 2064.320 2863.070 ;
        RECT 2063.720 2849.470 2064.320 2849.610 ;
        RECT 2063.720 2815.870 2063.860 2849.470 ;
        RECT 2063.660 2815.550 2063.920 2815.870 ;
        RECT 2063.660 2814.870 2063.920 2815.190 ;
        RECT 2063.720 2801.250 2063.860 2814.870 ;
        RECT 2063.660 2800.930 2063.920 2801.250 ;
        RECT 2064.580 2752.990 2064.840 2753.310 ;
        RECT 2064.640 2718.290 2064.780 2752.990 ;
        RECT 2063.660 2717.970 2063.920 2718.290 ;
        RECT 2064.580 2717.970 2064.840 2718.290 ;
        RECT 2063.720 2670.350 2063.860 2717.970 ;
        RECT 2063.660 2670.030 2063.920 2670.350 ;
        RECT 2064.580 2670.030 2064.840 2670.350 ;
        RECT 2064.640 2622.410 2064.780 2670.030 ;
        RECT 2064.580 2622.090 2064.840 2622.410 ;
        RECT 2065.040 2621.750 2065.300 2622.070 ;
        RECT 2065.100 2608.325 2065.240 2621.750 ;
        RECT 2064.110 2607.955 2064.390 2608.325 ;
        RECT 2065.030 2607.955 2065.310 2608.325 ;
        RECT 2064.180 2560.190 2064.320 2607.955 ;
        RECT 2064.120 2559.870 2064.380 2560.190 ;
        RECT 2065.500 2559.870 2065.760 2560.190 ;
        RECT 1503.380 2517.710 1503.640 2518.030 ;
        RECT 1503.440 2500.000 1503.580 2517.710 ;
        RECT 2065.560 2517.690 2065.700 2559.870 ;
        RECT 2065.500 2517.370 2065.760 2517.690 ;
        RECT 1503.370 2496.000 1503.650 2500.000 ;
      LAYER via2 ;
        RECT 2064.110 2608.000 2064.390 2608.280 ;
        RECT 2065.030 2608.000 2065.310 2608.280 ;
      LAYER met3 ;
        RECT 2064.085 2608.290 2064.415 2608.305 ;
        RECT 2065.005 2608.290 2065.335 2608.305 ;
        RECT 2064.085 2607.990 2065.335 2608.290 ;
        RECT 2064.085 2607.975 2064.415 2607.990 ;
        RECT 2065.005 2607.975 2065.335 2607.990 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2068.320 3500.970 2068.460 3517.600 ;
        RECT 1496.940 3500.650 1497.200 3500.970 ;
        RECT 2068.260 3500.650 2068.520 3500.970 ;
        RECT 1495.090 2499.410 1495.370 2500.000 ;
        RECT 1497.000 2499.410 1497.140 3500.650 ;
        RECT 1495.090 2499.270 1497.140 2499.410 ;
        RECT 1495.090 2496.000 1495.370 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1517.610 3499.520 1517.930 3499.580 ;
        RECT 1743.930 3499.520 1744.250 3499.580 ;
        RECT 1517.610 3499.380 1744.250 3499.520 ;
        RECT 1517.610 3499.320 1517.930 3499.380 ;
        RECT 1743.930 3499.320 1744.250 3499.380 ;
      LAYER via ;
        RECT 1517.640 3499.320 1517.900 3499.580 ;
        RECT 1743.960 3499.320 1744.220 3499.580 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1743.810 3519.700 1744.370 3524.800 ;
=======
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3499.610 1744.160 3517.600 ;
        RECT 1517.640 3499.290 1517.900 3499.610 ;
        RECT 1743.960 3499.290 1744.220 3499.610 ;
<<<<<<< HEAD
        RECT 1523.150 2499.410 1523.430 2500.000 ;
        RECT 1524.600 2499.410 1524.740 3499.290 ;
        RECT 1523.150 2499.270 1524.740 2499.410 ;
        RECT 1523.150 2496.000 1523.430 2499.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1517.700 2500.090 1517.840 3499.290 ;
        RECT 1514.410 2499.410 1514.690 2500.000 ;
        RECT 1515.860 2499.950 1517.840 2500.090 ;
        RECT 1515.860 2499.410 1516.000 2499.950 ;
        RECT 1514.410 2499.270 1516.000 2499.410 ;
        RECT 1514.410 2496.000 1514.690 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1468.925 3496.985 1469.095 3499.535 ;
        RECT 1496.985 3496.985 1497.155 3497.835 ;
        RECT 1497.445 3494.265 1497.615 3498.175 ;
      LAYER mcon ;
        RECT 1468.925 3499.365 1469.095 3499.535 ;
        RECT 1497.445 3498.005 1497.615 3498.175 ;
        RECT 1496.985 3497.665 1497.155 3497.835 ;
      LAYER met1 ;
        RECT 1419.170 3499.520 1419.490 3499.580 ;
        RECT 1468.865 3499.520 1469.155 3499.565 ;
        RECT 1419.170 3499.380 1469.155 3499.520 ;
        RECT 1419.170 3499.320 1419.490 3499.380 ;
        RECT 1468.865 3499.335 1469.155 3499.380 ;
        RECT 1497.385 3498.160 1497.675 3498.205 ;
        RECT 1497.000 3498.020 1497.675 3498.160 ;
        RECT 1497.000 3497.865 1497.140 3498.020 ;
        RECT 1497.385 3497.975 1497.675 3498.020 ;
        RECT 1496.925 3497.635 1497.215 3497.865 ;
        RECT 1468.865 3497.140 1469.155 3497.185 ;
        RECT 1496.925 3497.140 1497.215 3497.185 ;
        RECT 1468.865 3497.000 1497.215 3497.140 ;
        RECT 1468.865 3496.955 1469.155 3497.000 ;
        RECT 1496.925 3496.955 1497.215 3497.000 ;
        RECT 1497.385 3494.420 1497.675 3494.465 ;
        RECT 1531.870 3494.420 1532.190 3494.480 ;
        RECT 1497.385 3494.280 1532.190 3494.420 ;
        RECT 1497.385 3494.235 1497.675 3494.280 ;
        RECT 1531.870 3494.220 1532.190 3494.280 ;
      LAYER via ;
        RECT 1419.200 3499.320 1419.460 3499.580 ;
        RECT 1531.900 3494.220 1532.160 3494.480 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1419.050 3519.700 1419.610 3524.800 ;
=======
        RECT 1419.050 3517.600 1419.610 3524.800 ;
<<<<<<< HEAD
        RECT 1419.260 3517.370 1419.400 3517.600 ;
        RECT 1418.800 3517.230 1419.400 3517.370 ;
        RECT 1418.800 3478.190 1418.940 3517.230 ;
        RECT 1418.740 3477.870 1419.000 3478.190 ;
        RECT 1419.660 3477.870 1419.920 3478.190 ;
        RECT 1419.720 3443.170 1419.860 3477.870 ;
        RECT 1419.660 3442.850 1419.920 3443.170 ;
        RECT 1420.580 3442.850 1420.840 3443.170 ;
        RECT 1420.640 3429.230 1420.780 3442.850 ;
        RECT 1420.580 3428.910 1420.840 3429.230 ;
        RECT 1420.120 3380.970 1420.380 3381.290 ;
        RECT 1420.180 3367.690 1420.320 3380.970 ;
        RECT 1420.120 3367.370 1420.380 3367.690 ;
        RECT 1421.040 3367.370 1421.300 3367.690 ;
        RECT 1421.100 3318.810 1421.240 3367.370 ;
        RECT 1420.180 3318.670 1421.240 3318.810 ;
        RECT 1420.180 3270.790 1420.320 3318.670 ;
        RECT 1420.120 3270.470 1420.380 3270.790 ;
        RECT 1421.040 3270.470 1421.300 3270.790 ;
        RECT 1421.100 3222.170 1421.240 3270.470 ;
        RECT 1419.660 3221.850 1419.920 3222.170 ;
        RECT 1421.040 3221.850 1421.300 3222.170 ;
        RECT 1419.720 3174.230 1419.860 3221.850 ;
        RECT 1419.660 3173.910 1419.920 3174.230 ;
        RECT 1421.040 3173.910 1421.300 3174.230 ;
        RECT 1421.100 3125.610 1421.240 3173.910 ;
        RECT 1419.660 3125.290 1419.920 3125.610 ;
        RECT 1421.040 3125.290 1421.300 3125.610 ;
        RECT 1419.720 3077.670 1419.860 3125.290 ;
        RECT 1419.660 3077.350 1419.920 3077.670 ;
        RECT 1421.040 3077.350 1421.300 3077.670 ;
        RECT 1421.100 3029.050 1421.240 3077.350 ;
        RECT 1419.660 3028.730 1419.920 3029.050 ;
        RECT 1421.040 3028.730 1421.300 3029.050 ;
        RECT 1419.720 2981.110 1419.860 3028.730 ;
        RECT 1419.660 2980.790 1419.920 2981.110 ;
        RECT 1421.040 2980.790 1421.300 2981.110 ;
        RECT 1421.100 2932.490 1421.240 2980.790 ;
        RECT 1419.660 2932.170 1419.920 2932.490 ;
        RECT 1421.040 2932.170 1421.300 2932.490 ;
        RECT 1419.720 2884.550 1419.860 2932.170 ;
        RECT 1419.660 2884.230 1419.920 2884.550 ;
        RECT 1421.040 2884.230 1421.300 2884.550 ;
        RECT 1421.100 2835.930 1421.240 2884.230 ;
        RECT 1419.660 2835.610 1419.920 2835.930 ;
        RECT 1421.040 2835.610 1421.300 2835.930 ;
        RECT 1419.720 2787.990 1419.860 2835.610 ;
        RECT 1419.660 2787.670 1419.920 2787.990 ;
        RECT 1421.040 2787.670 1421.300 2787.990 ;
        RECT 1421.100 2739.370 1421.240 2787.670 ;
        RECT 1419.660 2739.050 1419.920 2739.370 ;
        RECT 1421.040 2739.050 1421.300 2739.370 ;
        RECT 1419.720 2691.285 1419.860 2739.050 ;
        RECT 1419.650 2690.915 1419.930 2691.285 ;
        RECT 1421.030 2690.915 1421.310 2691.285 ;
        RECT 1421.100 2642.810 1421.240 2690.915 ;
        RECT 1419.660 2642.490 1419.920 2642.810 ;
        RECT 1421.040 2642.490 1421.300 2642.810 ;
        RECT 1419.720 2594.870 1419.860 2642.490 ;
        RECT 1419.660 2594.550 1419.920 2594.870 ;
        RECT 1421.040 2594.550 1421.300 2594.870 ;
        RECT 1421.100 2546.250 1421.240 2594.550 ;
        RECT 1420.120 2545.930 1420.380 2546.250 ;
        RECT 1421.040 2545.930 1421.300 2546.250 ;
        RECT 1420.180 2518.370 1420.320 2545.930 ;
        RECT 1541.100 2518.390 1541.360 2518.710 ;
        RECT 1420.120 2518.050 1420.380 2518.370 ;
        RECT 1541.160 2499.410 1541.300 2518.390 ;
        RECT 1542.930 2499.410 1543.210 2500.000 ;
        RECT 1541.160 2499.270 1543.210 2499.410 ;
        RECT 1542.930 2496.000 1543.210 2499.270 ;
      LAYER via2 ;
        RECT 1419.650 2690.960 1419.930 2691.240 ;
        RECT 1421.030 2690.960 1421.310 2691.240 ;
      LAYER met3 ;
        RECT 1419.625 2691.250 1419.955 2691.265 ;
        RECT 1421.005 2691.250 1421.335 2691.265 ;
        RECT 1419.625 2690.950 1421.335 2691.250 ;
        RECT 1419.625 2690.935 1419.955 2690.950 ;
        RECT 1421.005 2690.935 1421.335 2690.950 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1419.260 3499.610 1419.400 3517.600 ;
        RECT 1419.200 3499.290 1419.460 3499.610 ;
        RECT 1531.900 3494.190 1532.160 3494.510 ;
        RECT 1531.960 2499.410 1532.100 3494.190 ;
        RECT 1533.730 2499.410 1534.010 2500.000 ;
        RECT 1531.960 2499.270 1534.010 2499.410 ;
        RECT 1533.730 2496.000 1534.010 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1457.350 380.700 1457.670 380.760 ;
        RECT 1496.910 380.700 1497.230 380.760 ;
        RECT 1457.350 380.560 1497.230 380.700 ;
        RECT 1457.350 380.500 1457.670 380.560 ;
        RECT 1496.910 380.500 1497.230 380.560 ;
        RECT 2090.310 380.700 2090.630 380.760 ;
        RECT 2124.810 380.700 2125.130 380.760 ;
        RECT 2090.310 380.560 2125.130 380.700 ;
        RECT 2090.310 380.500 2090.630 380.560 ;
        RECT 2124.810 380.500 2125.130 380.560 ;
        RECT 2476.710 380.700 2477.030 380.760 ;
        RECT 2528.690 380.700 2529.010 380.760 ;
        RECT 2476.710 380.560 2529.010 380.700 ;
        RECT 2476.710 380.500 2477.030 380.560 ;
        RECT 2528.690 380.500 2529.010 380.560 ;
        RECT 1799.130 380.360 1799.450 380.420 ;
        RECT 1801.890 380.360 1802.210 380.420 ;
        RECT 1799.130 380.220 1802.210 380.360 ;
        RECT 1799.130 380.160 1799.450 380.220 ;
        RECT 1801.890 380.160 1802.210 380.220 ;
        RECT 2621.610 380.360 2621.930 380.420 ;
        RECT 2625.750 380.360 2626.070 380.420 ;
        RECT 2621.610 380.220 2626.070 380.360 ;
        RECT 2621.610 380.160 2621.930 380.220 ;
        RECT 2625.750 380.160 2626.070 380.220 ;
        RECT 1642.270 380.020 1642.590 380.080 ;
        RECT 1690.110 380.020 1690.430 380.080 ;
        RECT 1642.270 379.880 1690.430 380.020 ;
        RECT 1642.270 379.820 1642.590 379.880 ;
        RECT 1690.110 379.820 1690.430 379.880 ;
        RECT 1973.470 380.020 1973.790 380.080 ;
        RECT 1994.630 380.020 1994.950 380.080 ;
        RECT 1973.470 379.880 1994.950 380.020 ;
        RECT 1973.470 379.820 1973.790 379.880 ;
        RECT 1994.630 379.820 1994.950 379.880 ;
        RECT 2649.670 380.020 2649.990 380.080 ;
        RECT 2697.510 380.020 2697.830 380.080 ;
        RECT 2649.670 379.880 2697.830 380.020 ;
        RECT 2649.670 379.820 2649.990 379.880 ;
        RECT 2697.510 379.820 2697.830 379.880 ;
      LAYER via ;
        RECT 1457.380 380.500 1457.640 380.760 ;
        RECT 1496.940 380.500 1497.200 380.760 ;
        RECT 2090.340 380.500 2090.600 380.760 ;
        RECT 2124.840 380.500 2125.100 380.760 ;
        RECT 2476.740 380.500 2477.000 380.760 ;
        RECT 2528.720 380.500 2528.980 380.760 ;
        RECT 1799.160 380.160 1799.420 380.420 ;
        RECT 1801.920 380.160 1802.180 380.420 ;
        RECT 2621.640 380.160 2621.900 380.420 ;
        RECT 2625.780 380.160 2626.040 380.420 ;
        RECT 1642.300 379.820 1642.560 380.080 ;
        RECT 1690.140 379.820 1690.400 380.080 ;
        RECT 1973.500 379.820 1973.760 380.080 ;
        RECT 1994.660 379.820 1994.920 380.080 ;
        RECT 2649.700 379.820 2649.960 380.080 ;
        RECT 2697.540 379.820 2697.800 380.080 ;
      LAYER met2 ;
        RECT 1185.510 2496.690 1185.790 2500.000 ;
        RECT 1185.970 2496.690 1186.250 2496.805 ;
        RECT 1185.510 2496.550 1186.250 2496.690 ;
        RECT 1185.510 2496.000 1185.790 2496.550 ;
        RECT 1185.970 2496.435 1186.250 2496.550 ;
        RECT 1562.710 382.315 1562.990 382.685 ;
        RECT 1562.780 381.325 1562.920 382.315 ;
        RECT 2069.170 381.635 2069.450 382.005 ;
        RECT 1496.930 380.955 1497.210 381.325 ;
        RECT 1562.710 380.955 1562.990 381.325 ;
        RECT 1690.130 380.955 1690.410 381.325 ;
        RECT 1497.000 380.790 1497.140 380.955 ;
        RECT 1457.380 380.470 1457.640 380.790 ;
        RECT 1496.940 380.470 1497.200 380.790 ;
        RECT 1457.440 379.965 1457.580 380.470 ;
        RECT 1606.410 380.275 1606.690 380.645 ;
        RECT 1457.370 379.595 1457.650 379.965 ;
        RECT 1606.480 378.605 1606.620 380.275 ;
        RECT 1690.200 380.110 1690.340 380.955 ;
        RECT 1799.150 380.275 1799.430 380.645 ;
        RECT 1801.910 380.275 1802.190 380.645 ;
        RECT 1994.650 380.275 1994.930 380.645 ;
        RECT 1799.160 380.130 1799.420 380.275 ;
        RECT 1801.920 380.130 1802.180 380.275 ;
        RECT 1994.720 380.110 1994.860 380.275 ;
        RECT 1642.300 379.965 1642.560 380.110 ;
        RECT 1642.290 379.595 1642.570 379.965 ;
        RECT 1690.140 379.790 1690.400 380.110 ;
        RECT 1973.500 379.965 1973.760 380.110 ;
        RECT 1973.490 379.595 1973.770 379.965 ;
        RECT 1994.660 379.790 1994.920 380.110 ;
        RECT 2069.240 379.850 2069.380 381.635 ;
        RECT 2124.830 380.955 2125.110 381.325 ;
        RECT 2697.530 380.955 2697.810 381.325 ;
        RECT 2124.900 380.790 2125.040 380.955 ;
        RECT 2090.340 380.645 2090.600 380.790 ;
        RECT 2090.330 380.275 2090.610 380.645 ;
        RECT 2124.840 380.470 2125.100 380.790 ;
        RECT 2476.740 380.645 2477.000 380.790 ;
        RECT 2528.720 380.645 2528.980 380.790 ;
        RECT 2476.730 380.275 2477.010 380.645 ;
        RECT 2528.710 380.275 2528.990 380.645 ;
        RECT 2573.330 380.530 2573.610 380.645 ;
        RECT 2574.250 380.530 2574.530 380.645 ;
        RECT 2573.330 380.390 2574.530 380.530 ;
        RECT 2573.330 380.275 2573.610 380.390 ;
        RECT 2574.250 380.275 2574.530 380.390 ;
        RECT 2621.630 380.275 2621.910 380.645 ;
        RECT 2621.640 380.130 2621.900 380.275 ;
        RECT 2625.780 380.130 2626.040 380.450 ;
        RECT 2625.840 379.965 2625.980 380.130 ;
        RECT 2697.600 380.110 2697.740 380.955 ;
        RECT 2649.700 379.965 2649.960 380.110 ;
        RECT 2069.630 379.850 2069.910 379.965 ;
        RECT 2069.240 379.710 2069.910 379.850 ;
        RECT 2069.630 379.595 2069.910 379.710 ;
        RECT 2625.770 379.595 2626.050 379.965 ;
        RECT 2649.690 379.595 2649.970 379.965 ;
        RECT 2697.540 379.790 2697.800 380.110 ;
        RECT 1606.410 378.235 1606.690 378.605 ;
      LAYER via2 ;
        RECT 1185.970 2496.480 1186.250 2496.760 ;
        RECT 1562.710 382.360 1562.990 382.640 ;
        RECT 2069.170 381.680 2069.450 381.960 ;
        RECT 1496.930 381.000 1497.210 381.280 ;
        RECT 1562.710 381.000 1562.990 381.280 ;
        RECT 1690.130 381.000 1690.410 381.280 ;
        RECT 1606.410 380.320 1606.690 380.600 ;
        RECT 1457.370 379.640 1457.650 379.920 ;
        RECT 1799.150 380.320 1799.430 380.600 ;
        RECT 1801.910 380.320 1802.190 380.600 ;
        RECT 1994.650 380.320 1994.930 380.600 ;
        RECT 1642.290 379.640 1642.570 379.920 ;
        RECT 1973.490 379.640 1973.770 379.920 ;
        RECT 2124.830 381.000 2125.110 381.280 ;
        RECT 2697.530 381.000 2697.810 381.280 ;
        RECT 2090.330 380.320 2090.610 380.600 ;
        RECT 2476.730 380.320 2477.010 380.600 ;
        RECT 2528.710 380.320 2528.990 380.600 ;
        RECT 2573.330 380.320 2573.610 380.600 ;
        RECT 2574.250 380.320 2574.530 380.600 ;
        RECT 2621.630 380.320 2621.910 380.600 ;
        RECT 2069.630 379.640 2069.910 379.920 ;
        RECT 2625.770 379.640 2626.050 379.920 ;
        RECT 2649.690 379.640 2649.970 379.920 ;
        RECT 1606.410 378.280 1606.690 378.560 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 380.540 2924.800 381.740 ;
=======
        RECT 1186.405 2498.140 1186.735 2498.145 ;
        RECT 1186.150 2498.130 1186.735 2498.140 ;
        RECT 1185.950 2497.830 1186.735 2498.130 ;
        RECT 1186.150 2497.820 1186.735 2497.830 ;
        RECT 1186.405 2497.815 1186.735 2497.820 ;
        RECT 1186.150 404.410 1186.530 404.420 ;
        RECT 1200.205 404.410 1200.535 404.425 ;
        RECT 1186.150 404.110 1200.535 404.410 ;
        RECT 1186.150 404.100 1186.530 404.110 ;
        RECT 1200.205 404.095 1200.535 404.110 ;
        RECT 1980.110 382.650 1980.490 382.660 ;
        RECT 2028.205 382.650 2028.535 382.665 ;
        RECT 1980.110 382.350 2028.535 382.650 ;
        RECT 1980.110 382.340 1980.490 382.350 ;
        RECT 2028.205 382.335 2028.535 382.350 ;
        RECT 2052.585 381.970 2052.915 381.985 ;
        RECT 2028.910 381.670 2052.915 381.970 ;
        RECT 1296.805 381.290 1297.135 381.305 ;
        RECT 1399.845 381.290 1400.175 381.305 ;
        RECT 1248.750 380.990 1297.135 381.290 ;
        RECT 1200.205 380.610 1200.535 380.625 ;
        RECT 1200.205 380.310 1225.130 380.610 ;
        RECT 1200.205 380.295 1200.535 380.310 ;
        RECT 1224.830 379.930 1225.130 380.310 ;
        RECT 1248.750 379.930 1249.050 380.990 ;
        RECT 1296.805 380.975 1297.135 380.990 ;
        RECT 1366.510 380.990 1400.175 381.290 ;
        RECT 1224.830 379.630 1249.050 379.930 ;
        RECT 1296.805 379.930 1297.135 379.945 ;
        RECT 1366.510 379.930 1366.810 380.990 ;
        RECT 1399.845 380.975 1400.175 380.990 ;
        RECT 1405.825 381.290 1406.155 381.305 ;
        RECT 1593.045 381.290 1593.375 381.305 ;
        RECT 1405.825 380.990 1593.375 381.290 ;
        RECT 1405.825 380.975 1406.155 380.990 ;
        RECT 1593.045 380.975 1593.375 380.990 ;
        RECT 1946.325 381.290 1946.655 381.305 ;
        RECT 1980.110 381.290 1980.490 381.300 ;
        RECT 1946.325 380.990 1980.490 381.290 ;
        RECT 1946.325 380.975 1946.655 380.990 ;
        RECT 1980.110 380.980 1980.490 380.990 ;
        RECT 1702.065 380.610 1702.395 380.625 ;
        RECT 1656.310 380.310 1702.395 380.610 ;
        RECT 1296.805 379.630 1366.810 379.930 ;
        RECT 1593.045 379.930 1593.375 379.945 ;
        RECT 1656.310 379.930 1656.610 380.310 ;
        RECT 1702.065 380.295 1702.395 380.310 ;
        RECT 1711.725 380.610 1712.055 380.625 ;
        RECT 1798.665 380.610 1798.995 380.625 ;
        RECT 1711.725 380.310 1738.490 380.610 ;
        RECT 1711.725 380.295 1712.055 380.310 ;
        RECT 1593.045 379.630 1656.610 379.930 ;
        RECT 1738.190 379.930 1738.490 380.310 ;
        RECT 1752.910 380.310 1798.995 380.610 ;
=======
        RECT 1185.945 2496.780 1186.275 2496.785 ;
        RECT 1185.945 2496.770 1186.530 2496.780 ;
        RECT 1185.945 2496.470 1186.730 2496.770 ;
        RECT 1185.945 2496.460 1186.530 2496.470 ;
        RECT 1185.945 2496.455 1186.275 2496.460 ;
        RECT 1538.510 382.650 1538.890 382.660 ;
        RECT 1562.685 382.650 1563.015 382.665 ;
        RECT 1538.510 382.350 1563.015 382.650 ;
        RECT 1538.510 382.340 1538.890 382.350 ;
        RECT 1562.685 382.335 1563.015 382.350 ;
        RECT 2069.145 381.970 2069.475 381.985 ;
        RECT 2021.550 381.670 2069.475 381.970 ;
        RECT 1496.905 381.290 1497.235 381.305 ;
        RECT 1538.510 381.290 1538.890 381.300 ;
        RECT 1266.230 380.990 1318.970 381.290 ;
        RECT 1186.150 380.610 1186.530 380.620 ;
        RECT 1266.230 380.610 1266.530 380.990 ;
        RECT 1186.150 380.310 1200.290 380.610 ;
        RECT 1186.150 380.300 1186.530 380.310 ;
        RECT 1199.990 379.930 1200.290 380.310 ;
        RECT 1225.750 380.310 1266.530 380.610 ;
        RECT 1225.750 379.930 1226.050 380.310 ;
        RECT 1199.990 379.630 1226.050 379.930 ;
        RECT 1318.670 379.930 1318.970 380.990 ;
        RECT 1496.905 380.990 1538.890 381.290 ;
        RECT 1496.905 380.975 1497.235 380.990 ;
        RECT 1538.510 380.980 1538.890 380.990 ;
        RECT 1562.685 381.290 1563.015 381.305 ;
        RECT 1690.105 381.290 1690.435 381.305 ;
        RECT 1924.910 381.290 1925.290 381.300 ;
        RECT 1562.685 380.990 1586.690 381.290 ;
        RECT 1562.685 380.975 1563.015 380.990 ;
        RECT 1586.390 380.610 1586.690 380.990 ;
        RECT 1690.105 380.990 1704.450 381.290 ;
        RECT 1690.105 380.975 1690.435 380.990 ;
        RECT 1606.385 380.610 1606.715 380.625 ;
        RECT 1586.390 380.310 1606.715 380.610 ;
        RECT 1606.385 380.295 1606.715 380.310 ;
        RECT 1457.345 379.930 1457.675 379.945 ;
        RECT 1642.265 379.930 1642.595 379.945 ;
        RECT 1318.670 379.630 1457.675 379.930 ;
        RECT 1457.345 379.615 1457.675 379.630 ;
        RECT 1641.590 379.630 1642.595 379.930 ;
        RECT 1704.150 379.930 1704.450 380.990 ;
        RECT 1849.510 380.990 1925.290 381.290 ;
        RECT 1799.125 380.610 1799.455 380.625 ;
        RECT 1752.910 380.310 1799.455 380.610 ;
>>>>>>> re-updated local openlane
        RECT 1752.910 379.930 1753.210 380.310 ;
        RECT 1799.125 380.295 1799.455 380.310 ;
        RECT 1801.885 380.610 1802.215 380.625 ;
        RECT 1801.885 380.310 1835.090 380.610 ;
        RECT 1801.885 380.295 1802.215 380.310 ;
        RECT 1704.150 379.630 1753.210 379.930 ;
        RECT 1834.790 379.930 1835.090 380.310 ;
        RECT 1849.510 379.930 1849.810 380.990 ;
        RECT 1924.910 380.980 1925.290 380.990 ;
        RECT 1994.625 380.610 1994.955 380.625 ;
        RECT 2021.550 380.610 2021.850 381.670 ;
        RECT 2069.145 381.655 2069.475 381.670 ;
        RECT 2124.805 381.290 2125.135 381.305 ;
        RECT 2697.505 381.290 2697.835 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2124.805 380.990 2235.290 381.290 ;
        RECT 2124.805 380.975 2125.135 380.990 ;
        RECT 2090.305 380.610 2090.635 380.625 ;
        RECT 1994.625 380.310 2021.850 380.610 ;
        RECT 2076.750 380.310 2090.635 380.610 ;
        RECT 1994.625 380.295 1994.955 380.310 ;
        RECT 1834.790 379.630 1849.810 379.930 ;
        RECT 1924.910 379.930 1925.290 379.940 ;
        RECT 1973.465 379.930 1973.795 379.945 ;
        RECT 1924.910 379.630 1973.795 379.930 ;
        RECT 1606.385 378.570 1606.715 378.585 ;
        RECT 1641.590 378.570 1641.890 379.630 ;
        RECT 1642.265 379.615 1642.595 379.630 ;
        RECT 1924.910 379.620 1925.290 379.630 ;
        RECT 1973.465 379.615 1973.795 379.630 ;
        RECT 2069.605 379.930 2069.935 379.945 ;
        RECT 2076.750 379.930 2077.050 380.310 ;
        RECT 2090.305 380.295 2090.635 380.310 ;
        RECT 2069.605 379.630 2077.050 379.930 ;
        RECT 2069.605 379.615 2069.935 379.630 ;
        RECT 2234.990 379.250 2235.290 380.990 ;
        RECT 2304.910 380.990 2353.050 381.290 ;
        RECT 2304.910 379.930 2305.210 380.990 ;
        RECT 2352.750 380.610 2353.050 380.990 ;
        RECT 2401.510 380.990 2429.410 381.290 ;
        RECT 2352.750 380.310 2400.890 380.610 ;
        RECT 2269.950 379.630 2305.210 379.930 ;
        RECT 2400.590 379.930 2400.890 380.310 ;
        RECT 2401.510 379.930 2401.810 380.990 ;
        RECT 2429.110 380.610 2429.410 380.990 ;
        RECT 2697.505 380.990 2739.450 381.290 ;
        RECT 2697.505 380.975 2697.835 380.990 ;
        RECT 2476.705 380.610 2477.035 380.625 ;
        RECT 2429.110 380.310 2477.035 380.610 ;
        RECT 2476.705 380.295 2477.035 380.310 ;
        RECT 2528.685 380.610 2529.015 380.625 ;
        RECT 2573.305 380.610 2573.635 380.625 ;
        RECT 2528.685 380.310 2573.635 380.610 ;
        RECT 2528.685 380.295 2529.015 380.310 ;
        RECT 2573.305 380.295 2573.635 380.310 ;
        RECT 2574.225 380.610 2574.555 380.625 ;
        RECT 2621.605 380.610 2621.935 380.625 ;
        RECT 2574.225 380.310 2621.935 380.610 ;
        RECT 2739.150 380.610 2739.450 380.990 ;
        RECT 2787.910 380.990 2836.050 381.290 ;
        RECT 2739.150 380.310 2787.290 380.610 ;
        RECT 2574.225 380.295 2574.555 380.310 ;
        RECT 2621.605 380.295 2621.935 380.310 ;
        RECT 2400.590 379.630 2401.810 379.930 ;
        RECT 2625.745 379.930 2626.075 379.945 ;
        RECT 2649.665 379.930 2649.995 379.945 ;
        RECT 2625.745 379.630 2649.995 379.930 ;
        RECT 2786.990 379.930 2787.290 380.310 ;
        RECT 2787.910 379.930 2788.210 380.990 ;
        RECT 2835.750 380.610 2836.050 380.990 ;
        RECT 2916.710 380.990 2924.800 381.290 ;
        RECT 2916.710 380.610 2917.010 380.990 ;
        RECT 2835.750 380.310 2883.890 380.610 ;
        RECT 2786.990 379.630 2788.210 379.930 ;
        RECT 2883.590 379.930 2883.890 380.310 ;
        RECT 2884.510 380.310 2917.010 380.610 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2884.510 379.930 2884.810 380.310 ;
        RECT 2883.590 379.630 2884.810 379.930 ;
        RECT 2269.950 379.250 2270.250 379.630 ;
        RECT 2625.745 379.615 2626.075 379.630 ;
        RECT 2649.665 379.615 2649.995 379.630 ;
        RECT 2234.990 378.950 2270.250 379.250 ;
        RECT 1606.385 378.270 1641.890 378.570 ;
        RECT 1606.385 378.255 1606.715 378.270 ;
      LAYER via3 ;
        RECT 1186.180 2496.460 1186.500 2496.780 ;
        RECT 1538.540 382.340 1538.860 382.660 ;
        RECT 1186.180 380.300 1186.500 380.620 ;
        RECT 1538.540 380.980 1538.860 381.300 ;
        RECT 1924.940 380.980 1925.260 381.300 ;
        RECT 1924.940 379.620 1925.260 379.940 ;
      LAYER met4 ;
<<<<<<< HEAD
        RECT 1186.175 2497.815 1186.505 2498.145 ;
        RECT 1186.190 404.425 1186.490 2497.815 ;
        RECT 1186.175 404.095 1186.505 404.425 ;
        RECT 1980.135 382.335 1980.465 382.665 ;
        RECT 1980.150 381.305 1980.450 382.335 ;
        RECT 1980.135 380.975 1980.465 381.305 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1186.175 2496.455 1186.505 2496.785 ;
        RECT 1186.190 380.625 1186.490 2496.455 ;
        RECT 1538.535 382.335 1538.865 382.665 ;
        RECT 1538.550 381.305 1538.850 382.335 ;
        RECT 1538.535 380.975 1538.865 381.305 ;
        RECT 1924.935 380.975 1925.265 381.305 ;
        RECT 1186.175 380.295 1186.505 380.625 ;
        RECT 1924.950 379.945 1925.250 380.975 ;
        RECT 1924.935 379.615 1925.265 379.945 ;
>>>>>>> re-updated local openlane
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3499.860 1095.190 3499.920 ;
        RECT 1552.570 3499.860 1552.890 3499.920 ;
        RECT 1094.870 3499.720 1552.890 3499.860 ;
        RECT 1094.870 3499.660 1095.190 3499.720 ;
        RECT 1552.570 3499.660 1552.890 3499.720 ;
      LAYER via ;
        RECT 1094.900 3499.660 1095.160 3499.920 ;
        RECT 1552.600 3499.660 1552.860 3499.920 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1094.750 3519.700 1095.310 3524.800 ;
=======
        RECT 1094.750 3517.600 1095.310 3524.800 ;
<<<<<<< HEAD
        RECT 1094.960 3500.630 1095.100 3517.600 ;
        RECT 1094.900 3500.310 1095.160 3500.630 ;
        RECT 1542.020 3500.310 1542.280 3500.630 ;
        RECT 1542.080 2517.690 1542.220 3500.310 ;
        RECT 1563.180 2517.710 1563.440 2518.030 ;
        RECT 1542.020 2517.370 1542.280 2517.690 ;
        RECT 1563.240 2500.000 1563.380 2517.710 ;
        RECT 1563.170 2496.000 1563.450 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1094.960 3499.950 1095.100 3517.600 ;
        RECT 1094.900 3499.630 1095.160 3499.950 ;
        RECT 1552.600 3499.630 1552.860 3499.950 ;
        RECT 1552.660 2499.410 1552.800 3499.630 ;
        RECT 1553.050 2499.410 1553.330 2500.000 ;
        RECT 1552.660 2499.270 1553.330 2499.410 ;
        RECT 1553.050 2496.000 1553.330 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 770.570 3504.960 770.890 3505.020 ;
        RECT 1566.370 3504.960 1566.690 3505.020 ;
        RECT 770.570 3504.820 1566.690 3504.960 ;
        RECT 770.570 3504.760 770.890 3504.820 ;
        RECT 1566.370 3504.760 1566.690 3504.820 ;
      LAYER via ;
        RECT 770.600 3504.760 770.860 3505.020 ;
        RECT 1566.400 3504.760 1566.660 3505.020 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 770.450 3519.700 771.010 3524.800 ;
=======
        RECT 770.450 3517.600 771.010 3524.800 ;
<<<<<<< HEAD
        RECT 770.660 3504.710 770.800 3517.600 ;
        RECT 770.600 3504.390 770.860 3504.710 ;
        RECT 1562.720 3504.390 1562.980 3504.710 ;
        RECT 1562.780 2518.450 1562.920 3504.390 ;
        RECT 1562.780 2518.310 1563.840 2518.450 ;
        RECT 1563.700 2517.770 1563.840 2518.310 ;
        RECT 1564.560 2518.050 1564.820 2518.370 ;
        RECT 1582.960 2518.050 1583.220 2518.370 ;
        RECT 1564.620 2517.770 1564.760 2518.050 ;
        RECT 1563.700 2517.630 1564.760 2517.770 ;
        RECT 1583.020 2500.000 1583.160 2518.050 ;
        RECT 1582.950 2496.000 1583.230 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 770.660 3505.050 770.800 3517.600 ;
        RECT 770.600 3504.730 770.860 3505.050 ;
        RECT 1566.400 3504.730 1566.660 3505.050 ;
        RECT 1566.460 2500.090 1566.600 3504.730 ;
        RECT 1566.460 2499.950 1570.280 2500.090 ;
        RECT 1570.140 2499.410 1570.280 2499.950 ;
        RECT 1572.370 2499.410 1572.650 2500.000 ;
        RECT 1570.140 2499.270 1572.650 2499.410 ;
        RECT 1572.370 2496.000 1572.650 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.810 3503.260 446.130 3503.320 ;
        RECT 1587.070 3503.260 1587.390 3503.320 ;
        RECT 445.810 3503.120 1587.390 3503.260 ;
        RECT 445.810 3503.060 446.130 3503.120 ;
        RECT 1587.070 3503.060 1587.390 3503.120 ;
      LAYER via ;
        RECT 445.840 3503.060 446.100 3503.320 ;
        RECT 1587.100 3503.060 1587.360 3503.320 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 445.690 3519.700 446.250 3524.800 ;
=======
        RECT 445.690 3517.600 446.250 3524.800 ;
<<<<<<< HEAD
        RECT 445.900 3503.010 446.040 3517.600 ;
        RECT 445.840 3502.690 446.100 3503.010 ;
        RECT 1583.420 3502.690 1583.680 3503.010 ;
        RECT 1583.480 2518.370 1583.620 3502.690 ;
        RECT 1583.420 2518.050 1583.680 2518.370 ;
        RECT 1602.740 2518.050 1603.000 2518.370 ;
        RECT 1602.800 2500.000 1602.940 2518.050 ;
        RECT 1602.730 2496.000 1603.010 2500.000 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 445.900 3503.350 446.040 3517.600 ;
        RECT 445.840 3503.030 446.100 3503.350 ;
        RECT 1587.100 3503.030 1587.360 3503.350 ;
        RECT 1587.160 2500.770 1587.300 3503.030 ;
        RECT 1587.160 2500.630 1589.600 2500.770 ;
        RECT 1589.460 2499.410 1589.600 2500.630 ;
        RECT 1591.690 2499.410 1591.970 2500.000 ;
        RECT 1589.460 2499.270 1591.970 2499.410 ;
        RECT 1591.690 2496.000 1591.970 2499.270 ;
>>>>>>> re-updated local openlane
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 1607.770 3501.560 1608.090 3501.620 ;
        RECT 121.510 3501.420 1608.090 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 1607.770 3501.360 1608.090 3501.420 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 1607.800 3501.360 1608.060 3501.620 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 121.390 3519.700 121.950 3524.800 ;
=======
        RECT 121.390 3517.600 121.950 3524.800 ;
<<<<<<< HEAD
        RECT 121.600 3502.525 121.740 3517.600 ;
        RECT 121.530 3502.155 121.810 3502.525 ;
        RECT 1604.110 3502.155 1604.390 3502.525 ;
        RECT 1604.180 2518.370 1604.320 3502.155 ;
        RECT 1604.120 2518.050 1604.380 2518.370 ;
        RECT 1622.520 2518.050 1622.780 2518.370 ;
        RECT 1622.580 2500.000 1622.720 2518.050 ;
        RECT 1622.510 2496.000 1622.790 2500.000 ;
      LAYER via2 ;
        RECT 121.530 3502.200 121.810 3502.480 ;
        RECT 1604.110 3502.200 1604.390 3502.480 ;
      LAYER met3 ;
        RECT 121.505 3502.490 121.835 3502.505 ;
        RECT 1604.085 3502.490 1604.415 3502.505 ;
        RECT 121.505 3502.190 1604.415 3502.490 ;
        RECT 121.505 3502.175 121.835 3502.190 ;
        RECT 1604.085 3502.175 1604.415 3502.190 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 1607.800 3501.330 1608.060 3501.650 ;
        RECT 1607.860 2499.410 1608.000 3501.330 ;
        RECT 1607.860 2499.270 1608.460 2499.410 ;
        RECT 1608.320 2498.730 1608.460 2499.270 ;
        RECT 1611.010 2498.730 1611.290 2500.000 ;
        RECT 1608.320 2498.590 1611.290 2498.730 ;
        RECT 1611.010 2496.000 1611.290 2498.590 ;
>>>>>>> re-updated local openlane
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 1628.470 3339.720 1628.790 3339.780 ;
        RECT 17.090 3339.580 1628.790 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 1628.470 3339.520 1628.790 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 1628.500 3339.520 1628.760 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 1628.500 3339.490 1628.760 3339.810 ;
        RECT 1628.560 2499.410 1628.700 3339.490 ;
        RECT 1630.330 2499.410 1630.610 2500.000 ;
        RECT 1628.560 2499.270 1630.610 2499.410 ;
        RECT 1630.330 2496.000 1630.610 2499.270 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3339.220 0.300 3340.420 ;
=======
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 3050.040 16.950 3050.100 ;
        RECT 1649.170 3050.040 1649.490 3050.100 ;
        RECT 16.630 3049.900 1649.490 3050.040 ;
        RECT 16.630 3049.840 16.950 3049.900 ;
        RECT 1649.170 3049.840 1649.490 3049.900 ;
      LAYER via ;
        RECT 16.660 3049.840 16.920 3050.100 ;
        RECT 1649.200 3049.840 1649.460 3050.100 ;
      LAYER met2 ;
        RECT 16.650 3051.995 16.930 3052.365 ;
        RECT 16.720 3050.130 16.860 3051.995 ;
        RECT 16.660 3049.810 16.920 3050.130 ;
        RECT 1649.200 3049.810 1649.460 3050.130 ;
        RECT 1649.260 2499.410 1649.400 3049.810 ;
        RECT 1649.650 2499.410 1649.930 2500.000 ;
        RECT 1649.260 2499.270 1649.930 2499.410 ;
        RECT 1649.650 2496.000 1649.930 2499.270 ;
      LAYER via2 ;
        RECT 16.650 3052.040 16.930 3052.320 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3051.580 0.300 3052.780 ;
=======
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 16.625 3052.330 16.955 3052.345 ;
        RECT -4.800 3052.030 16.955 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
<<<<<<< HEAD
        RECT 17.085 3052.015 17.415 3052.030 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 3052.015 16.955 3052.030 ;
>>>>>>> re-updated local openlane
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2760.360 16.950 2760.420 ;
        RECT 1662.970 2760.360 1663.290 2760.420 ;
        RECT 16.630 2760.220 1663.290 2760.360 ;
        RECT 16.630 2760.160 16.950 2760.220 ;
        RECT 1662.970 2760.160 1663.290 2760.220 ;
      LAYER via ;
        RECT 16.660 2760.160 16.920 2760.420 ;
        RECT 1663.000 2760.160 1663.260 2760.420 ;
      LAYER met2 ;
        RECT 16.650 2765.035 16.930 2765.405 ;
        RECT 16.720 2760.450 16.860 2765.035 ;
        RECT 16.660 2760.130 16.920 2760.450 ;
        RECT 1663.000 2760.130 1663.260 2760.450 ;
        RECT 1663.060 2500.090 1663.200 2760.130 ;
        RECT 1663.060 2499.950 1667.340 2500.090 ;
        RECT 1667.200 2499.410 1667.340 2499.950 ;
        RECT 1668.970 2499.410 1669.250 2500.000 ;
        RECT 1667.200 2499.270 1669.250 2499.410 ;
        RECT 1668.970 2496.000 1669.250 2499.270 ;
      LAYER via2 ;
        RECT 16.650 2765.080 16.930 2765.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2764.620 0.300 2765.820 ;
=======
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 16.625 2765.370 16.955 2765.385 ;
        RECT -4.800 2765.070 16.955 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
<<<<<<< HEAD
        RECT 15.705 2765.055 16.035 2765.070 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 2765.055 16.955 2765.070 ;
>>>>>>> re-updated local openlane
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1687.425 2491.945 1687.595 2497.215 ;
      LAYER mcon ;
        RECT 1687.425 2497.045 1687.595 2497.215 ;
      LAYER met1 ;
        RECT 1687.350 2497.200 1687.670 2497.260 ;
        RECT 1687.155 2497.060 1687.670 2497.200 ;
        RECT 1687.350 2497.000 1687.670 2497.060 ;
        RECT 15.710 2492.100 16.030 2492.160 ;
        RECT 1687.365 2492.100 1687.655 2492.145 ;
        RECT 15.710 2491.960 1687.655 2492.100 ;
        RECT 15.710 2491.900 16.030 2491.960 ;
        RECT 1687.365 2491.915 1687.655 2491.960 ;
      LAYER via ;
        RECT 1687.380 2497.000 1687.640 2497.260 ;
        RECT 15.740 2491.900 16.000 2492.160 ;
      LAYER met2 ;
        RECT 1688.750 2497.370 1689.030 2500.000 ;
        RECT 1687.440 2497.290 1689.030 2497.370 ;
        RECT 1687.380 2497.230 1689.030 2497.290 ;
        RECT 1687.380 2496.970 1687.640 2497.230 ;
        RECT 1688.750 2496.000 1689.030 2497.230 ;
        RECT 15.740 2491.870 16.000 2492.190 ;
        RECT 15.800 2477.765 15.940 2491.870 ;
        RECT 15.730 2477.395 16.010 2477.765 ;
      LAYER via2 ;
        RECT 15.730 2477.440 16.010 2477.720 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2476.980 0.300 2478.180 ;
=======
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 15.705 2477.730 16.035 2477.745 ;
        RECT -4.800 2477.430 16.035 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
<<<<<<< HEAD
        RECT 13.865 2477.415 14.195 2477.430 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 15.705 2477.415 16.035 2477.430 ;
>>>>>>> re-updated local openlane
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.890 2512.160 31.210 2512.220 ;
        RECT 1708.050 2512.160 1708.370 2512.220 ;
        RECT 30.890 2512.020 1708.370 2512.160 ;
        RECT 30.890 2511.960 31.210 2512.020 ;
        RECT 1708.050 2511.960 1708.370 2512.020 ;
        RECT 13.870 2191.880 14.190 2191.940 ;
        RECT 30.890 2191.880 31.210 2191.940 ;
        RECT 13.870 2191.740 31.210 2191.880 ;
        RECT 13.870 2191.680 14.190 2191.740 ;
        RECT 30.890 2191.680 31.210 2191.740 ;
      LAYER via ;
        RECT 30.920 2511.960 31.180 2512.220 ;
        RECT 1708.080 2511.960 1708.340 2512.220 ;
        RECT 13.900 2191.680 14.160 2191.940 ;
        RECT 30.920 2191.680 31.180 2191.940 ;
      LAYER met2 ;
        RECT 30.920 2511.930 31.180 2512.250 ;
        RECT 1708.080 2511.930 1708.340 2512.250 ;
        RECT 30.980 2191.970 31.120 2511.930 ;
        RECT 1708.140 2500.000 1708.280 2511.930 ;
        RECT 1708.070 2496.000 1708.350 2500.000 ;
        RECT 13.900 2191.650 14.160 2191.970 ;
        RECT 30.920 2191.650 31.180 2191.970 ;
        RECT 13.960 2190.125 14.100 2191.650 ;
        RECT 13.890 2189.755 14.170 2190.125 ;
      LAYER via2 ;
        RECT 13.890 2189.800 14.170 2190.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2189.340 0.300 2190.540 ;
=======
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 13.865 2190.090 14.195 2190.105 ;
        RECT -4.800 2189.790 14.195 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 13.865 2189.775 14.195 2189.790 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 79.190 2512.840 79.510 2512.900 ;
        RECT 1727.370 2512.840 1727.690 2512.900 ;
        RECT 79.190 2512.700 1727.690 2512.840 ;
        RECT 79.190 2512.640 79.510 2512.700 ;
        RECT 1727.370 2512.640 1727.690 2512.700 ;
        RECT 16.630 1904.240 16.950 1904.300 ;
        RECT 79.190 1904.240 79.510 1904.300 ;
        RECT 16.630 1904.100 79.510 1904.240 ;
        RECT 16.630 1904.040 16.950 1904.100 ;
        RECT 79.190 1904.040 79.510 1904.100 ;
      LAYER via ;
        RECT 79.220 2512.640 79.480 2512.900 ;
        RECT 1727.400 2512.640 1727.660 2512.900 ;
        RECT 16.660 1904.040 16.920 1904.300 ;
        RECT 79.220 1904.040 79.480 1904.300 ;
      LAYER met2 ;
        RECT 79.220 2512.610 79.480 2512.930 ;
        RECT 1727.400 2512.610 1727.660 2512.930 ;
        RECT 79.280 1904.330 79.420 2512.610 ;
        RECT 1727.460 2500.000 1727.600 2512.610 ;
        RECT 1727.390 2496.000 1727.670 2500.000 ;
        RECT 16.660 1904.010 16.920 1904.330 ;
        RECT 79.220 1904.010 79.480 1904.330 ;
        RECT 16.720 1903.165 16.860 1904.010 ;
        RECT 16.650 1902.795 16.930 1903.165 ;
      LAYER via2 ;
        RECT 16.650 1902.840 16.930 1903.120 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1902.380 0.300 1903.580 ;
=======
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.625 1903.130 16.955 1903.145 ;
        RECT -4.800 1902.830 16.955 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
<<<<<<< HEAD
        RECT 15.245 1902.815 15.575 1902.830 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 1902.815 16.955 1902.830 ;
>>>>>>> re-updated local openlane
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2456.470 615.300 2456.790 615.360 ;
        RECT 2504.310 615.300 2504.630 615.360 ;
        RECT 2456.470 615.160 2504.630 615.300 ;
        RECT 2456.470 615.100 2456.790 615.160 ;
        RECT 2504.310 615.100 2504.630 615.160 ;
        RECT 1799.130 614.960 1799.450 615.020 ;
        RECT 1801.890 614.960 1802.210 615.020 ;
        RECT 1799.130 614.820 1802.210 614.960 ;
        RECT 1799.130 614.760 1799.450 614.820 ;
        RECT 1801.890 614.760 1802.210 614.820 ;
        RECT 2621.610 614.960 2621.930 615.020 ;
        RECT 2622.530 614.960 2622.850 615.020 ;
        RECT 2621.610 614.820 2622.850 614.960 ;
        RECT 2621.610 614.760 2621.930 614.820 ;
        RECT 2622.530 614.760 2622.850 614.820 ;
        RECT 1642.270 614.620 1642.590 614.680 ;
        RECT 1690.110 614.620 1690.430 614.680 ;
        RECT 1642.270 614.480 1690.430 614.620 ;
        RECT 1642.270 614.420 1642.590 614.480 ;
        RECT 1690.110 614.420 1690.430 614.480 ;
        RECT 2070.070 614.620 2070.390 614.680 ;
        RECT 2117.910 614.620 2118.230 614.680 ;
        RECT 2070.070 614.480 2118.230 614.620 ;
        RECT 2070.070 614.420 2070.390 614.480 ;
        RECT 2117.910 614.420 2118.230 614.480 ;
        RECT 2649.670 614.620 2649.990 614.680 ;
        RECT 2697.510 614.620 2697.830 614.680 ;
        RECT 2649.670 614.480 2697.830 614.620 ;
        RECT 2649.670 614.420 2649.990 614.480 ;
        RECT 2697.510 614.420 2697.830 614.480 ;
        RECT 1959.670 614.280 1959.990 614.340 ;
        RECT 2007.510 614.280 2007.830 614.340 ;
        RECT 1959.670 614.140 2007.830 614.280 ;
        RECT 1959.670 614.080 1959.990 614.140 ;
        RECT 2007.510 614.080 2007.830 614.140 ;
        RECT 2021.310 613.260 2021.630 613.320 ;
        RECT 2055.810 613.260 2056.130 613.320 ;
        RECT 2021.310 613.120 2056.130 613.260 ;
        RECT 2021.310 613.060 2021.630 613.120 ;
        RECT 2055.810 613.060 2056.130 613.120 ;
      LAYER via ;
        RECT 2456.500 615.100 2456.760 615.360 ;
        RECT 2504.340 615.100 2504.600 615.360 ;
        RECT 1799.160 614.760 1799.420 615.020 ;
        RECT 1801.920 614.760 1802.180 615.020 ;
        RECT 2621.640 614.760 2621.900 615.020 ;
        RECT 2622.560 614.760 2622.820 615.020 ;
        RECT 1642.300 614.420 1642.560 614.680 ;
        RECT 1690.140 614.420 1690.400 614.680 ;
        RECT 2070.100 614.420 2070.360 614.680 ;
        RECT 2117.940 614.420 2118.200 614.680 ;
        RECT 2649.700 614.420 2649.960 614.680 ;
        RECT 2697.540 614.420 2697.800 614.680 ;
        RECT 1959.700 614.080 1959.960 614.340 ;
        RECT 2007.540 614.080 2007.800 614.340 ;
        RECT 2021.340 613.060 2021.600 613.320 ;
        RECT 2055.840 613.060 2056.100 613.320 ;
      LAYER met2 ;
        RECT 1204.830 2498.050 1205.110 2500.000 ;
        RECT 1206.210 2498.050 1206.490 2498.165 ;
        RECT 1204.830 2497.910 1206.490 2498.050 ;
        RECT 1204.830 2496.000 1205.110 2497.910 ;
        RECT 1206.210 2497.795 1206.490 2497.910 ;
        RECT 2294.110 616.915 2294.390 617.285 ;
        RECT 2186.930 616.490 2187.210 616.605 ;
        RECT 2187.850 616.490 2188.130 616.605 ;
        RECT 2186.930 616.350 2188.130 616.490 ;
        RECT 2186.930 616.235 2187.210 616.350 ;
        RECT 2187.850 616.235 2188.130 616.350 ;
        RECT 2294.180 615.925 2294.320 616.915 ;
        RECT 1424.710 615.555 1424.990 615.925 ;
        RECT 1690.130 615.555 1690.410 615.925 ;
        RECT 2117.930 615.555 2118.210 615.925 ;
        RECT 2294.110 615.555 2294.390 615.925 ;
        RECT 2504.330 615.555 2504.610 615.925 ;
        RECT 2697.530 615.555 2697.810 615.925 ;
        RECT 1424.780 614.565 1424.920 615.555 ;
        RECT 1606.410 614.875 1606.690 615.245 ;
        RECT 1424.710 614.195 1424.990 614.565 ;
        RECT 1606.480 613.205 1606.620 614.875 ;
        RECT 1690.200 614.710 1690.340 615.555 ;
        RECT 1799.150 614.875 1799.430 615.245 ;
        RECT 1801.910 614.875 1802.190 615.245 ;
        RECT 1799.160 614.730 1799.420 614.875 ;
        RECT 1801.920 614.730 1802.180 614.875 ;
        RECT 2118.000 614.710 2118.140 615.555 ;
        RECT 2504.400 615.390 2504.540 615.555 ;
        RECT 2456.500 615.245 2456.760 615.390 ;
        RECT 2456.490 614.875 2456.770 615.245 ;
        RECT 2504.340 615.070 2504.600 615.390 ;
        RECT 2574.250 615.130 2574.530 615.245 ;
        RECT 2573.400 614.990 2574.530 615.130 ;
        RECT 1642.300 614.565 1642.560 614.710 ;
        RECT 1642.290 614.195 1642.570 614.565 ;
        RECT 1690.140 614.390 1690.400 614.710 ;
        RECT 2070.100 614.565 2070.360 614.710 ;
        RECT 1959.690 614.195 1959.970 614.565 ;
        RECT 1959.700 614.050 1959.960 614.195 ;
        RECT 2007.540 614.050 2007.800 614.370 ;
        RECT 2055.830 614.195 2056.110 614.565 ;
        RECT 2070.090 614.195 2070.370 614.565 ;
        RECT 2117.940 614.390 2118.200 614.710 ;
        RECT 2573.400 614.565 2573.540 614.990 ;
        RECT 2574.250 614.875 2574.530 614.990 ;
        RECT 2621.630 614.875 2621.910 615.245 ;
        RECT 2621.640 614.730 2621.900 614.875 ;
        RECT 2622.560 614.730 2622.820 615.050 ;
        RECT 2622.620 614.565 2622.760 614.730 ;
        RECT 2697.600 614.710 2697.740 615.555 ;
        RECT 2649.700 614.565 2649.960 614.710 ;
        RECT 2573.330 614.195 2573.610 614.565 ;
        RECT 2622.550 614.195 2622.830 614.565 ;
        RECT 2649.690 614.195 2649.970 614.565 ;
        RECT 2697.540 614.390 2697.800 614.710 ;
        RECT 2007.600 613.885 2007.740 614.050 ;
        RECT 2007.530 613.515 2007.810 613.885 ;
        RECT 2055.900 613.350 2056.040 614.195 ;
        RECT 2021.340 613.205 2021.600 613.350 ;
        RECT 1606.410 612.835 1606.690 613.205 ;
        RECT 2021.330 612.835 2021.610 613.205 ;
        RECT 2055.840 613.030 2056.100 613.350 ;
      LAYER via2 ;
        RECT 1206.210 2497.840 1206.490 2498.120 ;
        RECT 2294.110 616.960 2294.390 617.240 ;
        RECT 2186.930 616.280 2187.210 616.560 ;
        RECT 2187.850 616.280 2188.130 616.560 ;
        RECT 1424.710 615.600 1424.990 615.880 ;
        RECT 1690.130 615.600 1690.410 615.880 ;
        RECT 2117.930 615.600 2118.210 615.880 ;
        RECT 2294.110 615.600 2294.390 615.880 ;
        RECT 2504.330 615.600 2504.610 615.880 ;
        RECT 2697.530 615.600 2697.810 615.880 ;
        RECT 1606.410 614.920 1606.690 615.200 ;
        RECT 1424.710 614.240 1424.990 614.520 ;
        RECT 1799.150 614.920 1799.430 615.200 ;
        RECT 1801.910 614.920 1802.190 615.200 ;
        RECT 2456.490 614.920 2456.770 615.200 ;
        RECT 1642.290 614.240 1642.570 614.520 ;
        RECT 1959.690 614.240 1959.970 614.520 ;
        RECT 2055.830 614.240 2056.110 614.520 ;
        RECT 2070.090 614.240 2070.370 614.520 ;
        RECT 2574.250 614.920 2574.530 615.200 ;
        RECT 2621.630 614.920 2621.910 615.200 ;
        RECT 2573.330 614.240 2573.610 614.520 ;
        RECT 2622.550 614.240 2622.830 614.520 ;
        RECT 2649.690 614.240 2649.970 614.520 ;
        RECT 2007.530 613.560 2007.810 613.840 ;
        RECT 1606.410 612.880 1606.690 613.160 ;
        RECT 2021.330 612.880 2021.610 613.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 615.140 2924.800 616.340 ;
=======
        RECT 1206.185 2498.140 1206.515 2498.145 ;
        RECT 1206.185 2498.130 1206.770 2498.140 ;
        RECT 1206.185 2497.830 1206.970 2498.130 ;
        RECT 1206.185 2497.820 1206.770 2497.830 ;
        RECT 1206.185 2497.815 1206.515 2497.820 ;
        RECT 2269.910 617.250 2270.290 617.260 ;
        RECT 2294.085 617.250 2294.415 617.265 ;
        RECT 2269.910 616.950 2294.415 617.250 ;
        RECT 2269.910 616.940 2270.290 616.950 ;
        RECT 2294.085 616.935 2294.415 616.950 ;
        RECT 2173.310 616.570 2173.690 616.580 ;
        RECT 2186.905 616.570 2187.235 616.585 ;
        RECT 1268.990 616.270 1318.970 616.570 ;
        RECT 1206.390 615.210 1206.770 615.220 ;
        RECT 1268.990 615.210 1269.290 616.270 ;
        RECT 1206.390 614.910 1269.290 615.210 ;
        RECT 1318.670 615.210 1318.970 616.270 ;
        RECT 2173.310 616.270 2187.235 616.570 ;
        RECT 2173.310 616.260 2173.690 616.270 ;
        RECT 2186.905 616.255 2187.235 616.270 ;
        RECT 2187.825 616.570 2188.155 616.585 ;
        RECT 2187.825 616.270 2236.210 616.570 ;
        RECT 2187.825 616.255 2188.155 616.270 ;
        RECT 1424.685 615.890 1425.015 615.905 ;
        RECT 1369.270 615.590 1425.015 615.890 ;
        RECT 1369.270 615.210 1369.570 615.590 ;
        RECT 1424.685 615.575 1425.015 615.590 ;
        RECT 1441.910 615.890 1442.290 615.900 ;
        RECT 1690.105 615.890 1690.435 615.905 ;
        RECT 1911.110 615.890 1911.490 615.900 ;
        RECT 1441.910 615.590 1511.250 615.890 ;
        RECT 1441.910 615.580 1442.290 615.590 ;
        RECT 1318.670 614.910 1369.570 615.210 ;
        RECT 1206.390 614.900 1206.770 614.910 ;
        RECT 1424.685 614.530 1425.015 614.545 ;
        RECT 1441.910 614.530 1442.290 614.540 ;
        RECT 1424.685 614.230 1442.290 614.530 ;
        RECT 1510.950 614.530 1511.250 615.590 ;
        RECT 1690.105 615.590 1704.450 615.890 ;
        RECT 1690.105 615.575 1690.435 615.590 ;
        RECT 1606.385 615.210 1606.715 615.225 ;
        RECT 1559.710 614.910 1606.715 615.210 ;
        RECT 1559.710 614.530 1560.010 614.910 ;
        RECT 1606.385 614.895 1606.715 614.910 ;
        RECT 1642.265 614.530 1642.595 614.545 ;
        RECT 1510.950 614.230 1560.010 614.530 ;
        RECT 1641.590 614.230 1642.595 614.530 ;
        RECT 1704.150 614.530 1704.450 615.590 ;
        RECT 1849.510 615.590 1911.490 615.890 ;
        RECT 1799.125 615.210 1799.455 615.225 ;
        RECT 1752.910 614.910 1799.455 615.210 ;
        RECT 1752.910 614.530 1753.210 614.910 ;
        RECT 1799.125 614.895 1799.455 614.910 ;
        RECT 1801.885 615.210 1802.215 615.225 ;
        RECT 1801.885 614.910 1835.090 615.210 ;
        RECT 1801.885 614.895 1802.215 614.910 ;
        RECT 1704.150 614.230 1753.210 614.530 ;
        RECT 1834.790 614.530 1835.090 614.910 ;
        RECT 1849.510 614.530 1849.810 615.590 ;
        RECT 1911.110 615.580 1911.490 615.590 ;
        RECT 2117.905 615.890 2118.235 615.905 ;
        RECT 2235.910 615.890 2236.210 616.270 ;
        RECT 2269.910 615.890 2270.290 615.900 ;
        RECT 2117.905 615.590 2163.530 615.890 ;
        RECT 2235.910 615.590 2270.290 615.890 ;
        RECT 2117.905 615.575 2118.235 615.590 ;
        RECT 1834.790 614.230 1849.810 614.530 ;
        RECT 1911.110 614.530 1911.490 614.540 ;
        RECT 1959.665 614.530 1959.995 614.545 ;
        RECT 1911.110 614.230 1959.995 614.530 ;
        RECT 1424.685 614.215 1425.015 614.230 ;
        RECT 1441.910 614.220 1442.290 614.230 ;
        RECT 1606.385 613.170 1606.715 613.185 ;
        RECT 1641.590 613.170 1641.890 614.230 ;
        RECT 1642.265 614.215 1642.595 614.230 ;
        RECT 1911.110 614.220 1911.490 614.230 ;
        RECT 1959.665 614.215 1959.995 614.230 ;
        RECT 2055.805 614.530 2056.135 614.545 ;
        RECT 2070.065 614.530 2070.395 614.545 ;
        RECT 2055.805 614.230 2070.395 614.530 ;
        RECT 2163.230 614.530 2163.530 615.590 ;
        RECT 2269.910 615.580 2270.290 615.590 ;
        RECT 2294.085 615.890 2294.415 615.905 ;
        RECT 2504.305 615.890 2504.635 615.905 ;
        RECT 2697.505 615.890 2697.835 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2294.085 615.590 2353.050 615.890 ;
        RECT 2294.085 615.575 2294.415 615.590 ;
        RECT 2352.750 615.210 2353.050 615.590 ;
        RECT 2401.510 615.590 2429.410 615.890 ;
        RECT 2352.750 614.910 2400.890 615.210 ;
        RECT 2173.310 614.530 2173.690 614.540 ;
        RECT 2163.230 614.230 2173.690 614.530 ;
        RECT 2400.590 614.530 2400.890 614.910 ;
        RECT 2401.510 614.530 2401.810 615.590 ;
        RECT 2429.110 615.210 2429.410 615.590 ;
        RECT 2504.305 615.590 2526.010 615.890 ;
        RECT 2504.305 615.575 2504.635 615.590 ;
        RECT 2456.465 615.210 2456.795 615.225 ;
        RECT 2429.110 614.910 2456.795 615.210 ;
        RECT 2456.465 614.895 2456.795 614.910 ;
        RECT 2400.590 614.230 2401.810 614.530 ;
        RECT 2525.710 614.530 2526.010 615.590 ;
        RECT 2697.505 615.590 2739.450 615.890 ;
        RECT 2697.505 615.575 2697.835 615.590 ;
        RECT 2574.225 615.210 2574.555 615.225 ;
        RECT 2621.605 615.210 2621.935 615.225 ;
        RECT 2574.225 614.910 2621.935 615.210 ;
        RECT 2739.150 615.210 2739.450 615.590 ;
        RECT 2787.910 615.590 2836.050 615.890 ;
        RECT 2739.150 614.910 2787.290 615.210 ;
        RECT 2574.225 614.895 2574.555 614.910 ;
        RECT 2621.605 614.895 2621.935 614.910 ;
        RECT 2573.305 614.530 2573.635 614.545 ;
        RECT 2525.710 614.230 2573.635 614.530 ;
        RECT 2055.805 614.215 2056.135 614.230 ;
        RECT 2070.065 614.215 2070.395 614.230 ;
        RECT 2173.310 614.220 2173.690 614.230 ;
        RECT 2573.305 614.215 2573.635 614.230 ;
        RECT 2622.525 614.530 2622.855 614.545 ;
        RECT 2649.665 614.530 2649.995 614.545 ;
        RECT 2622.525 614.230 2649.995 614.530 ;
        RECT 2786.990 614.530 2787.290 614.910 ;
        RECT 2787.910 614.530 2788.210 615.590 ;
        RECT 2835.750 615.210 2836.050 615.590 ;
        RECT 2916.710 615.590 2924.800 615.890 ;
        RECT 2916.710 615.210 2917.010 615.590 ;
        RECT 2835.750 614.910 2883.890 615.210 ;
        RECT 2786.990 614.230 2788.210 614.530 ;
        RECT 2883.590 614.530 2883.890 614.910 ;
        RECT 2884.510 614.910 2917.010 615.210 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
        RECT 2884.510 614.530 2884.810 614.910 ;
        RECT 2883.590 614.230 2884.810 614.530 ;
        RECT 2622.525 614.215 2622.855 614.230 ;
        RECT 2649.665 614.215 2649.995 614.230 ;
        RECT 2007.505 613.850 2007.835 613.865 ;
        RECT 2007.100 613.550 2008.050 613.850 ;
        RECT 2007.505 613.535 2008.050 613.550 ;
        RECT 1606.385 612.870 1641.890 613.170 ;
        RECT 2007.750 613.170 2008.050 613.535 ;
        RECT 2021.305 613.170 2021.635 613.185 ;
        RECT 2007.750 612.870 2021.635 613.170 ;
        RECT 1606.385 612.855 1606.715 612.870 ;
        RECT 2021.305 612.855 2021.635 612.870 ;
      LAYER via3 ;
        RECT 1206.420 2497.820 1206.740 2498.140 ;
        RECT 2269.940 616.940 2270.260 617.260 ;
        RECT 1206.420 614.900 1206.740 615.220 ;
        RECT 2173.340 616.260 2173.660 616.580 ;
        RECT 1441.940 615.580 1442.260 615.900 ;
        RECT 1441.940 614.220 1442.260 614.540 ;
        RECT 1911.140 615.580 1911.460 615.900 ;
        RECT 1911.140 614.220 1911.460 614.540 ;
        RECT 2269.940 615.580 2270.260 615.900 ;
        RECT 2173.340 614.220 2173.660 614.540 ;
      LAYER met4 ;
        RECT 1206.415 2497.815 1206.745 2498.145 ;
        RECT 1206.430 615.225 1206.730 2497.815 ;
        RECT 2269.935 616.935 2270.265 617.265 ;
        RECT 2173.335 616.255 2173.665 616.585 ;
        RECT 1441.935 615.575 1442.265 615.905 ;
        RECT 1911.135 615.575 1911.465 615.905 ;
        RECT 1206.415 614.895 1206.745 615.225 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1441.950 614.545 1442.250 615.575 ;
        RECT 1911.150 614.545 1911.450 615.575 ;
        RECT 2173.350 614.545 2173.650 616.255 ;
        RECT 2269.950 615.905 2270.250 616.935 ;
        RECT 2269.935 615.575 2270.265 615.905 ;
        RECT 1441.935 614.215 1442.265 614.545 ;
        RECT 1911.135 614.215 1911.465 614.545 ;
        RECT 2173.335 614.215 2173.665 614.545 ;
>>>>>>> re-updated local openlane
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 86.090 2512.500 86.410 2512.560 ;
        RECT 1746.690 2512.500 1747.010 2512.560 ;
        RECT 86.090 2512.360 1747.010 2512.500 ;
        RECT 86.090 2512.300 86.410 2512.360 ;
        RECT 1746.690 2512.300 1747.010 2512.360 ;
        RECT 15.250 1621.360 15.570 1621.420 ;
        RECT 86.090 1621.360 86.410 1621.420 ;
        RECT 15.250 1621.220 86.410 1621.360 ;
        RECT 15.250 1621.160 15.570 1621.220 ;
        RECT 86.090 1621.160 86.410 1621.220 ;
      LAYER via ;
        RECT 86.120 2512.300 86.380 2512.560 ;
        RECT 1746.720 2512.300 1746.980 2512.560 ;
        RECT 15.280 1621.160 15.540 1621.420 ;
        RECT 86.120 1621.160 86.380 1621.420 ;
      LAYER met2 ;
        RECT 86.120 2512.270 86.380 2512.590 ;
        RECT 1746.720 2512.270 1746.980 2512.590 ;
        RECT 86.180 1621.450 86.320 2512.270 ;
        RECT 1746.780 2500.000 1746.920 2512.270 ;
        RECT 1746.710 2496.000 1746.990 2500.000 ;
        RECT 15.280 1621.130 15.540 1621.450 ;
        RECT 86.120 1621.130 86.380 1621.450 ;
        RECT 15.340 1615.525 15.480 1621.130 ;
        RECT 15.270 1615.155 15.550 1615.525 ;
      LAYER via2 ;
        RECT 15.270 1615.200 15.550 1615.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1614.740 0.300 1615.940 ;
=======
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 15.245 1615.490 15.575 1615.505 ;
        RECT -4.800 1615.190 15.575 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
<<<<<<< HEAD
        RECT 13.865 1615.175 14.195 1615.190 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 15.245 1615.175 15.575 1615.190 ;
>>>>>>> re-updated local openlane
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 121.050 2513.520 121.370 2513.580 ;
        RECT 1766.010 2513.520 1766.330 2513.580 ;
        RECT 121.050 2513.380 1766.330 2513.520 ;
        RECT 121.050 2513.320 121.370 2513.380 ;
        RECT 1766.010 2513.320 1766.330 2513.380 ;
        RECT 16.630 1400.700 16.950 1400.760 ;
        RECT 121.050 1400.700 121.370 1400.760 ;
        RECT 16.630 1400.560 121.370 1400.700 ;
        RECT 16.630 1400.500 16.950 1400.560 ;
        RECT 121.050 1400.500 121.370 1400.560 ;
      LAYER via ;
        RECT 121.080 2513.320 121.340 2513.580 ;
        RECT 1766.040 2513.320 1766.300 2513.580 ;
        RECT 16.660 1400.500 16.920 1400.760 ;
        RECT 121.080 1400.500 121.340 1400.760 ;
      LAYER met2 ;
        RECT 121.080 2513.290 121.340 2513.610 ;
        RECT 1766.040 2513.290 1766.300 2513.610 ;
        RECT 121.140 1400.790 121.280 2513.290 ;
        RECT 1766.100 2500.000 1766.240 2513.290 ;
        RECT 1766.030 2496.000 1766.310 2500.000 ;
        RECT 16.660 1400.645 16.920 1400.790 ;
        RECT 16.650 1400.275 16.930 1400.645 ;
        RECT 121.080 1400.470 121.340 1400.790 ;
      LAYER via2 ;
        RECT 16.650 1400.320 16.930 1400.600 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1399.860 0.300 1401.060 ;
=======
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 16.625 1400.610 16.955 1400.625 ;
        RECT -4.800 1400.310 16.955 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
<<<<<<< HEAD
        RECT 13.865 1400.295 14.195 1400.310 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 1400.295 16.955 1400.310 ;
>>>>>>> re-updated local openlane
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1784.025 2491.605 1784.195 2496.875 ;
      LAYER mcon ;
        RECT 1784.025 2496.705 1784.195 2496.875 ;
      LAYER met1 ;
        RECT 1783.950 2496.860 1784.270 2496.920 ;
        RECT 1783.755 2496.720 1784.270 2496.860 ;
        RECT 1783.950 2496.660 1784.270 2496.720 ;
        RECT 18.010 2491.760 18.330 2491.820 ;
        RECT 1783.965 2491.760 1784.255 2491.805 ;
        RECT 18.010 2491.620 1784.255 2491.760 ;
        RECT 18.010 2491.560 18.330 2491.620 ;
        RECT 1783.965 2491.575 1784.255 2491.620 ;
      LAYER via ;
        RECT 1783.980 2496.660 1784.240 2496.920 ;
        RECT 18.040 2491.560 18.300 2491.820 ;
      LAYER met2 ;
        RECT 1783.980 2496.690 1784.240 2496.950 ;
        RECT 1785.350 2496.690 1785.630 2500.000 ;
        RECT 1783.980 2496.630 1785.630 2496.690 ;
        RECT 1784.040 2496.550 1785.630 2496.630 ;
        RECT 1785.350 2496.000 1785.630 2496.550 ;
        RECT 18.040 2491.530 18.300 2491.850 ;
        RECT 18.100 1185.085 18.240 2491.530 ;
        RECT 18.030 1184.715 18.310 1185.085 ;
      LAYER via2 ;
        RECT 18.030 1184.760 18.310 1185.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 1184.300 0.300 1185.500 ;
=======
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 18.005 1185.050 18.335 1185.065 ;
        RECT -4.800 1184.750 18.335 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
<<<<<<< HEAD
        RECT 13.865 1184.735 14.195 1184.750 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 18.005 1184.735 18.335 1184.750 ;
>>>>>>> re-updated local openlane
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 155.550 2513.180 155.870 2513.240 ;
        RECT 1804.650 2513.180 1804.970 2513.240 ;
        RECT 155.550 2513.040 1804.970 2513.180 ;
        RECT 155.550 2512.980 155.870 2513.040 ;
        RECT 1804.650 2512.980 1804.970 2513.040 ;
        RECT 16.630 972.640 16.950 972.700 ;
        RECT 155.550 972.640 155.870 972.700 ;
        RECT 16.630 972.500 155.870 972.640 ;
        RECT 16.630 972.440 16.950 972.500 ;
        RECT 155.550 972.440 155.870 972.500 ;
      LAYER via ;
        RECT 155.580 2512.980 155.840 2513.240 ;
        RECT 1804.680 2512.980 1804.940 2513.240 ;
        RECT 16.660 972.440 16.920 972.700 ;
        RECT 155.580 972.440 155.840 972.700 ;
      LAYER met2 ;
        RECT 155.580 2512.950 155.840 2513.270 ;
        RECT 1804.680 2512.950 1804.940 2513.270 ;
        RECT 155.640 972.730 155.780 2512.950 ;
        RECT 1804.740 2500.000 1804.880 2512.950 ;
        RECT 1804.670 2496.000 1804.950 2500.000 ;
        RECT 16.660 972.410 16.920 972.730 ;
        RECT 155.580 972.410 155.840 972.730 ;
        RECT 16.720 969.525 16.860 972.410 ;
        RECT 16.650 969.155 16.930 969.525 ;
      LAYER via2 ;
        RECT 16.650 969.200 16.930 969.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 968.740 0.300 969.940 ;
=======
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 16.625 969.490 16.955 969.505 ;
        RECT -4.800 969.190 16.955 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
<<<<<<< HEAD
        RECT 16.165 969.175 16.495 969.190 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.625 969.175 16.955 969.190 ;
>>>>>>> re-updated local openlane
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1822.665 2491.265 1822.835 2496.535 ;
      LAYER mcon ;
        RECT 1822.665 2496.365 1822.835 2496.535 ;
      LAYER met1 ;
        RECT 1822.590 2496.520 1822.910 2496.580 ;
        RECT 1822.395 2496.380 1822.910 2496.520 ;
        RECT 1822.590 2496.320 1822.910 2496.380 ;
        RECT 17.550 2491.420 17.870 2491.480 ;
        RECT 1822.605 2491.420 1822.895 2491.465 ;
        RECT 17.550 2491.280 1822.895 2491.420 ;
        RECT 17.550 2491.220 17.870 2491.280 ;
        RECT 1822.605 2491.235 1822.895 2491.280 ;
      LAYER via ;
        RECT 1822.620 2496.320 1822.880 2496.580 ;
        RECT 17.580 2491.220 17.840 2491.480 ;
      LAYER met2 ;
        RECT 1823.990 2496.690 1824.270 2500.000 ;
        RECT 1822.680 2496.610 1824.270 2496.690 ;
        RECT 1822.620 2496.550 1824.270 2496.610 ;
        RECT 1822.620 2496.290 1822.880 2496.550 ;
        RECT 1823.990 2496.000 1824.270 2496.550 ;
        RECT 17.580 2491.190 17.840 2491.510 ;
        RECT 17.640 753.965 17.780 2491.190 ;
        RECT 17.570 753.595 17.850 753.965 ;
      LAYER via2 ;
        RECT 17.570 753.640 17.850 753.920 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 753.180 0.300 754.380 ;
=======
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 17.545 753.930 17.875 753.945 ;
        RECT -4.800 753.630 17.875 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
<<<<<<< HEAD
        RECT 13.865 753.615 14.195 753.630 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 17.545 753.615 17.875 753.630 ;
>>>>>>> re-updated local openlane
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.990 2511.820 162.310 2511.880 ;
        RECT 1843.290 2511.820 1843.610 2511.880 ;
        RECT 161.990 2511.680 1843.610 2511.820 ;
        RECT 161.990 2511.620 162.310 2511.680 ;
        RECT 1843.290 2511.620 1843.610 2511.680 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 161.990 544.920 162.310 544.980 ;
        RECT 16.170 544.780 162.310 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 161.990 544.720 162.310 544.780 ;
      LAYER via ;
        RECT 162.020 2511.620 162.280 2511.880 ;
        RECT 1843.320 2511.620 1843.580 2511.880 ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 162.020 544.720 162.280 544.980 ;
      LAYER met2 ;
        RECT 162.020 2511.590 162.280 2511.910 ;
        RECT 1843.320 2511.590 1843.580 2511.910 ;
        RECT 162.080 545.010 162.220 2511.590 ;
        RECT 1843.380 2500.000 1843.520 2511.590 ;
        RECT 1843.310 2496.000 1843.590 2500.000 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 162.020 544.690 162.280 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 537.620 0.300 538.820 ;
=======
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
<<<<<<< HEAD
        RECT 17.545 538.055 17.875 538.070 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 16.165 538.055 16.495 538.070 ;
>>>>>>> re-updated local openlane
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1861.305 2490.925 1861.475 2496.535 ;
      LAYER mcon ;
        RECT 1861.305 2496.365 1861.475 2496.535 ;
      LAYER met1 ;
        RECT 1861.230 2496.520 1861.550 2496.580 ;
        RECT 1861.035 2496.380 1861.550 2496.520 ;
        RECT 1861.230 2496.320 1861.550 2496.380 ;
        RECT 17.090 2491.080 17.410 2491.140 ;
        RECT 1861.245 2491.080 1861.535 2491.125 ;
        RECT 17.090 2490.940 1861.535 2491.080 ;
        RECT 17.090 2490.880 17.410 2490.940 ;
        RECT 1861.245 2490.895 1861.535 2490.940 ;
      LAYER via ;
        RECT 1861.260 2496.320 1861.520 2496.580 ;
        RECT 17.120 2490.880 17.380 2491.140 ;
      LAYER met2 ;
        RECT 1862.630 2496.690 1862.910 2500.000 ;
        RECT 1861.320 2496.610 1862.910 2496.690 ;
        RECT 1861.260 2496.550 1862.910 2496.610 ;
        RECT 1861.260 2496.290 1861.520 2496.550 ;
        RECT 1862.630 2496.000 1862.910 2496.550 ;
        RECT 17.120 2490.850 17.380 2491.170 ;
        RECT 17.180 322.845 17.320 2490.850 ;
        RECT 17.110 322.475 17.390 322.845 ;
      LAYER via2 ;
        RECT 17.110 322.520 17.390 322.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 322.060 0.300 323.260 ;
=======
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 17.085 322.810 17.415 322.825 ;
        RECT -4.800 322.510 17.415 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
<<<<<<< HEAD
        RECT 15.705 322.495 16.035 322.510 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 17.085 322.495 17.415 322.510 ;
>>>>>>> re-updated local openlane
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 168.890 110.400 169.210 110.460 ;
        RECT 15.710 110.260 169.210 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 168.890 110.200 169.210 110.260 ;
      LAYER via ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 168.920 110.200 169.180 110.460 ;
      LAYER met2 ;
        RECT 168.910 2512.755 169.190 2513.125 ;
        RECT 1881.950 2512.755 1882.230 2513.125 ;
        RECT 168.980 110.490 169.120 2512.755 ;
        RECT 1882.020 2500.000 1882.160 2512.755 ;
        RECT 1881.950 2496.000 1882.230 2500.000 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 168.920 110.170 169.180 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 168.910 2512.800 169.190 2513.080 ;
        RECT 1881.950 2512.800 1882.230 2513.080 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT -4.800 106.500 0.300 107.700 ;
=======
=======
        RECT 168.885 2513.090 169.215 2513.105 ;
        RECT 1881.925 2513.090 1882.255 2513.105 ;
        RECT 168.885 2512.790 1882.255 2513.090 ;
        RECT 168.885 2512.775 169.215 2512.790 ;
        RECT 1881.925 2512.775 1882.255 2512.790 ;
>>>>>>> re-updated local openlane
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
<<<<<<< HEAD
        RECT 14.785 106.935 15.115 106.950 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 15.705 106.935 16.035 106.950 ;
>>>>>>> re-updated local openlane
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1448.610 849.900 1448.930 849.960 ;
        RECT 1490.010 849.900 1490.330 849.960 ;
        RECT 1448.610 849.760 1490.330 849.900 ;
        RECT 1448.610 849.700 1448.930 849.760 ;
        RECT 1490.010 849.700 1490.330 849.760 ;
        RECT 1932.070 849.900 1932.390 849.960 ;
        RECT 1956.450 849.900 1956.770 849.960 ;
        RECT 1932.070 849.760 1956.770 849.900 ;
        RECT 1932.070 849.700 1932.390 849.760 ;
        RECT 1956.450 849.700 1956.770 849.760 ;
        RECT 2476.710 849.900 2477.030 849.960 ;
        RECT 2511.210 849.900 2511.530 849.960 ;
        RECT 2476.710 849.760 2511.530 849.900 ;
        RECT 2476.710 849.700 2477.030 849.760 ;
        RECT 2511.210 849.700 2511.530 849.760 ;
        RECT 1799.130 849.560 1799.450 849.620 ;
        RECT 1801.890 849.560 1802.210 849.620 ;
        RECT 1799.130 849.420 1802.210 849.560 ;
        RECT 1799.130 849.360 1799.450 849.420 ;
        RECT 1801.890 849.360 1802.210 849.420 ;
        RECT 1642.270 849.220 1642.590 849.280 ;
        RECT 1690.110 849.220 1690.430 849.280 ;
        RECT 1642.270 849.080 1690.430 849.220 ;
        RECT 1642.270 849.020 1642.590 849.080 ;
        RECT 1690.110 849.020 1690.430 849.080 ;
        RECT 2621.610 849.220 2621.930 849.280 ;
        RECT 2625.290 849.220 2625.610 849.280 ;
        RECT 2621.610 849.080 2625.610 849.220 ;
        RECT 2621.610 849.020 2621.930 849.080 ;
        RECT 2625.290 849.020 2625.610 849.080 ;
        RECT 2649.670 849.220 2649.990 849.280 ;
        RECT 2697.510 849.220 2697.830 849.280 ;
        RECT 2649.670 849.080 2697.830 849.220 ;
        RECT 2649.670 849.020 2649.990 849.080 ;
        RECT 2697.510 849.020 2697.830 849.080 ;
      LAYER via ;
        RECT 1448.640 849.700 1448.900 849.960 ;
        RECT 1490.040 849.700 1490.300 849.960 ;
        RECT 1932.100 849.700 1932.360 849.960 ;
        RECT 1956.480 849.700 1956.740 849.960 ;
        RECT 2476.740 849.700 2477.000 849.960 ;
        RECT 2511.240 849.700 2511.500 849.960 ;
        RECT 1799.160 849.360 1799.420 849.620 ;
        RECT 1801.920 849.360 1802.180 849.620 ;
        RECT 1642.300 849.020 1642.560 849.280 ;
        RECT 1690.140 849.020 1690.400 849.280 ;
        RECT 2621.640 849.020 2621.900 849.280 ;
        RECT 2625.320 849.020 2625.580 849.280 ;
        RECT 2649.700 849.020 2649.960 849.280 ;
        RECT 2697.540 849.020 2697.800 849.280 ;
      LAYER met2 ;
        RECT 1224.150 2498.050 1224.430 2500.000 ;
        RECT 1225.990 2498.050 1226.270 2498.165 ;
        RECT 1224.150 2497.910 1226.270 2498.050 ;
        RECT 1224.150 2496.000 1224.430 2497.910 ;
        RECT 1225.990 2497.795 1226.270 2497.910 ;
        RECT 1994.650 851.090 1994.930 851.205 ;
        RECT 1993.800 850.950 1994.930 851.090 ;
        RECT 1993.800 850.525 1993.940 850.950 ;
        RECT 1994.650 850.835 1994.930 850.950 ;
        RECT 2187.390 850.835 2187.670 851.205 ;
        RECT 1393.890 850.155 1394.170 850.525 ;
        RECT 1490.030 850.155 1490.310 850.525 ;
        RECT 1690.130 850.155 1690.410 850.525 ;
        RECT 1956.470 850.155 1956.750 850.525 ;
        RECT 1993.730 850.155 1994.010 850.525 ;
        RECT 2090.790 850.410 2091.070 850.525 ;
        RECT 2090.400 850.270 2091.070 850.410 ;
        RECT 1393.960 849.845 1394.100 850.155 ;
        RECT 1490.100 849.990 1490.240 850.155 ;
        RECT 1448.640 849.845 1448.900 849.990 ;
        RECT 1393.890 849.475 1394.170 849.845 ;
        RECT 1448.630 849.475 1448.910 849.845 ;
        RECT 1490.040 849.670 1490.300 849.990 ;
        RECT 1606.410 849.475 1606.690 849.845 ;
        RECT 1606.480 847.805 1606.620 849.475 ;
        RECT 1690.200 849.310 1690.340 850.155 ;
        RECT 1956.540 849.990 1956.680 850.155 ;
        RECT 1932.100 849.845 1932.360 849.990 ;
        RECT 1799.150 849.475 1799.430 849.845 ;
        RECT 1801.910 849.475 1802.190 849.845 ;
        RECT 1932.090 849.475 1932.370 849.845 ;
        RECT 1956.480 849.670 1956.740 849.990 ;
        RECT 2090.400 849.845 2090.540 850.270 ;
        RECT 2090.790 850.155 2091.070 850.270 ;
        RECT 2090.330 849.475 2090.610 849.845 ;
        RECT 1799.160 849.330 1799.420 849.475 ;
        RECT 1801.920 849.330 1802.180 849.475 ;
        RECT 1642.300 849.165 1642.560 849.310 ;
        RECT 1642.290 848.795 1642.570 849.165 ;
        RECT 1690.140 848.990 1690.400 849.310 ;
        RECT 2186.930 849.050 2187.210 849.165 ;
        RECT 2187.460 849.050 2187.600 850.835 ;
        RECT 2283.070 850.410 2283.350 850.525 ;
        RECT 2283.990 850.410 2284.270 850.525 ;
        RECT 2283.070 850.270 2284.270 850.410 ;
        RECT 2283.070 850.155 2283.350 850.270 ;
        RECT 2283.990 850.155 2284.270 850.270 ;
        RECT 2511.230 850.155 2511.510 850.525 ;
        RECT 2697.530 850.155 2697.810 850.525 ;
        RECT 2511.300 849.990 2511.440 850.155 ;
        RECT 2476.740 849.845 2477.000 849.990 ;
        RECT 2476.730 849.475 2477.010 849.845 ;
        RECT 2511.240 849.670 2511.500 849.990 ;
        RECT 2697.600 849.310 2697.740 850.155 ;
        RECT 2621.640 849.165 2621.900 849.310 ;
        RECT 2625.320 849.165 2625.580 849.310 ;
        RECT 2649.700 849.165 2649.960 849.310 ;
        RECT 2186.930 848.910 2187.600 849.050 ;
        RECT 2186.930 848.795 2187.210 848.910 ;
        RECT 2621.630 848.795 2621.910 849.165 ;
        RECT 2625.310 848.795 2625.590 849.165 ;
        RECT 2649.690 848.795 2649.970 849.165 ;
        RECT 2697.540 848.990 2697.800 849.310 ;
        RECT 1606.410 847.435 1606.690 847.805 ;
      LAYER via2 ;
        RECT 1225.990 2497.840 1226.270 2498.120 ;
        RECT 1994.650 850.880 1994.930 851.160 ;
        RECT 2187.390 850.880 2187.670 851.160 ;
        RECT 1393.890 850.200 1394.170 850.480 ;
        RECT 1490.030 850.200 1490.310 850.480 ;
        RECT 1690.130 850.200 1690.410 850.480 ;
        RECT 1956.470 850.200 1956.750 850.480 ;
        RECT 1993.730 850.200 1994.010 850.480 ;
        RECT 1393.890 849.520 1394.170 849.800 ;
        RECT 1448.630 849.520 1448.910 849.800 ;
        RECT 1606.410 849.520 1606.690 849.800 ;
        RECT 1799.150 849.520 1799.430 849.800 ;
        RECT 1801.910 849.520 1802.190 849.800 ;
        RECT 1932.090 849.520 1932.370 849.800 ;
        RECT 2090.790 850.200 2091.070 850.480 ;
        RECT 2090.330 849.520 2090.610 849.800 ;
        RECT 1642.290 848.840 1642.570 849.120 ;
        RECT 2186.930 848.840 2187.210 849.120 ;
        RECT 2283.070 850.200 2283.350 850.480 ;
        RECT 2283.990 850.200 2284.270 850.480 ;
        RECT 2511.230 850.200 2511.510 850.480 ;
        RECT 2697.530 850.200 2697.810 850.480 ;
        RECT 2476.730 849.520 2477.010 849.800 ;
        RECT 2621.630 848.840 2621.910 849.120 ;
        RECT 2625.310 848.840 2625.590 849.120 ;
        RECT 2649.690 848.840 2649.970 849.120 ;
        RECT 1606.410 847.480 1606.690 847.760 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 849.740 2924.800 850.940 ;
=======
        RECT 1226.425 2498.140 1226.755 2498.145 ;
        RECT 1226.425 2498.130 1227.010 2498.140 ;
        RECT 1226.425 2497.830 1227.210 2498.130 ;
        RECT 1226.425 2497.820 1227.010 2497.830 ;
        RECT 1226.425 2497.815 1226.755 2497.820 ;
        RECT 1226.630 860.010 1227.010 860.020 ;
        RECT 1255.405 860.010 1255.735 860.025 ;
        RECT 1226.630 859.710 1255.735 860.010 ;
        RECT 1226.630 859.700 1227.010 859.710 ;
        RECT 1255.405 859.695 1255.735 859.710 ;
        RECT 1980.110 851.850 1980.490 851.860 ;
        RECT 2028.205 851.850 2028.535 851.865 ;
        RECT 1980.110 851.550 2028.535 851.850 ;
        RECT 1980.110 851.540 1980.490 851.550 ;
        RECT 2028.205 851.535 2028.535 851.550 ;
        RECT 1325.325 851.170 1325.655 851.185 ;
=======
        RECT 1225.965 2498.130 1226.295 2498.145 ;
        RECT 1226.630 2498.130 1227.010 2498.140 ;
        RECT 1225.965 2497.830 1227.010 2498.130 ;
        RECT 1225.965 2497.815 1226.295 2497.830 ;
        RECT 1226.630 2497.820 1227.010 2497.830 ;
>>>>>>> re-updated local openlane
        RECT 1345.310 851.170 1345.690 851.180 ;
        RECT 1994.625 851.170 1994.955 851.185 ;
        RECT 2187.365 851.170 2187.695 851.185 ;
        RECT 1269.910 850.870 1318.970 851.170 ;
        RECT 1226.630 850.490 1227.010 850.500 ;
        RECT 1269.910 850.490 1270.210 850.870 ;
        RECT 1226.630 850.190 1270.210 850.490 ;
        RECT 1226.630 850.180 1227.010 850.190 ;
        RECT 1318.670 849.810 1318.970 850.870 ;
        RECT 1345.310 850.870 1370.490 851.170 ;
        RECT 1345.310 850.860 1345.690 850.870 ;
        RECT 1370.190 850.490 1370.490 850.870 ;
        RECT 1994.625 850.870 2043.010 851.170 ;
        RECT 1994.625 850.855 1994.955 850.870 ;
        RECT 1393.865 850.490 1394.195 850.505 ;
        RECT 1370.190 850.190 1394.195 850.490 ;
        RECT 1393.865 850.175 1394.195 850.190 ;
        RECT 1490.005 850.490 1490.335 850.505 ;
        RECT 1690.105 850.490 1690.435 850.505 ;
        RECT 1883.510 850.490 1883.890 850.500 ;
        RECT 1490.005 850.190 1511.250 850.490 ;
        RECT 1490.005 850.175 1490.335 850.190 ;
        RECT 1345.310 849.810 1345.690 849.820 ;
        RECT 1318.670 849.510 1345.690 849.810 ;
        RECT 1345.310 849.500 1345.690 849.510 ;
        RECT 1393.865 849.810 1394.195 849.825 ;
        RECT 1448.605 849.810 1448.935 849.825 ;
        RECT 1393.865 849.510 1448.935 849.810 ;
        RECT 1393.865 849.495 1394.195 849.510 ;
        RECT 1448.605 849.495 1448.935 849.510 ;
        RECT 1510.950 849.130 1511.250 850.190 ;
        RECT 1690.105 850.190 1704.450 850.490 ;
        RECT 1690.105 850.175 1690.435 850.190 ;
        RECT 1606.385 849.810 1606.715 849.825 ;
        RECT 1559.710 849.510 1606.715 849.810 ;
        RECT 1559.710 849.130 1560.010 849.510 ;
        RECT 1606.385 849.495 1606.715 849.510 ;
        RECT 1642.265 849.130 1642.595 849.145 ;
        RECT 1510.950 848.830 1560.010 849.130 ;
        RECT 1641.590 848.830 1642.595 849.130 ;
        RECT 1704.150 849.130 1704.450 850.190 ;
        RECT 1849.510 850.190 1883.890 850.490 ;
        RECT 1799.125 849.810 1799.455 849.825 ;
        RECT 1752.910 849.510 1799.455 849.810 ;
        RECT 1752.910 849.130 1753.210 849.510 ;
        RECT 1799.125 849.495 1799.455 849.510 ;
        RECT 1801.885 849.810 1802.215 849.825 ;
        RECT 1801.885 849.510 1835.090 849.810 ;
        RECT 1801.885 849.495 1802.215 849.510 ;
        RECT 1704.150 848.830 1753.210 849.130 ;
        RECT 1834.790 849.130 1835.090 849.510 ;
        RECT 1849.510 849.130 1849.810 850.190 ;
        RECT 1883.510 850.180 1883.890 850.190 ;
        RECT 1956.445 850.490 1956.775 850.505 ;
        RECT 1993.705 850.490 1994.035 850.505 ;
        RECT 1956.445 850.190 1994.035 850.490 ;
        RECT 2042.710 850.490 2043.010 850.870 ;
        RECT 2187.365 850.870 2236.210 851.170 ;
        RECT 2187.365 850.855 2187.695 850.870 ;
        RECT 2090.765 850.490 2091.095 850.505 ;
        RECT 2235.910 850.490 2236.210 850.870 ;
        RECT 2283.045 850.490 2283.375 850.505 ;
        RECT 2042.710 850.190 2077.050 850.490 ;
        RECT 1956.445 850.175 1956.775 850.190 ;
        RECT 1993.705 850.175 1994.035 850.190 ;
        RECT 1932.065 849.810 1932.395 849.825 ;
        RECT 1834.790 848.830 1849.810 849.130 ;
        RECT 1931.390 849.510 1932.395 849.810 ;
        RECT 2076.750 849.810 2077.050 850.190 ;
        RECT 2090.765 850.190 2163.530 850.490 ;
        RECT 2235.910 850.190 2283.375 850.490 ;
        RECT 2090.765 850.175 2091.095 850.190 ;
        RECT 2090.305 849.810 2090.635 849.825 ;
        RECT 2076.750 849.510 2090.635 849.810 ;
        RECT 1606.385 847.770 1606.715 847.785 ;
        RECT 1641.590 847.770 1641.890 848.830 ;
        RECT 1642.265 848.815 1642.595 848.830 ;
        RECT 1883.510 848.450 1883.890 848.460 ;
        RECT 1931.390 848.450 1931.690 849.510 ;
        RECT 1932.065 849.495 1932.395 849.510 ;
        RECT 2090.305 849.495 2090.635 849.510 ;
        RECT 2163.230 849.130 2163.530 850.190 ;
        RECT 2283.045 850.175 2283.375 850.190 ;
        RECT 2283.965 850.490 2284.295 850.505 ;
        RECT 2511.205 850.490 2511.535 850.505 ;
        RECT 2697.505 850.490 2697.835 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2283.965 850.190 2353.050 850.490 ;
        RECT 2283.965 850.175 2284.295 850.190 ;
        RECT 2352.750 849.810 2353.050 850.190 ;
        RECT 2401.510 850.190 2429.410 850.490 ;
        RECT 2352.750 849.510 2400.890 849.810 ;
        RECT 2186.905 849.130 2187.235 849.145 ;
        RECT 2163.230 848.830 2187.235 849.130 ;
        RECT 2400.590 849.130 2400.890 849.510 ;
        RECT 2401.510 849.130 2401.810 850.190 ;
        RECT 2429.110 849.810 2429.410 850.190 ;
        RECT 2511.205 850.190 2526.010 850.490 ;
        RECT 2511.205 850.175 2511.535 850.190 ;
        RECT 2476.705 849.810 2477.035 849.825 ;
        RECT 2429.110 849.510 2477.035 849.810 ;
        RECT 2476.705 849.495 2477.035 849.510 ;
        RECT 2400.590 848.830 2401.810 849.130 ;
        RECT 2525.710 849.130 2526.010 850.190 ;
        RECT 2697.505 850.190 2739.450 850.490 ;
        RECT 2697.505 850.175 2697.835 850.190 ;
        RECT 2739.150 849.810 2739.450 850.190 ;
        RECT 2787.910 850.190 2836.050 850.490 ;
        RECT 2739.150 849.510 2787.290 849.810 ;
        RECT 2621.605 849.130 2621.935 849.145 ;
        RECT 2525.710 848.830 2621.935 849.130 ;
        RECT 2186.905 848.815 2187.235 848.830 ;
        RECT 2621.605 848.815 2621.935 848.830 ;
        RECT 2625.285 849.130 2625.615 849.145 ;
        RECT 2649.665 849.130 2649.995 849.145 ;
        RECT 2625.285 848.830 2649.995 849.130 ;
        RECT 2786.990 849.130 2787.290 849.510 ;
        RECT 2787.910 849.130 2788.210 850.190 ;
        RECT 2835.750 849.810 2836.050 850.190 ;
        RECT 2916.710 850.190 2924.800 850.490 ;
        RECT 2916.710 849.810 2917.010 850.190 ;
        RECT 2835.750 849.510 2883.890 849.810 ;
        RECT 2786.990 848.830 2788.210 849.130 ;
        RECT 2883.590 849.130 2883.890 849.510 ;
        RECT 2884.510 849.510 2917.010 849.810 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
        RECT 2884.510 849.130 2884.810 849.510 ;
        RECT 2883.590 848.830 2884.810 849.130 ;
        RECT 2625.285 848.815 2625.615 848.830 ;
        RECT 2649.665 848.815 2649.995 848.830 ;
        RECT 1883.510 848.150 1931.690 848.450 ;
        RECT 1883.510 848.140 1883.890 848.150 ;
        RECT 1606.385 847.470 1641.890 847.770 ;
        RECT 1606.385 847.455 1606.715 847.470 ;
      LAYER via3 ;
        RECT 1226.660 2497.820 1226.980 2498.140 ;
        RECT 1226.660 850.180 1226.980 850.500 ;
        RECT 1345.340 850.860 1345.660 851.180 ;
        RECT 1345.340 849.500 1345.660 849.820 ;
        RECT 1883.540 850.180 1883.860 850.500 ;
        RECT 1883.540 848.140 1883.860 848.460 ;
      LAYER met4 ;
        RECT 1226.655 2497.815 1226.985 2498.145 ;
        RECT 1226.670 850.505 1226.970 2497.815 ;
        RECT 1345.335 850.855 1345.665 851.185 ;
        RECT 1226.655 850.175 1226.985 850.505 ;
        RECT 1345.350 849.825 1345.650 850.855 ;
        RECT 1883.535 850.175 1883.865 850.505 ;
        RECT 1345.335 849.495 1345.665 849.825 ;
<<<<<<< HEAD
        RECT 1441.935 849.495 1442.265 849.825 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1883.550 848.465 1883.850 850.175 ;
        RECT 1883.535 848.135 1883.865 848.465 ;
>>>>>>> re-updated local openlane
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1245.290 2498.900 1245.610 2498.960 ;
        RECT 2031.890 2498.900 2032.210 2498.960 ;
        RECT 1245.290 2498.760 2032.210 2498.900 ;
        RECT 1245.290 2498.700 1245.610 2498.760 ;
        RECT 2031.890 2498.700 2032.210 2498.760 ;
        RECT 2031.890 1089.940 2032.210 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2031.890 1089.800 2901.150 1089.940 ;
        RECT 2031.890 1089.740 2032.210 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 1245.320 2498.700 1245.580 2498.960 ;
        RECT 2031.920 2498.700 2032.180 2498.960 ;
        RECT 2031.920 1089.740 2032.180 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 1243.470 2498.730 1243.750 2500.000 ;
        RECT 1245.320 2498.730 1245.580 2498.990 ;
        RECT 1243.470 2498.670 1245.580 2498.730 ;
        RECT 2031.920 2498.670 2032.180 2498.990 ;
        RECT 1243.470 2498.590 1245.520 2498.670 ;
        RECT 1243.470 2496.000 1243.750 2498.590 ;
        RECT 2031.980 1090.030 2032.120 2498.670 ;
        RECT 2031.920 1089.710 2032.180 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1084.340 2924.800 1085.540 ;
=======
        RECT 1246.665 2498.140 1246.995 2498.145 ;
        RECT 1246.665 2498.130 1247.250 2498.140 ;
        RECT 1246.665 2497.830 1247.450 2498.130 ;
        RECT 1246.665 2497.820 1247.250 2497.830 ;
        RECT 1246.665 2497.815 1246.995 2497.820 ;
        RECT 1579.245 1086.450 1579.575 1086.465 ;
        RECT 1532.110 1086.150 1579.575 1086.450 ;
        RECT 1331.510 1085.090 1331.890 1085.100 ;
        RECT 1355.685 1085.090 1356.015 1085.105 ;
        RECT 1272.670 1084.790 1314.370 1085.090 ;
        RECT 1246.870 1084.410 1247.250 1084.420 ;
        RECT 1272.670 1084.410 1272.970 1084.790 ;
        RECT 1246.870 1084.110 1272.970 1084.410 ;
        RECT 1246.870 1084.100 1247.250 1084.110 ;
        RECT 1314.070 1083.730 1314.370 1084.790 ;
        RECT 1331.510 1084.790 1356.015 1085.090 ;
        RECT 1331.510 1084.780 1331.890 1084.790 ;
        RECT 1355.685 1084.775 1356.015 1084.790 ;
        RECT 1483.105 1085.090 1483.435 1085.105 ;
        RECT 1532.110 1085.090 1532.410 1086.150 ;
        RECT 1579.245 1086.135 1579.575 1086.150 ;
        RECT 1980.110 1086.450 1980.490 1086.460 ;
        RECT 2028.205 1086.450 2028.535 1086.465 ;
        RECT 1980.110 1086.150 2028.535 1086.450 ;
        RECT 1980.110 1086.140 1980.490 1086.150 ;
        RECT 2028.205 1086.135 2028.535 1086.150 ;
        RECT 2052.585 1085.770 2052.915 1085.785 ;
        RECT 2028.910 1085.470 2052.915 1085.770 ;
        RECT 1483.105 1084.790 1532.410 1085.090 ;
        RECT 1946.325 1085.090 1946.655 1085.105 ;
        RECT 1980.110 1085.090 1980.490 1085.100 ;
        RECT 1946.325 1084.790 1980.490 1085.090 ;
        RECT 1483.105 1084.775 1483.435 1084.790 ;
        RECT 1946.325 1084.775 1946.655 1084.790 ;
        RECT 1980.110 1084.780 1980.490 1084.790 ;
        RECT 1483.105 1084.410 1483.435 1084.425 ;
        RECT 1435.510 1084.110 1483.435 1084.410 ;
        RECT 1331.510 1083.730 1331.890 1083.740 ;
        RECT 1435.510 1083.730 1435.810 1084.110 ;
        RECT 1483.105 1084.095 1483.435 1084.110 ;
        RECT 1579.245 1084.410 1579.575 1084.425 ;
        RECT 1606.385 1084.410 1606.715 1084.425 ;
        RECT 1579.245 1084.110 1606.715 1084.410 ;
        RECT 1579.245 1084.095 1579.575 1084.110 ;
        RECT 1606.385 1084.095 1606.715 1084.110 ;
        RECT 1607.765 1084.410 1608.095 1084.425 ;
        RECT 1702.065 1084.410 1702.395 1084.425 ;
        RECT 1607.765 1084.110 1641.890 1084.410 ;
        RECT 1607.765 1084.095 1608.095 1084.110 ;
        RECT 1314.070 1083.430 1331.890 1083.730 ;
        RECT 1331.510 1083.420 1331.890 1083.430 ;
        RECT 1399.630 1083.430 1400.850 1083.730 ;
        RECT 1355.685 1083.050 1356.015 1083.065 ;
        RECT 1399.630 1083.050 1399.930 1083.430 ;
        RECT 1355.685 1082.750 1399.930 1083.050 ;
        RECT 1400.550 1083.050 1400.850 1083.430 ;
        RECT 1415.270 1083.430 1435.810 1083.730 ;
        RECT 1641.590 1083.730 1641.890 1084.110 ;
        RECT 1656.310 1084.110 1702.395 1084.410 ;
        RECT 1656.310 1083.730 1656.610 1084.110 ;
        RECT 1702.065 1084.095 1702.395 1084.110 ;
        RECT 1711.725 1084.410 1712.055 1084.425 ;
        RECT 1798.665 1084.410 1798.995 1084.425 ;
        RECT 1711.725 1084.110 1738.490 1084.410 ;
        RECT 1711.725 1084.095 1712.055 1084.110 ;
        RECT 1641.590 1083.430 1656.610 1083.730 ;
        RECT 1738.190 1083.730 1738.490 1084.110 ;
        RECT 1752.910 1084.110 1798.995 1084.410 ;
        RECT 1752.910 1083.730 1753.210 1084.110 ;
        RECT 1798.665 1084.095 1798.995 1084.110 ;
        RECT 1801.885 1084.410 1802.215 1084.425 ;
        RECT 1895.265 1084.410 1895.595 1084.425 ;
        RECT 1801.885 1084.110 1835.090 1084.410 ;
        RECT 1801.885 1084.095 1802.215 1084.110 ;
        RECT 1738.190 1083.430 1753.210 1083.730 ;
        RECT 1834.790 1083.730 1835.090 1084.110 ;
        RECT 1849.510 1084.110 1895.595 1084.410 ;
        RECT 1849.510 1083.730 1849.810 1084.110 ;
        RECT 1895.265 1084.095 1895.595 1084.110 ;
        RECT 2028.205 1084.410 2028.535 1084.425 ;
        RECT 2028.910 1084.410 2029.210 1085.470 ;
        RECT 2052.585 1085.455 2052.915 1085.470 ;
        RECT 2124.805 1085.090 2125.135 1085.105 ;
=======
        RECT 2900.825 1085.090 2901.155 1085.105 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
<<<<<<< HEAD
        RECT 2884.510 1083.730 2884.810 1084.110 ;
        RECT 2883.590 1083.430 2884.810 1083.730 ;
        RECT 2052.585 1083.415 2052.915 1083.430 ;
        RECT 1895.265 1082.070 1931.690 1082.370 ;
        RECT 1895.265 1082.055 1895.595 1082.070 ;
      LAYER via3 ;
        RECT 1246.900 2497.820 1247.220 2498.140 ;
        RECT 1246.900 1084.100 1247.220 1084.420 ;
        RECT 1331.540 1084.780 1331.860 1085.100 ;
        RECT 1980.140 1086.140 1980.460 1086.460 ;
        RECT 1980.140 1084.780 1980.460 1085.100 ;
        RECT 1331.540 1083.420 1331.860 1083.740 ;
      LAYER met4 ;
        RECT 1246.895 2497.815 1247.225 2498.145 ;
        RECT 1246.910 1084.425 1247.210 2497.815 ;
        RECT 1980.135 1086.135 1980.465 1086.465 ;
        RECT 1980.150 1085.105 1980.450 1086.135 ;
        RECT 1331.535 1084.775 1331.865 1085.105 ;
        RECT 1980.135 1084.775 1980.465 1085.105 ;
        RECT 1246.895 1084.095 1247.225 1084.425 ;
        RECT 1331.550 1083.745 1331.850 1084.775 ;
        RECT 1331.535 1083.415 1331.865 1083.745 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1264.685 2492.625 1264.855 2496.535 ;
      LAYER mcon ;
        RECT 1264.685 2496.365 1264.855 2496.535 ;
      LAYER met1 ;
        RECT 1264.610 2496.520 1264.930 2496.580 ;
        RECT 1264.415 2496.380 1264.930 2496.520 ;
        RECT 1264.610 2496.320 1264.930 2496.380 ;
        RECT 1264.625 2492.780 1264.915 2492.825 ;
        RECT 2100.890 2492.780 2101.210 2492.840 ;
        RECT 1264.625 2492.640 2101.210 2492.780 ;
        RECT 1264.625 2492.595 1264.915 2492.640 ;
        RECT 2100.890 2492.580 2101.210 2492.640 ;
        RECT 2100.890 1324.540 2101.210 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 2100.890 1324.400 2901.150 1324.540 ;
        RECT 2100.890 1324.340 2101.210 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 1264.640 2496.320 1264.900 2496.580 ;
        RECT 2100.920 2492.580 2101.180 2492.840 ;
        RECT 2100.920 1324.340 2101.180 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 1262.790 2496.690 1263.070 2500.000 ;
        RECT 1262.790 2496.610 1264.840 2496.690 ;
        RECT 1262.790 2496.550 1264.900 2496.610 ;
        RECT 1262.790 2496.000 1263.070 2496.550 ;
        RECT 1264.640 2496.290 1264.900 2496.550 ;
        RECT 2100.920 2492.550 2101.180 2492.870 ;
        RECT 2100.980 1324.630 2101.120 2492.550 ;
        RECT 2100.920 1324.310 2101.180 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2919.700 1318.940 2924.800 1320.140 ;
=======
        RECT 1267.365 2498.130 1267.695 2498.145 ;
        RECT 1268.950 2498.130 1269.330 2498.140 ;
        RECT 1267.365 2497.830 1269.330 2498.130 ;
        RECT 1267.365 2497.815 1267.695 2497.830 ;
        RECT 1268.950 2497.820 1269.330 2497.830 ;
        RECT 1980.110 1321.050 1980.490 1321.060 ;
        RECT 2028.205 1321.050 2028.535 1321.065 ;
        RECT 1980.110 1320.750 2028.535 1321.050 ;
        RECT 1980.110 1320.740 1980.490 1320.750 ;
        RECT 2028.205 1320.735 2028.535 1320.750 ;
        RECT 1268.950 1320.370 1269.330 1320.380 ;
        RECT 2052.585 1320.370 2052.915 1320.385 ;
        RECT 1268.950 1320.070 1365.890 1320.370 ;
        RECT 1268.950 1320.060 1269.330 1320.070 ;
        RECT 1365.590 1319.010 1365.890 1320.070 ;
        RECT 2028.910 1320.070 2052.915 1320.370 ;
        RECT 1448.605 1319.690 1448.935 1319.705 ;
        RECT 1946.325 1319.690 1946.655 1319.705 ;
        RECT 1980.110 1319.690 1980.490 1319.700 ;
        RECT 1448.605 1319.390 1511.250 1319.690 ;
        RECT 1448.605 1319.375 1448.935 1319.390 ;
        RECT 1448.605 1319.010 1448.935 1319.025 ;
        RECT 1365.590 1318.710 1448.935 1319.010 ;
        RECT 1448.605 1318.695 1448.935 1318.710 ;
        RECT 1510.950 1318.330 1511.250 1319.390 ;
        RECT 1946.325 1319.390 1980.490 1319.690 ;
        RECT 1946.325 1319.375 1946.655 1319.390 ;
        RECT 1980.110 1319.380 1980.490 1319.390 ;
        RECT 1606.385 1319.010 1606.715 1319.025 ;
        RECT 1559.710 1318.710 1606.715 1319.010 ;
        RECT 1559.710 1318.330 1560.010 1318.710 ;
        RECT 1606.385 1318.695 1606.715 1318.710 ;
        RECT 1607.765 1319.010 1608.095 1319.025 ;
        RECT 1702.065 1319.010 1702.395 1319.025 ;
        RECT 1607.765 1318.710 1641.890 1319.010 ;
        RECT 1607.765 1318.695 1608.095 1318.710 ;
        RECT 1510.950 1318.030 1560.010 1318.330 ;
        RECT 1641.590 1318.330 1641.890 1318.710 ;
        RECT 1656.310 1318.710 1702.395 1319.010 ;
        RECT 1656.310 1318.330 1656.610 1318.710 ;
        RECT 1702.065 1318.695 1702.395 1318.710 ;
        RECT 1711.725 1319.010 1712.055 1319.025 ;
        RECT 1798.665 1319.010 1798.995 1319.025 ;
        RECT 1711.725 1318.710 1738.490 1319.010 ;
        RECT 1711.725 1318.695 1712.055 1318.710 ;
        RECT 1641.590 1318.030 1656.610 1318.330 ;
        RECT 1738.190 1318.330 1738.490 1318.710 ;
        RECT 1752.910 1318.710 1798.995 1319.010 ;
        RECT 1752.910 1318.330 1753.210 1318.710 ;
        RECT 1798.665 1318.695 1798.995 1318.710 ;
        RECT 1801.885 1319.010 1802.215 1319.025 ;
        RECT 1895.265 1319.010 1895.595 1319.025 ;
        RECT 1801.885 1318.710 1835.090 1319.010 ;
        RECT 1801.885 1318.695 1802.215 1318.710 ;
        RECT 1738.190 1318.030 1753.210 1318.330 ;
        RECT 1834.790 1318.330 1835.090 1318.710 ;
        RECT 1849.510 1318.710 1895.595 1319.010 ;
        RECT 1849.510 1318.330 1849.810 1318.710 ;
        RECT 1895.265 1318.695 1895.595 1318.710 ;
        RECT 2028.205 1319.010 2028.535 1319.025 ;
        RECT 2028.910 1319.010 2029.210 1320.070 ;
        RECT 2052.585 1320.055 2052.915 1320.070 ;
        RECT 2124.805 1319.690 2125.135 1319.705 ;
=======
        RECT 2900.825 1319.690 2901.155 1319.705 ;
>>>>>>> re-updated local openlane
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
<<<<<<< HEAD
        RECT 2884.510 1318.330 2884.810 1318.710 ;
        RECT 2883.590 1318.030 2884.810 1318.330 ;
        RECT 2052.585 1318.015 2052.915 1318.030 ;
        RECT 1895.265 1316.670 1931.690 1316.970 ;
        RECT 1895.265 1316.655 1895.595 1316.670 ;
      LAYER via3 ;
        RECT 1268.980 2497.820 1269.300 2498.140 ;
        RECT 1980.140 1320.740 1980.460 1321.060 ;
        RECT 1268.980 1320.060 1269.300 1320.380 ;
        RECT 1980.140 1319.380 1980.460 1319.700 ;
      LAYER met4 ;
        RECT 1268.975 2497.815 1269.305 2498.145 ;
        RECT 1268.990 1320.385 1269.290 2497.815 ;
        RECT 1980.135 1320.735 1980.465 1321.065 ;
        RECT 1268.975 1320.055 1269.305 1320.385 ;
        RECT 1980.150 1319.705 1980.450 1320.735 ;
        RECT 1980.135 1319.375 1980.465 1319.705 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1282.090 2507.060 1282.410 2507.120 ;
        RECT 2080.190 2507.060 2080.510 2507.120 ;
        RECT 1282.090 2506.920 2080.510 2507.060 ;
        RECT 1282.090 2506.860 1282.410 2506.920 ;
        RECT 2080.190 2506.860 2080.510 2506.920 ;
        RECT 2080.190 1559.140 2080.510 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2080.190 1559.000 2901.150 1559.140 ;
        RECT 2080.190 1558.940 2080.510 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 1282.120 2506.860 1282.380 2507.120 ;
        RECT 2080.220 2506.860 2080.480 2507.120 ;
        RECT 2080.220 1558.940 2080.480 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 1282.120 2506.830 1282.380 2507.150 ;
        RECT 2080.220 2506.830 2080.480 2507.150 ;
        RECT 1282.180 2500.000 1282.320 2506.830 ;
        RECT 1282.110 2496.000 1282.390 2500.000 ;
        RECT 2080.280 1559.230 2080.420 2506.830 ;
        RECT 2080.220 1558.910 2080.480 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1553.540 2924.800 1554.740 ;
=======
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1301.410 2513.860 1301.730 2513.920 ;
        RECT 1942.190 2513.860 1942.510 2513.920 ;
        RECT 1301.410 2513.720 1942.510 2513.860 ;
        RECT 1301.410 2513.660 1301.730 2513.720 ;
        RECT 1942.190 2513.660 1942.510 2513.720 ;
        RECT 1945.410 1793.740 1945.730 1793.800 ;
        RECT 2900.830 1793.740 2901.150 1793.800 ;
        RECT 1945.410 1793.600 2901.150 1793.740 ;
        RECT 1945.410 1793.540 1945.730 1793.600 ;
        RECT 2900.830 1793.540 2901.150 1793.600 ;
      LAYER via ;
        RECT 1301.440 2513.660 1301.700 2513.920 ;
        RECT 1942.220 2513.660 1942.480 2513.920 ;
        RECT 1945.440 1793.540 1945.700 1793.800 ;
        RECT 2900.860 1793.540 2901.120 1793.800 ;
      LAYER met2 ;
        RECT 1301.440 2513.630 1301.700 2513.950 ;
        RECT 1942.220 2513.630 1942.480 2513.950 ;
        RECT 1301.500 2500.000 1301.640 2513.630 ;
        RECT 1301.430 2496.000 1301.710 2500.000 ;
        RECT 1942.280 1793.570 1942.420 2513.630 ;
        RECT 1945.440 1793.570 1945.700 1793.830 ;
        RECT 1942.280 1793.510 1945.700 1793.570 ;
        RECT 2900.860 1793.510 2901.120 1793.830 ;
        RECT 1942.280 1793.430 1945.640 1793.510 ;
        RECT 2900.920 1789.605 2901.060 1793.510 ;
        RECT 2900.850 1789.235 2901.130 1789.605 ;
      LAYER via2 ;
        RECT 2900.850 1789.280 2901.130 1789.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 1788.820 2924.800 1790.020 ;
=======
        RECT 2900.825 1789.570 2901.155 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.825 1789.270 2924.800 1789.570 ;
        RECT 2900.825 1789.255 2901.155 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1320.730 2514.200 1321.050 2514.260 ;
        RECT 1942.650 2514.200 1942.970 2514.260 ;
        RECT 1320.730 2514.060 1942.970 2514.200 ;
        RECT 1320.730 2514.000 1321.050 2514.060 ;
        RECT 1942.650 2514.000 1942.970 2514.060 ;
        RECT 1945.410 2028.340 1945.730 2028.400 ;
        RECT 2900.830 2028.340 2901.150 2028.400 ;
        RECT 1945.410 2028.200 2901.150 2028.340 ;
        RECT 1945.410 2028.140 1945.730 2028.200 ;
        RECT 2900.830 2028.140 2901.150 2028.200 ;
      LAYER via ;
        RECT 1320.760 2514.000 1321.020 2514.260 ;
        RECT 1942.680 2514.000 1942.940 2514.260 ;
        RECT 1945.440 2028.140 1945.700 2028.400 ;
        RECT 2900.860 2028.140 2901.120 2028.400 ;
      LAYER met2 ;
        RECT 1320.760 2513.970 1321.020 2514.290 ;
        RECT 1942.680 2513.970 1942.940 2514.290 ;
        RECT 1320.820 2500.000 1320.960 2513.970 ;
        RECT 1320.750 2496.000 1321.030 2500.000 ;
        RECT 1942.740 2069.650 1942.880 2513.970 ;
        RECT 1942.740 2069.510 1943.800 2069.650 ;
        RECT 1943.660 2028.170 1943.800 2069.510 ;
        RECT 1945.440 2028.170 1945.700 2028.430 ;
        RECT 1943.660 2028.110 1945.700 2028.170 ;
        RECT 2900.860 2028.110 2901.120 2028.430 ;
        RECT 1943.660 2028.030 1945.640 2028.110 ;
        RECT 2900.920 2024.205 2901.060 2028.110 ;
        RECT 2900.850 2023.835 2901.130 2024.205 ;
      LAYER via2 ;
        RECT 2900.850 2023.880 2901.130 2024.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2023.420 2924.800 2024.620 ;
=======
        RECT 2900.825 2024.170 2901.155 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.825 2023.870 2924.800 2024.170 ;
        RECT 2900.825 2023.855 2901.155 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1340.050 2517.260 1340.370 2517.320 ;
        RECT 1943.110 2517.260 1943.430 2517.320 ;
        RECT 1340.050 2517.120 1943.430 2517.260 ;
        RECT 1340.050 2517.060 1340.370 2517.120 ;
        RECT 1943.110 2517.060 1943.430 2517.120 ;
        RECT 1945.410 2262.940 1945.730 2263.000 ;
        RECT 2900.830 2262.940 2901.150 2263.000 ;
        RECT 1945.410 2262.800 2901.150 2262.940 ;
        RECT 1945.410 2262.740 1945.730 2262.800 ;
        RECT 2900.830 2262.740 2901.150 2262.800 ;
      LAYER via ;
        RECT 1340.080 2517.060 1340.340 2517.320 ;
        RECT 1943.140 2517.060 1943.400 2517.320 ;
        RECT 1945.440 2262.740 1945.700 2263.000 ;
        RECT 2900.860 2262.740 2901.120 2263.000 ;
      LAYER met2 ;
        RECT 1340.080 2517.030 1340.340 2517.350 ;
        RECT 1943.140 2517.030 1943.400 2517.350 ;
        RECT 1340.140 2500.000 1340.280 2517.030 ;
        RECT 1340.070 2496.000 1340.350 2500.000 ;
        RECT 1943.200 2262.770 1943.340 2517.030 ;
        RECT 1945.440 2262.770 1945.700 2263.030 ;
        RECT 1943.200 2262.710 1945.700 2262.770 ;
        RECT 2900.860 2262.710 2901.120 2263.030 ;
        RECT 1943.200 2262.630 1945.640 2262.710 ;
        RECT 2900.920 2258.805 2901.060 2262.710 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2919.700 2258.020 2924.800 2259.220 ;
=======
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 0.300 ;
=======
      LAYER met1 ;
        RECT 634.410 1680.180 634.730 1680.240 ;
        RECT 1321.190 1680.180 1321.510 1680.240 ;
        RECT 634.410 1680.040 1321.510 1680.180 ;
        RECT 634.410 1679.980 634.730 1680.040 ;
        RECT 1321.190 1679.980 1321.510 1680.040 ;
      LAYER via ;
        RECT 634.440 1679.980 634.700 1680.240 ;
        RECT 1321.220 1679.980 1321.480 1680.240 ;
      LAYER met2 ;
        RECT 1321.210 1700.000 1321.490 1704.000 ;
        RECT 1321.280 1680.270 1321.420 1700.000 ;
        RECT 634.440 1679.950 634.700 1680.270 ;
        RECT 1321.220 1679.950 1321.480 1680.270 ;
        RECT 634.500 17.410 634.640 1679.950 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1802.350 1683.920 1802.670 1683.980 ;
        RECT 1806.950 1683.920 1807.270 1683.980 ;
        RECT 1802.350 1683.780 1807.270 1683.920 ;
        RECT 1802.350 1683.720 1802.670 1683.780 ;
        RECT 1806.950 1683.720 1807.270 1683.780 ;
        RECT 1806.950 44.780 1807.270 44.840 ;
        RECT 2417.370 44.780 2417.690 44.840 ;
        RECT 1806.950 44.640 2417.690 44.780 ;
        RECT 1806.950 44.580 1807.270 44.640 ;
        RECT 2417.370 44.580 2417.690 44.640 ;
      LAYER via ;
        RECT 1802.380 1683.720 1802.640 1683.980 ;
        RECT 1806.980 1683.720 1807.240 1683.980 ;
        RECT 1806.980 44.580 1807.240 44.840 ;
        RECT 2417.400 44.580 2417.660 44.840 ;
      LAYER met2 ;
        RECT 1802.370 1700.000 1802.650 1704.000 ;
        RECT 1802.440 1684.010 1802.580 1700.000 ;
        RECT 1802.380 1683.690 1802.640 1684.010 ;
        RECT 1806.980 1683.690 1807.240 1684.010 ;
        RECT 1807.040 44.870 1807.180 1683.690 ;
        RECT 1806.980 44.550 1807.240 44.870 ;
        RECT 2417.400 44.550 2417.660 44.870 ;
        RECT 2417.460 2.400 2417.600 44.550 ;
=======
      LAYER li1 ;
        RECT 2415.145 48.365 2415.315 96.475 ;
      LAYER mcon ;
        RECT 2415.145 96.305 2415.315 96.475 ;
      LAYER met1 ;
        RECT 1805.110 1680.180 1805.430 1680.240 ;
        RECT 2415.070 1680.180 2415.390 1680.240 ;
        RECT 1805.110 1680.040 2415.390 1680.180 ;
        RECT 1805.110 1679.980 1805.430 1680.040 ;
        RECT 2415.070 1679.980 2415.390 1680.040 ;
        RECT 2415.070 96.460 2415.390 96.520 ;
        RECT 2415.070 96.320 2415.585 96.460 ;
        RECT 2415.070 96.260 2415.390 96.320 ;
        RECT 2415.085 48.520 2415.375 48.565 ;
        RECT 2417.370 48.520 2417.690 48.580 ;
        RECT 2415.085 48.380 2417.690 48.520 ;
        RECT 2415.085 48.335 2415.375 48.380 ;
        RECT 2417.370 48.320 2417.690 48.380 ;
        RECT 2416.910 2.960 2417.230 3.020 ;
        RECT 2417.370 2.960 2417.690 3.020 ;
        RECT 2416.910 2.820 2417.690 2.960 ;
        RECT 2416.910 2.760 2417.230 2.820 ;
        RECT 2417.370 2.760 2417.690 2.820 ;
      LAYER via ;
        RECT 1805.140 1679.980 1805.400 1680.240 ;
        RECT 2415.100 1679.980 2415.360 1680.240 ;
        RECT 2415.100 96.260 2415.360 96.520 ;
        RECT 2417.400 48.320 2417.660 48.580 ;
        RECT 2416.940 2.760 2417.200 3.020 ;
        RECT 2417.400 2.760 2417.660 3.020 ;
      LAYER met2 ;
        RECT 1805.130 1700.000 1805.410 1704.000 ;
        RECT 1805.200 1680.270 1805.340 1700.000 ;
        RECT 1805.140 1679.950 1805.400 1680.270 ;
        RECT 2415.100 1679.950 2415.360 1680.270 ;
        RECT 2415.160 96.550 2415.300 1679.950 ;
        RECT 2415.100 96.230 2415.360 96.550 ;
        RECT 2417.400 48.290 2417.660 48.610 ;
        RECT 2417.460 48.010 2417.600 48.290 ;
        RECT 2417.000 47.870 2417.600 48.010 ;
        RECT 2417.000 3.050 2417.140 47.870 ;
        RECT 2416.940 2.730 2417.200 3.050 ;
        RECT 2417.400 2.730 2417.660 3.050 ;
        RECT 2417.460 2.400 2417.600 2.730 ;
>>>>>>> re-updated local openlane
        RECT 2417.250 -4.800 2417.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2434.730 -4.800 2435.290 0.300 ;
=======
        RECT 1807.430 1700.410 1807.710 1704.000 ;
        RECT 1806.580 1700.270 1807.710 1700.410 ;
        RECT 1806.580 48.125 1806.720 1700.270 ;
        RECT 1807.430 1700.000 1807.710 1700.270 ;
        RECT 1806.510 47.755 1806.790 48.125 ;
        RECT 2434.870 47.755 2435.150 48.125 ;
        RECT 2434.940 2.400 2435.080 47.755 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
      LAYER via2 ;
        RECT 1806.510 47.800 1806.790 48.080 ;
        RECT 2434.870 47.800 2435.150 48.080 ;
      LAYER met3 ;
        RECT 1806.485 48.090 1806.815 48.105 ;
        RECT 2434.845 48.090 2435.175 48.105 ;
        RECT 1806.485 47.790 2435.175 48.090 ;
        RECT 1806.485 47.775 1806.815 47.790 ;
        RECT 2434.845 47.775 2435.175 47.790 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1807.870 1683.920 1808.190 1683.980 ;
        RECT 1809.710 1683.920 1810.030 1683.980 ;
        RECT 1807.870 1683.780 1810.030 1683.920 ;
        RECT 1807.870 1683.720 1808.190 1683.780 ;
        RECT 1809.710 1683.720 1810.030 1683.780 ;
        RECT 1807.870 1652.640 1808.190 1652.700 ;
        RECT 2428.870 1652.640 2429.190 1652.700 ;
        RECT 1807.870 1652.500 2429.190 1652.640 ;
        RECT 1807.870 1652.440 1808.190 1652.500 ;
        RECT 2428.870 1652.440 2429.190 1652.500 ;
        RECT 2428.870 35.940 2429.190 36.000 ;
        RECT 2434.850 35.940 2435.170 36.000 ;
        RECT 2428.870 35.800 2435.170 35.940 ;
        RECT 2428.870 35.740 2429.190 35.800 ;
        RECT 2434.850 35.740 2435.170 35.800 ;
      LAYER via ;
        RECT 1807.900 1683.720 1808.160 1683.980 ;
        RECT 1809.740 1683.720 1810.000 1683.980 ;
        RECT 1807.900 1652.440 1808.160 1652.700 ;
        RECT 2428.900 1652.440 2429.160 1652.700 ;
        RECT 2428.900 35.740 2429.160 36.000 ;
        RECT 2434.880 35.740 2435.140 36.000 ;
      LAYER met2 ;
        RECT 1809.730 1700.000 1810.010 1704.000 ;
        RECT 1809.800 1684.010 1809.940 1700.000 ;
        RECT 1807.900 1683.690 1808.160 1684.010 ;
        RECT 1809.740 1683.690 1810.000 1684.010 ;
        RECT 1807.960 1652.730 1808.100 1683.690 ;
        RECT 1807.900 1652.410 1808.160 1652.730 ;
        RECT 2428.900 1652.410 2429.160 1652.730 ;
        RECT 2428.960 36.030 2429.100 1652.410 ;
        RECT 2428.900 35.710 2429.160 36.030 ;
        RECT 2434.880 35.710 2435.140 36.030 ;
        RECT 2434.940 2.400 2435.080 35.710 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2452.670 -4.800 2453.230 0.300 ;
=======
        RECT 1812.030 1700.410 1812.310 1704.000 ;
        RECT 1812.030 1700.270 1813.620 1700.410 ;
        RECT 1812.030 1700.000 1812.310 1700.270 ;
        RECT 1813.480 47.445 1813.620 1700.270 ;
        RECT 1813.410 47.075 1813.690 47.445 ;
        RECT 2452.810 47.075 2453.090 47.445 ;
        RECT 2452.880 2.400 2453.020 47.075 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
      LAYER via2 ;
        RECT 1813.410 47.120 1813.690 47.400 ;
        RECT 2452.810 47.120 2453.090 47.400 ;
      LAYER met3 ;
        RECT 1813.385 47.410 1813.715 47.425 ;
        RECT 2452.785 47.410 2453.115 47.425 ;
        RECT 1813.385 47.110 2453.115 47.410 ;
        RECT 1813.385 47.095 1813.715 47.110 ;
        RECT 2452.785 47.095 2453.115 47.110 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1814.770 1666.580 1815.090 1666.640 ;
        RECT 2449.570 1666.580 2449.890 1666.640 ;
        RECT 1814.770 1666.440 2449.890 1666.580 ;
        RECT 1814.770 1666.380 1815.090 1666.440 ;
        RECT 2449.570 1666.380 2449.890 1666.440 ;
        RECT 2449.570 62.120 2449.890 62.180 ;
        RECT 2452.790 62.120 2453.110 62.180 ;
        RECT 2449.570 61.980 2453.110 62.120 ;
        RECT 2449.570 61.920 2449.890 61.980 ;
        RECT 2452.790 61.920 2453.110 61.980 ;
      LAYER via ;
        RECT 1814.800 1666.380 1815.060 1666.640 ;
        RECT 2449.600 1666.380 2449.860 1666.640 ;
        RECT 2449.600 61.920 2449.860 62.180 ;
        RECT 2452.820 61.920 2453.080 62.180 ;
      LAYER met2 ;
        RECT 1814.790 1700.000 1815.070 1704.000 ;
        RECT 1814.860 1666.670 1815.000 1700.000 ;
        RECT 1814.800 1666.350 1815.060 1666.670 ;
        RECT 2449.600 1666.350 2449.860 1666.670 ;
        RECT 2449.660 62.210 2449.800 1666.350 ;
        RECT 2449.600 61.890 2449.860 62.210 ;
        RECT 2452.820 61.890 2453.080 62.210 ;
        RECT 2452.880 2.400 2453.020 61.890 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1819.830 1683.920 1820.150 1683.980 ;
        RECT 1820.750 1683.920 1821.070 1683.980 ;
        RECT 1819.830 1683.780 1821.070 1683.920 ;
        RECT 1819.830 1683.720 1820.150 1683.780 ;
        RECT 1820.750 1683.720 1821.070 1683.780 ;
        RECT 1820.750 51.580 1821.070 51.640 ;
        RECT 2470.730 51.580 2471.050 51.640 ;
        RECT 1820.750 51.440 2471.050 51.580 ;
        RECT 1820.750 51.380 1821.070 51.440 ;
        RECT 2470.730 51.380 2471.050 51.440 ;
      LAYER via ;
        RECT 1819.860 1683.720 1820.120 1683.980 ;
        RECT 1820.780 1683.720 1821.040 1683.980 ;
        RECT 1820.780 51.380 1821.040 51.640 ;
        RECT 2470.760 51.380 2471.020 51.640 ;
      LAYER met2 ;
        RECT 1819.850 1700.000 1820.130 1704.000 ;
        RECT 1819.920 1684.010 1820.060 1700.000 ;
        RECT 1819.860 1683.690 1820.120 1684.010 ;
        RECT 1820.780 1683.690 1821.040 1684.010 ;
        RECT 1820.840 51.670 1820.980 1683.690 ;
        RECT 1820.780 51.350 1821.040 51.670 ;
        RECT 2470.760 51.350 2471.020 51.670 ;
        RECT 2470.820 2.400 2470.960 51.350 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 0.300 ;
=======
      LAYER li1 ;
        RECT 1873.725 21.165 1873.895 23.715 ;
      LAYER mcon ;
        RECT 1873.725 23.545 1873.895 23.715 ;
      LAYER met1 ;
        RECT 1823.050 1677.460 1823.370 1677.520 ;
        RECT 1827.650 1677.460 1827.970 1677.520 ;
        RECT 1823.050 1677.320 1827.970 1677.460 ;
        RECT 1823.050 1677.260 1823.370 1677.320 ;
        RECT 1827.650 1677.260 1827.970 1677.320 ;
        RECT 1873.665 23.700 1873.955 23.745 ;
        RECT 1833.260 23.560 1873.955 23.700 ;
        RECT 1827.650 23.360 1827.970 23.420 ;
        RECT 1833.260 23.360 1833.400 23.560 ;
        RECT 1873.665 23.515 1873.955 23.560 ;
        RECT 1827.650 23.220 1833.400 23.360 ;
        RECT 1827.650 23.160 1827.970 23.220 ;
        RECT 1873.665 21.320 1873.955 21.365 ;
        RECT 2488.670 21.320 2488.990 21.380 ;
        RECT 1873.665 21.180 2488.990 21.320 ;
        RECT 1873.665 21.135 1873.955 21.180 ;
        RECT 2488.670 21.120 2488.990 21.180 ;
      LAYER via ;
        RECT 1823.080 1677.260 1823.340 1677.520 ;
        RECT 1827.680 1677.260 1827.940 1677.520 ;
        RECT 1827.680 23.160 1827.940 23.420 ;
        RECT 2488.700 21.120 2488.960 21.380 ;
      LAYER met2 ;
        RECT 1821.690 1700.410 1821.970 1704.000 ;
        RECT 1821.690 1700.270 1823.280 1700.410 ;
        RECT 1821.690 1700.000 1821.970 1700.270 ;
        RECT 1823.140 1677.550 1823.280 1700.270 ;
        RECT 1823.080 1677.230 1823.340 1677.550 ;
        RECT 1827.680 1677.230 1827.940 1677.550 ;
        RECT 1827.740 23.450 1827.880 1677.230 ;
        RECT 1827.680 23.130 1827.940 23.450 ;
        RECT 2488.700 21.090 2488.960 21.410 ;
        RECT 2488.760 2.400 2488.900 21.090 ;
=======
      LAYER met1 ;
        RECT 1824.430 1659.440 1824.750 1659.500 ;
        RECT 2484.070 1659.440 2484.390 1659.500 ;
        RECT 1824.430 1659.300 2484.390 1659.440 ;
        RECT 1824.430 1659.240 1824.750 1659.300 ;
        RECT 2484.070 1659.240 2484.390 1659.300 ;
      LAYER via ;
        RECT 1824.460 1659.240 1824.720 1659.500 ;
        RECT 2484.100 1659.240 2484.360 1659.500 ;
      LAYER met2 ;
        RECT 1824.450 1700.000 1824.730 1704.000 ;
        RECT 1824.520 1659.530 1824.660 1700.000 ;
        RECT 1824.460 1659.210 1824.720 1659.530 ;
        RECT 2484.100 1659.210 2484.360 1659.530 ;
        RECT 2484.160 16.730 2484.300 1659.210 ;
        RECT 2484.160 16.590 2488.900 16.730 ;
        RECT 2488.760 2.400 2488.900 16.590 ;
>>>>>>> re-updated local openlane
        RECT 2488.550 -4.800 2489.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1829.490 1683.920 1829.810 1683.980 ;
        RECT 1833.630 1683.920 1833.950 1683.980 ;
        RECT 1829.490 1683.780 1833.950 1683.920 ;
        RECT 1829.490 1683.720 1829.810 1683.780 ;
        RECT 1833.630 1683.720 1833.950 1683.780 ;
        RECT 1833.630 1639.040 1833.950 1639.100 ;
        RECT 2504.770 1639.040 2505.090 1639.100 ;
        RECT 1833.630 1638.900 2505.090 1639.040 ;
        RECT 1833.630 1638.840 1833.950 1638.900 ;
        RECT 2504.770 1638.840 2505.090 1638.900 ;
      LAYER via ;
        RECT 1829.520 1683.720 1829.780 1683.980 ;
        RECT 1833.660 1683.720 1833.920 1683.980 ;
        RECT 1833.660 1638.840 1833.920 1639.100 ;
        RECT 2504.800 1638.840 2505.060 1639.100 ;
      LAYER met2 ;
        RECT 1829.510 1700.000 1829.790 1704.000 ;
        RECT 1829.580 1684.010 1829.720 1700.000 ;
        RECT 1829.520 1683.690 1829.780 1684.010 ;
        RECT 1833.660 1683.690 1833.920 1684.010 ;
        RECT 1833.720 1639.130 1833.860 1683.690 ;
        RECT 1833.660 1638.810 1833.920 1639.130 ;
        RECT 2504.800 1638.810 2505.060 1639.130 ;
        RECT 2504.860 16.730 2505.000 1638.810 ;
        RECT 2504.860 16.590 2506.380 16.730 ;
        RECT 2506.240 2.400 2506.380 16.590 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1834.090 1631.900 1834.410 1631.960 ;
        RECT 2518.570 1631.900 2518.890 1631.960 ;
        RECT 1834.090 1631.760 2518.890 1631.900 ;
        RECT 1834.090 1631.700 1834.410 1631.760 ;
        RECT 2518.570 1631.700 2518.890 1631.760 ;
      LAYER via ;
        RECT 1834.120 1631.700 1834.380 1631.960 ;
        RECT 2518.600 1631.700 2518.860 1631.960 ;
      LAYER met2 ;
        RECT 1834.110 1700.000 1834.390 1704.000 ;
        RECT 1834.180 1631.990 1834.320 1700.000 ;
        RECT 1834.120 1631.670 1834.380 1631.990 ;
        RECT 2518.600 1631.670 2518.860 1631.990 ;
        RECT 2518.660 16.730 2518.800 1631.670 ;
        RECT 2518.660 16.590 2524.320 16.730 ;
        RECT 2524.180 2.400 2524.320 16.590 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 0.300 ;
=======
      LAYER li1 ;
        RECT 2539.345 1635.485 2539.515 1645.855 ;
        RECT 2539.345 1538.925 2539.515 1587.035 ;
        RECT 2539.345 1442.025 2539.515 1490.475 ;
        RECT 2539.345 766.105 2539.515 814.215 ;
        RECT 2539.345 669.545 2539.515 717.655 ;
        RECT 2539.345 572.645 2539.515 620.755 ;
        RECT 2539.345 476.085 2539.515 524.195 ;
        RECT 2539.345 379.525 2539.515 427.635 ;
        RECT 2539.345 282.965 2539.515 331.075 ;
        RECT 2539.345 186.405 2539.515 234.515 ;
        RECT 2539.345 89.845 2539.515 137.955 ;
      LAYER mcon ;
        RECT 2539.345 1645.685 2539.515 1645.855 ;
        RECT 2539.345 1586.865 2539.515 1587.035 ;
        RECT 2539.345 1490.305 2539.515 1490.475 ;
        RECT 2539.345 814.045 2539.515 814.215 ;
        RECT 2539.345 717.485 2539.515 717.655 ;
        RECT 2539.345 620.585 2539.515 620.755 ;
        RECT 2539.345 524.025 2539.515 524.195 ;
        RECT 2539.345 427.465 2539.515 427.635 ;
        RECT 2539.345 330.905 2539.515 331.075 ;
        RECT 2539.345 234.345 2539.515 234.515 ;
        RECT 2539.345 137.785 2539.515 137.955 ;
      LAYER met1 ;
        RECT 1835.470 1683.920 1835.790 1683.980 ;
        RECT 1839.150 1683.920 1839.470 1683.980 ;
        RECT 1835.470 1683.780 1839.470 1683.920 ;
        RECT 1835.470 1683.720 1835.790 1683.780 ;
        RECT 1839.150 1683.720 1839.470 1683.780 ;
        RECT 1835.470 1645.840 1835.790 1645.900 ;
        RECT 2539.285 1645.840 2539.575 1645.885 ;
        RECT 1835.470 1645.700 2539.575 1645.840 ;
        RECT 1835.470 1645.640 1835.790 1645.700 ;
        RECT 2539.285 1645.655 2539.575 1645.700 ;
        RECT 2539.270 1635.640 2539.590 1635.700 ;
        RECT 2539.075 1635.500 2539.590 1635.640 ;
        RECT 2539.270 1635.440 2539.590 1635.500 ;
        RECT 2539.270 1587.020 2539.590 1587.080 ;
        RECT 2539.075 1586.880 2539.590 1587.020 ;
        RECT 2539.270 1586.820 2539.590 1586.880 ;
        RECT 2539.270 1539.080 2539.590 1539.140 ;
        RECT 2539.075 1538.940 2539.590 1539.080 ;
        RECT 2539.270 1538.880 2539.590 1538.940 ;
        RECT 2539.270 1490.460 2539.590 1490.520 ;
        RECT 2539.075 1490.320 2539.590 1490.460 ;
        RECT 2539.270 1490.260 2539.590 1490.320 ;
        RECT 2539.270 1442.180 2539.590 1442.240 ;
        RECT 2539.075 1442.040 2539.590 1442.180 ;
        RECT 2539.270 1441.980 2539.590 1442.040 ;
        RECT 2539.270 1345.620 2539.590 1345.680 ;
        RECT 2540.190 1345.620 2540.510 1345.680 ;
        RECT 2539.270 1345.480 2540.510 1345.620 ;
        RECT 2539.270 1345.420 2539.590 1345.480 ;
        RECT 2540.190 1345.420 2540.510 1345.480 ;
        RECT 2539.270 1249.060 2539.590 1249.120 ;
        RECT 2540.190 1249.060 2540.510 1249.120 ;
        RECT 2539.270 1248.920 2540.510 1249.060 ;
        RECT 2539.270 1248.860 2539.590 1248.920 ;
        RECT 2540.190 1248.860 2540.510 1248.920 ;
        RECT 2539.270 1152.500 2539.590 1152.560 ;
        RECT 2540.190 1152.500 2540.510 1152.560 ;
        RECT 2539.270 1152.360 2540.510 1152.500 ;
        RECT 2539.270 1152.300 2539.590 1152.360 ;
        RECT 2540.190 1152.300 2540.510 1152.360 ;
        RECT 2539.270 1007.320 2539.590 1007.380 ;
        RECT 2540.190 1007.320 2540.510 1007.380 ;
        RECT 2539.270 1007.180 2540.510 1007.320 ;
        RECT 2539.270 1007.120 2539.590 1007.180 ;
        RECT 2540.190 1007.120 2540.510 1007.180 ;
        RECT 2539.270 910.760 2539.590 910.820 ;
        RECT 2540.190 910.760 2540.510 910.820 ;
        RECT 2539.270 910.620 2540.510 910.760 ;
        RECT 2539.270 910.560 2539.590 910.620 ;
        RECT 2540.190 910.560 2540.510 910.620 ;
        RECT 2539.270 814.200 2539.590 814.260 ;
        RECT 2539.075 814.060 2539.590 814.200 ;
        RECT 2539.270 814.000 2539.590 814.060 ;
        RECT 2539.270 766.260 2539.590 766.320 ;
        RECT 2539.075 766.120 2539.590 766.260 ;
        RECT 2539.270 766.060 2539.590 766.120 ;
        RECT 2539.270 717.640 2539.590 717.700 ;
        RECT 2539.075 717.500 2539.590 717.640 ;
        RECT 2539.270 717.440 2539.590 717.500 ;
        RECT 2539.270 669.700 2539.590 669.760 ;
        RECT 2539.075 669.560 2539.590 669.700 ;
        RECT 2539.270 669.500 2539.590 669.560 ;
        RECT 2539.270 620.740 2539.590 620.800 ;
        RECT 2539.075 620.600 2539.590 620.740 ;
        RECT 2539.270 620.540 2539.590 620.600 ;
        RECT 2539.270 572.800 2539.590 572.860 ;
        RECT 2539.075 572.660 2539.590 572.800 ;
        RECT 2539.270 572.600 2539.590 572.660 ;
        RECT 2539.270 524.180 2539.590 524.240 ;
        RECT 2539.075 524.040 2539.590 524.180 ;
        RECT 2539.270 523.980 2539.590 524.040 ;
        RECT 2539.270 476.240 2539.590 476.300 ;
        RECT 2539.075 476.100 2539.590 476.240 ;
        RECT 2539.270 476.040 2539.590 476.100 ;
        RECT 2539.270 427.620 2539.590 427.680 ;
        RECT 2539.075 427.480 2539.590 427.620 ;
        RECT 2539.270 427.420 2539.590 427.480 ;
        RECT 2539.270 379.680 2539.590 379.740 ;
        RECT 2539.075 379.540 2539.590 379.680 ;
        RECT 2539.270 379.480 2539.590 379.540 ;
        RECT 2539.270 331.060 2539.590 331.120 ;
        RECT 2539.075 330.920 2539.590 331.060 ;
        RECT 2539.270 330.860 2539.590 330.920 ;
        RECT 2539.270 283.120 2539.590 283.180 ;
        RECT 2539.075 282.980 2539.590 283.120 ;
        RECT 2539.270 282.920 2539.590 282.980 ;
        RECT 2539.270 234.500 2539.590 234.560 ;
        RECT 2539.075 234.360 2539.590 234.500 ;
        RECT 2539.270 234.300 2539.590 234.360 ;
        RECT 2539.270 186.560 2539.590 186.620 ;
        RECT 2539.075 186.420 2539.590 186.560 ;
        RECT 2539.270 186.360 2539.590 186.420 ;
        RECT 2539.270 137.940 2539.590 138.000 ;
        RECT 2539.075 137.800 2539.590 137.940 ;
        RECT 2539.270 137.740 2539.590 137.800 ;
        RECT 2539.270 90.000 2539.590 90.060 ;
        RECT 2539.075 89.860 2539.590 90.000 ;
        RECT 2539.270 89.800 2539.590 89.860 ;
        RECT 2539.270 62.120 2539.590 62.180 ;
        RECT 2542.030 62.120 2542.350 62.180 ;
        RECT 2539.270 61.980 2542.350 62.120 ;
        RECT 2539.270 61.920 2539.590 61.980 ;
        RECT 2542.030 61.920 2542.350 61.980 ;
      LAYER via ;
        RECT 1835.500 1683.720 1835.760 1683.980 ;
        RECT 1839.180 1683.720 1839.440 1683.980 ;
        RECT 1835.500 1645.640 1835.760 1645.900 ;
        RECT 2539.300 1635.440 2539.560 1635.700 ;
        RECT 2539.300 1586.820 2539.560 1587.080 ;
        RECT 2539.300 1538.880 2539.560 1539.140 ;
        RECT 2539.300 1490.260 2539.560 1490.520 ;
        RECT 2539.300 1441.980 2539.560 1442.240 ;
        RECT 2539.300 1345.420 2539.560 1345.680 ;
        RECT 2540.220 1345.420 2540.480 1345.680 ;
        RECT 2539.300 1248.860 2539.560 1249.120 ;
        RECT 2540.220 1248.860 2540.480 1249.120 ;
        RECT 2539.300 1152.300 2539.560 1152.560 ;
        RECT 2540.220 1152.300 2540.480 1152.560 ;
        RECT 2539.300 1007.120 2539.560 1007.380 ;
        RECT 2540.220 1007.120 2540.480 1007.380 ;
        RECT 2539.300 910.560 2539.560 910.820 ;
        RECT 2540.220 910.560 2540.480 910.820 ;
        RECT 2539.300 814.000 2539.560 814.260 ;
        RECT 2539.300 766.060 2539.560 766.320 ;
        RECT 2539.300 717.440 2539.560 717.700 ;
        RECT 2539.300 669.500 2539.560 669.760 ;
        RECT 2539.300 620.540 2539.560 620.800 ;
        RECT 2539.300 572.600 2539.560 572.860 ;
        RECT 2539.300 523.980 2539.560 524.240 ;
        RECT 2539.300 476.040 2539.560 476.300 ;
        RECT 2539.300 427.420 2539.560 427.680 ;
        RECT 2539.300 379.480 2539.560 379.740 ;
        RECT 2539.300 330.860 2539.560 331.120 ;
        RECT 2539.300 282.920 2539.560 283.180 ;
        RECT 2539.300 234.300 2539.560 234.560 ;
        RECT 2539.300 186.360 2539.560 186.620 ;
        RECT 2539.300 137.740 2539.560 138.000 ;
        RECT 2539.300 89.800 2539.560 90.060 ;
        RECT 2539.300 61.920 2539.560 62.180 ;
        RECT 2542.060 61.920 2542.320 62.180 ;
      LAYER met2 ;
        RECT 1839.170 1700.000 1839.450 1704.000 ;
        RECT 1839.240 1684.010 1839.380 1700.000 ;
        RECT 1835.500 1683.690 1835.760 1684.010 ;
        RECT 1839.180 1683.690 1839.440 1684.010 ;
        RECT 1835.560 1645.930 1835.700 1683.690 ;
        RECT 1835.500 1645.610 1835.760 1645.930 ;
        RECT 2539.300 1635.410 2539.560 1635.730 ;
        RECT 2539.360 1587.110 2539.500 1635.410 ;
        RECT 2539.300 1586.790 2539.560 1587.110 ;
        RECT 2539.300 1538.850 2539.560 1539.170 ;
        RECT 2539.360 1490.550 2539.500 1538.850 ;
        RECT 2539.300 1490.230 2539.560 1490.550 ;
        RECT 2539.300 1441.950 2539.560 1442.270 ;
        RECT 2539.360 1393.845 2539.500 1441.950 ;
        RECT 2539.290 1393.475 2539.570 1393.845 ;
        RECT 2540.210 1393.475 2540.490 1393.845 ;
        RECT 2540.280 1345.710 2540.420 1393.475 ;
        RECT 2539.300 1345.390 2539.560 1345.710 ;
        RECT 2540.220 1345.390 2540.480 1345.710 ;
        RECT 2539.360 1297.285 2539.500 1345.390 ;
        RECT 2539.290 1296.915 2539.570 1297.285 ;
        RECT 2540.210 1296.915 2540.490 1297.285 ;
        RECT 2540.280 1249.150 2540.420 1296.915 ;
        RECT 2539.300 1248.830 2539.560 1249.150 ;
        RECT 2540.220 1248.830 2540.480 1249.150 ;
        RECT 2539.360 1200.725 2539.500 1248.830 ;
        RECT 2539.290 1200.355 2539.570 1200.725 ;
        RECT 2540.210 1200.355 2540.490 1200.725 ;
        RECT 2540.280 1152.590 2540.420 1200.355 ;
        RECT 2539.300 1152.270 2539.560 1152.590 ;
        RECT 2540.220 1152.270 2540.480 1152.590 ;
        RECT 2539.360 1104.165 2539.500 1152.270 ;
        RECT 2539.290 1103.795 2539.570 1104.165 ;
        RECT 2540.210 1103.795 2540.490 1104.165 ;
        RECT 2540.280 1055.885 2540.420 1103.795 ;
        RECT 2539.290 1055.515 2539.570 1055.885 ;
        RECT 2540.210 1055.515 2540.490 1055.885 ;
        RECT 2539.360 1007.410 2539.500 1055.515 ;
        RECT 2539.300 1007.090 2539.560 1007.410 ;
        RECT 2540.220 1007.090 2540.480 1007.410 ;
        RECT 2540.280 959.325 2540.420 1007.090 ;
        RECT 2539.290 958.955 2539.570 959.325 ;
        RECT 2540.210 958.955 2540.490 959.325 ;
        RECT 2539.360 910.850 2539.500 958.955 ;
        RECT 2539.300 910.530 2539.560 910.850 ;
        RECT 2540.220 910.530 2540.480 910.850 ;
        RECT 2540.280 862.765 2540.420 910.530 ;
        RECT 2539.290 862.395 2539.570 862.765 ;
        RECT 2540.210 862.395 2540.490 862.765 ;
        RECT 2539.360 814.290 2539.500 862.395 ;
        RECT 2539.300 813.970 2539.560 814.290 ;
        RECT 2539.300 766.030 2539.560 766.350 ;
        RECT 2539.360 717.730 2539.500 766.030 ;
        RECT 2539.300 717.410 2539.560 717.730 ;
        RECT 2539.300 669.470 2539.560 669.790 ;
        RECT 2539.360 620.830 2539.500 669.470 ;
        RECT 2539.300 620.510 2539.560 620.830 ;
        RECT 2539.300 572.570 2539.560 572.890 ;
        RECT 2539.360 524.270 2539.500 572.570 ;
        RECT 2539.300 523.950 2539.560 524.270 ;
        RECT 2539.300 476.010 2539.560 476.330 ;
        RECT 2539.360 427.710 2539.500 476.010 ;
        RECT 2539.300 427.390 2539.560 427.710 ;
        RECT 2539.300 379.450 2539.560 379.770 ;
        RECT 2539.360 331.150 2539.500 379.450 ;
        RECT 2539.300 330.830 2539.560 331.150 ;
        RECT 2539.300 282.890 2539.560 283.210 ;
        RECT 2539.360 234.590 2539.500 282.890 ;
        RECT 2539.300 234.270 2539.560 234.590 ;
        RECT 2539.300 186.330 2539.560 186.650 ;
        RECT 2539.360 138.030 2539.500 186.330 ;
        RECT 2539.300 137.710 2539.560 138.030 ;
        RECT 2539.300 89.770 2539.560 90.090 ;
        RECT 2539.360 62.210 2539.500 89.770 ;
        RECT 2539.300 61.890 2539.560 62.210 ;
        RECT 2542.060 61.890 2542.320 62.210 ;
        RECT 2542.120 2.400 2542.260 61.890 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 2539.290 1393.520 2539.570 1393.800 ;
        RECT 2540.210 1393.520 2540.490 1393.800 ;
        RECT 2539.290 1296.960 2539.570 1297.240 ;
        RECT 2540.210 1296.960 2540.490 1297.240 ;
        RECT 2539.290 1200.400 2539.570 1200.680 ;
        RECT 2540.210 1200.400 2540.490 1200.680 ;
        RECT 2539.290 1103.840 2539.570 1104.120 ;
        RECT 2540.210 1103.840 2540.490 1104.120 ;
        RECT 2539.290 1055.560 2539.570 1055.840 ;
        RECT 2540.210 1055.560 2540.490 1055.840 ;
        RECT 2539.290 959.000 2539.570 959.280 ;
        RECT 2540.210 959.000 2540.490 959.280 ;
        RECT 2539.290 862.440 2539.570 862.720 ;
        RECT 2540.210 862.440 2540.490 862.720 ;
      LAYER met3 ;
        RECT 2539.265 1393.810 2539.595 1393.825 ;
        RECT 2540.185 1393.810 2540.515 1393.825 ;
        RECT 2539.265 1393.510 2540.515 1393.810 ;
        RECT 2539.265 1393.495 2539.595 1393.510 ;
        RECT 2540.185 1393.495 2540.515 1393.510 ;
        RECT 2539.265 1297.250 2539.595 1297.265 ;
        RECT 2540.185 1297.250 2540.515 1297.265 ;
        RECT 2539.265 1296.950 2540.515 1297.250 ;
        RECT 2539.265 1296.935 2539.595 1296.950 ;
        RECT 2540.185 1296.935 2540.515 1296.950 ;
        RECT 2539.265 1200.690 2539.595 1200.705 ;
        RECT 2540.185 1200.690 2540.515 1200.705 ;
        RECT 2539.265 1200.390 2540.515 1200.690 ;
        RECT 2539.265 1200.375 2539.595 1200.390 ;
        RECT 2540.185 1200.375 2540.515 1200.390 ;
        RECT 2539.265 1104.130 2539.595 1104.145 ;
        RECT 2540.185 1104.130 2540.515 1104.145 ;
        RECT 2539.265 1103.830 2540.515 1104.130 ;
        RECT 2539.265 1103.815 2539.595 1103.830 ;
        RECT 2540.185 1103.815 2540.515 1103.830 ;
        RECT 2539.265 1055.850 2539.595 1055.865 ;
        RECT 2540.185 1055.850 2540.515 1055.865 ;
        RECT 2539.265 1055.550 2540.515 1055.850 ;
        RECT 2539.265 1055.535 2539.595 1055.550 ;
        RECT 2540.185 1055.535 2540.515 1055.550 ;
        RECT 2539.265 959.290 2539.595 959.305 ;
        RECT 2540.185 959.290 2540.515 959.305 ;
        RECT 2539.265 958.990 2540.515 959.290 ;
        RECT 2539.265 958.975 2539.595 958.990 ;
        RECT 2540.185 958.975 2540.515 958.990 ;
        RECT 2539.265 862.730 2539.595 862.745 ;
        RECT 2540.185 862.730 2540.515 862.745 ;
        RECT 2539.265 862.430 2540.515 862.730 ;
        RECT 2539.265 862.415 2539.595 862.430 ;
        RECT 2540.185 862.415 2540.515 862.430 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1843.750 1684.260 1844.070 1684.320 ;
        RECT 1848.350 1684.260 1848.670 1684.320 ;
        RECT 1843.750 1684.120 1848.670 1684.260 ;
        RECT 1843.750 1684.060 1844.070 1684.120 ;
        RECT 1848.350 1684.060 1848.670 1684.120 ;
        RECT 1848.350 20.980 1848.670 21.040 ;
        RECT 2559.970 20.980 2560.290 21.040 ;
        RECT 1848.350 20.840 2560.290 20.980 ;
        RECT 1848.350 20.780 1848.670 20.840 ;
        RECT 2559.970 20.780 2560.290 20.840 ;
      LAYER via ;
        RECT 1843.780 1684.060 1844.040 1684.320 ;
        RECT 1848.380 1684.060 1848.640 1684.320 ;
        RECT 1848.380 20.780 1848.640 21.040 ;
        RECT 2560.000 20.780 2560.260 21.040 ;
      LAYER met2 ;
        RECT 1843.770 1700.000 1844.050 1704.000 ;
        RECT 1843.840 1684.350 1843.980 1700.000 ;
        RECT 1843.780 1684.030 1844.040 1684.350 ;
        RECT 1848.380 1684.030 1848.640 1684.350 ;
        RECT 1848.440 21.070 1848.580 1684.030 ;
        RECT 1848.380 20.750 1848.640 21.070 ;
        RECT 2560.000 20.750 2560.260 21.070 ;
        RECT 2560.060 2.400 2560.200 20.750 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1848.810 21.320 1849.130 21.380 ;
        RECT 2577.910 21.320 2578.230 21.380 ;
        RECT 1848.810 21.180 2578.230 21.320 ;
        RECT 1848.810 21.120 1849.130 21.180 ;
        RECT 2577.910 21.120 2578.230 21.180 ;
      LAYER via ;
        RECT 1848.840 21.120 1849.100 21.380 ;
        RECT 2577.940 21.120 2578.200 21.380 ;
      LAYER met2 ;
        RECT 1848.830 1700.000 1849.110 1704.000 ;
        RECT 1848.900 21.410 1849.040 1700.000 ;
        RECT 1848.840 21.090 1849.100 21.410 ;
        RECT 2577.940 21.090 2578.200 21.410 ;
        RECT 2578.000 2.400 2578.140 21.090 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 0.300 ;
=======
      LAYER met1 ;
        RECT 1359.830 1689.360 1360.150 1689.420 ;
        RECT 1369.490 1689.360 1369.810 1689.420 ;
        RECT 1359.830 1689.220 1369.810 1689.360 ;
        RECT 1359.830 1689.160 1360.150 1689.220 ;
        RECT 1369.490 1689.160 1369.810 1689.220 ;
        RECT 813.810 1673.380 814.130 1673.440 ;
        RECT 1359.830 1673.380 1360.150 1673.440 ;
        RECT 813.810 1673.240 1360.150 1673.380 ;
        RECT 813.810 1673.180 814.130 1673.240 ;
        RECT 1359.830 1673.180 1360.150 1673.240 ;
      LAYER via ;
        RECT 1359.860 1689.160 1360.120 1689.420 ;
        RECT 1369.520 1689.160 1369.780 1689.420 ;
        RECT 813.840 1673.180 814.100 1673.440 ;
        RECT 1359.860 1673.180 1360.120 1673.440 ;
      LAYER met2 ;
        RECT 1369.510 1700.000 1369.790 1704.000 ;
        RECT 1369.580 1689.450 1369.720 1700.000 ;
        RECT 1359.860 1689.130 1360.120 1689.450 ;
        RECT 1369.520 1689.130 1369.780 1689.450 ;
        RECT 1359.920 1673.470 1360.060 1689.130 ;
        RECT 813.840 1673.150 814.100 1673.470 ;
        RECT 1359.860 1673.150 1360.120 1673.470 ;
        RECT 813.900 3.130 814.040 1673.150 ;
        RECT 811.600 2.990 814.040 3.130 ;
        RECT 811.600 2.400 811.740 2.990 ;
        RECT 811.390 -4.800 811.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 0.300 ;
=======
      LAYER li1 ;
        RECT 1869.125 22.355 1869.295 22.695 ;
        RECT 1869.125 22.185 1870.675 22.355 ;
      LAYER mcon ;
        RECT 1869.125 22.525 1869.295 22.695 ;
        RECT 1870.505 22.185 1870.675 22.355 ;
      LAYER met1 ;
        RECT 1850.650 1685.620 1850.970 1685.680 ;
        RECT 1854.790 1685.620 1855.110 1685.680 ;
        RECT 1850.650 1685.480 1855.110 1685.620 ;
        RECT 1850.650 1685.420 1850.970 1685.480 ;
        RECT 1854.790 1685.420 1855.110 1685.480 ;
        RECT 1874.570 23.360 1874.890 23.420 ;
        RECT 2595.390 23.360 2595.710 23.420 ;
        RECT 1874.570 23.220 2595.710 23.360 ;
        RECT 1874.570 23.160 1874.890 23.220 ;
        RECT 2595.390 23.160 2595.710 23.220 ;
        RECT 1854.790 22.680 1855.110 22.740 ;
        RECT 1869.065 22.680 1869.355 22.725 ;
        RECT 1854.790 22.540 1869.355 22.680 ;
        RECT 1854.790 22.480 1855.110 22.540 ;
        RECT 1869.065 22.495 1869.355 22.540 ;
        RECT 1870.445 22.340 1870.735 22.385 ;
        RECT 1872.730 22.340 1873.050 22.400 ;
        RECT 1870.445 22.200 1873.050 22.340 ;
        RECT 1870.445 22.155 1870.735 22.200 ;
        RECT 1872.730 22.140 1873.050 22.200 ;
      LAYER via ;
        RECT 1850.680 1685.420 1850.940 1685.680 ;
        RECT 1854.820 1685.420 1855.080 1685.680 ;
        RECT 1874.600 23.160 1874.860 23.420 ;
        RECT 2595.420 23.160 2595.680 23.420 ;
        RECT 1854.820 22.480 1855.080 22.740 ;
        RECT 1872.760 22.140 1873.020 22.400 ;
      LAYER met2 ;
        RECT 1850.670 1700.000 1850.950 1704.000 ;
        RECT 1850.740 1685.710 1850.880 1700.000 ;
        RECT 1850.680 1685.390 1850.940 1685.710 ;
        RECT 1854.820 1685.390 1855.080 1685.710 ;
        RECT 1854.880 22.770 1855.020 1685.390 ;
        RECT 1874.600 23.130 1874.860 23.450 ;
        RECT 2595.420 23.130 2595.680 23.450 ;
        RECT 1874.660 22.850 1874.800 23.130 ;
        RECT 1854.820 22.450 1855.080 22.770 ;
        RECT 1872.820 22.710 1874.800 22.850 ;
        RECT 1872.820 22.430 1872.960 22.710 ;
        RECT 1872.760 22.110 1873.020 22.430 ;
        RECT 2595.480 2.400 2595.620 23.130 ;
=======
      LAYER met1 ;
        RECT 1853.410 1684.600 1853.730 1684.660 ;
        RECT 1855.710 1684.600 1856.030 1684.660 ;
        RECT 1853.410 1684.460 1856.030 1684.600 ;
        RECT 1853.410 1684.400 1853.730 1684.460 ;
        RECT 1855.710 1684.400 1856.030 1684.460 ;
        RECT 1855.710 21.660 1856.030 21.720 ;
        RECT 2595.390 21.660 2595.710 21.720 ;
        RECT 1855.710 21.520 2595.710 21.660 ;
        RECT 1855.710 21.460 1856.030 21.520 ;
        RECT 2595.390 21.460 2595.710 21.520 ;
      LAYER via ;
        RECT 1853.440 1684.400 1853.700 1684.660 ;
        RECT 1855.740 1684.400 1856.000 1684.660 ;
        RECT 1855.740 21.460 1856.000 21.720 ;
        RECT 2595.420 21.460 2595.680 21.720 ;
      LAYER met2 ;
        RECT 1853.430 1700.000 1853.710 1704.000 ;
        RECT 1853.500 1684.690 1853.640 1700.000 ;
        RECT 1853.440 1684.370 1853.700 1684.690 ;
        RECT 1855.740 1684.370 1856.000 1684.690 ;
        RECT 1855.800 21.750 1855.940 1684.370 ;
        RECT 1855.740 21.430 1856.000 21.750 ;
        RECT 2595.420 21.430 2595.680 21.750 ;
        RECT 2595.480 2.400 2595.620 21.430 ;
>>>>>>> re-updated local openlane
        RECT 2595.270 -4.800 2595.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1858.470 1684.600 1858.790 1684.660 ;
        RECT 1860.770 1684.600 1861.090 1684.660 ;
        RECT 1858.470 1684.460 1861.090 1684.600 ;
        RECT 1858.470 1684.400 1858.790 1684.460 ;
        RECT 1860.770 1684.400 1861.090 1684.460 ;
        RECT 1861.230 22.000 1861.550 22.060 ;
        RECT 2613.330 22.000 2613.650 22.060 ;
        RECT 1861.230 21.860 2613.650 22.000 ;
        RECT 1861.230 21.800 1861.550 21.860 ;
        RECT 2613.330 21.800 2613.650 21.860 ;
      LAYER via ;
        RECT 1858.500 1684.400 1858.760 1684.660 ;
        RECT 1860.800 1684.400 1861.060 1684.660 ;
        RECT 1861.260 21.800 1861.520 22.060 ;
        RECT 2613.360 21.800 2613.620 22.060 ;
      LAYER met2 ;
        RECT 1858.490 1700.000 1858.770 1704.000 ;
        RECT 1858.560 1684.690 1858.700 1700.000 ;
        RECT 1858.500 1684.370 1858.760 1684.690 ;
        RECT 1860.800 1684.370 1861.060 1684.690 ;
        RECT 1860.860 1656.210 1861.000 1684.370 ;
        RECT 1860.860 1656.070 1861.460 1656.210 ;
        RECT 1861.320 22.090 1861.460 1656.070 ;
        RECT 1861.260 21.770 1861.520 22.090 ;
        RECT 2613.360 21.770 2613.620 22.090 ;
        RECT 2613.420 2.400 2613.560 21.770 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 0.300 ;
=======
      LAYER li1 ;
        RECT 1880.625 27.285 1881.715 27.455 ;
        RECT 1880.625 26.945 1880.795 27.285 ;
      LAYER mcon ;
        RECT 1881.545 27.285 1881.715 27.455 ;
      LAYER met1 ;
        RECT 1860.310 1686.640 1860.630 1686.700 ;
        RECT 1862.610 1686.640 1862.930 1686.700 ;
        RECT 1860.310 1686.500 1862.930 1686.640 ;
        RECT 1860.310 1686.440 1860.630 1686.500 ;
        RECT 1862.610 1686.440 1862.930 1686.500 ;
        RECT 1881.485 27.440 1881.775 27.485 ;
        RECT 2631.270 27.440 2631.590 27.500 ;
        RECT 1881.485 27.300 2631.590 27.440 ;
        RECT 1881.485 27.255 1881.775 27.300 ;
        RECT 2631.270 27.240 2631.590 27.300 ;
        RECT 1880.565 27.100 1880.855 27.145 ;
        RECT 1873.740 26.960 1880.855 27.100 ;
        RECT 1862.610 26.760 1862.930 26.820 ;
        RECT 1873.740 26.760 1873.880 26.960 ;
        RECT 1880.565 26.915 1880.855 26.960 ;
        RECT 1862.610 26.620 1873.880 26.760 ;
        RECT 1862.610 26.560 1862.930 26.620 ;
      LAYER via ;
        RECT 1860.340 1686.440 1860.600 1686.700 ;
        RECT 1862.640 1686.440 1862.900 1686.700 ;
        RECT 2631.300 27.240 2631.560 27.500 ;
        RECT 1862.640 26.560 1862.900 26.820 ;
      LAYER met2 ;
        RECT 1860.330 1700.000 1860.610 1704.000 ;
        RECT 1860.400 1686.730 1860.540 1700.000 ;
        RECT 1860.340 1686.410 1860.600 1686.730 ;
        RECT 1862.640 1686.410 1862.900 1686.730 ;
        RECT 1862.700 26.850 1862.840 1686.410 ;
        RECT 2631.300 27.210 2631.560 27.530 ;
        RECT 1862.640 26.530 1862.900 26.850 ;
        RECT 2631.360 2.400 2631.500 27.210 ;
=======
      LAYER met1 ;
        RECT 1863.070 1684.940 1863.390 1685.000 ;
        RECT 1869.050 1684.940 1869.370 1685.000 ;
        RECT 1863.070 1684.800 1869.370 1684.940 ;
        RECT 1863.070 1684.740 1863.390 1684.800 ;
        RECT 1869.050 1684.740 1869.370 1684.800 ;
        RECT 1869.050 22.340 1869.370 22.400 ;
        RECT 2631.270 22.340 2631.590 22.400 ;
        RECT 1869.050 22.200 2631.590 22.340 ;
        RECT 1869.050 22.140 1869.370 22.200 ;
        RECT 2631.270 22.140 2631.590 22.200 ;
      LAYER via ;
        RECT 1863.100 1684.740 1863.360 1685.000 ;
        RECT 1869.080 1684.740 1869.340 1685.000 ;
        RECT 1869.080 22.140 1869.340 22.400 ;
        RECT 2631.300 22.140 2631.560 22.400 ;
      LAYER met2 ;
        RECT 1863.090 1700.000 1863.370 1704.000 ;
        RECT 1863.160 1685.030 1863.300 1700.000 ;
        RECT 1863.100 1684.710 1863.360 1685.030 ;
        RECT 1869.080 1684.710 1869.340 1685.030 ;
        RECT 1869.140 22.430 1869.280 1684.710 ;
        RECT 1869.080 22.110 1869.340 22.430 ;
        RECT 2631.300 22.110 2631.560 22.430 ;
        RECT 2631.360 2.400 2631.500 22.110 ;
>>>>>>> re-updated local openlane
        RECT 2631.150 -4.800 2631.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1868.130 1684.600 1868.450 1684.660 ;
        RECT 1869.510 1684.600 1869.830 1684.660 ;
        RECT 1868.130 1684.460 1869.830 1684.600 ;
        RECT 1868.130 1684.400 1868.450 1684.460 ;
        RECT 1869.510 1684.400 1869.830 1684.460 ;
        RECT 1869.510 22.680 1869.830 22.740 ;
        RECT 2649.210 22.680 2649.530 22.740 ;
        RECT 1869.510 22.540 2649.530 22.680 ;
        RECT 1869.510 22.480 1869.830 22.540 ;
        RECT 2649.210 22.480 2649.530 22.540 ;
      LAYER via ;
        RECT 1868.160 1684.400 1868.420 1684.660 ;
        RECT 1869.540 1684.400 1869.800 1684.660 ;
        RECT 1869.540 22.480 1869.800 22.740 ;
        RECT 2649.240 22.480 2649.500 22.740 ;
      LAYER met2 ;
        RECT 1868.150 1700.000 1868.430 1704.000 ;
        RECT 1868.220 1684.690 1868.360 1700.000 ;
        RECT 1868.160 1684.370 1868.420 1684.690 ;
        RECT 1869.540 1684.370 1869.800 1684.690 ;
        RECT 1869.600 22.770 1869.740 1684.370 ;
        RECT 1869.540 22.450 1869.800 22.770 ;
        RECT 2649.240 22.450 2649.500 22.770 ;
        RECT 2649.300 2.400 2649.440 22.450 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1872.730 1684.940 1873.050 1685.000 ;
        RECT 1876.410 1684.940 1876.730 1685.000 ;
        RECT 1872.730 1684.800 1876.730 1684.940 ;
        RECT 1872.730 1684.740 1873.050 1684.800 ;
        RECT 1876.410 1684.740 1876.730 1684.800 ;
        RECT 1876.410 23.020 1876.730 23.080 ;
        RECT 2667.150 23.020 2667.470 23.080 ;
        RECT 1876.410 22.880 2667.470 23.020 ;
        RECT 1876.410 22.820 1876.730 22.880 ;
        RECT 2667.150 22.820 2667.470 22.880 ;
      LAYER via ;
        RECT 1872.760 1684.740 1873.020 1685.000 ;
        RECT 1876.440 1684.740 1876.700 1685.000 ;
        RECT 1876.440 22.820 1876.700 23.080 ;
        RECT 2667.180 22.820 2667.440 23.080 ;
      LAYER met2 ;
        RECT 1872.750 1700.000 1873.030 1704.000 ;
        RECT 1872.820 1685.030 1872.960 1700.000 ;
        RECT 1872.760 1684.710 1873.020 1685.030 ;
        RECT 1876.440 1684.710 1876.700 1685.030 ;
        RECT 1876.500 23.110 1876.640 1684.710 ;
        RECT 1876.440 22.790 1876.700 23.110 ;
        RECT 2667.180 22.790 2667.440 23.110 ;
        RECT 2667.240 2.400 2667.380 22.790 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 0.300 ;
=======
      LAYER li1 ;
        RECT 1916.965 26.265 1918.055 26.435 ;
        RECT 1916.965 25.245 1917.135 26.265 ;
      LAYER mcon ;
        RECT 1917.885 26.265 1918.055 26.435 ;
      LAYER met1 ;
        RECT 1917.825 26.420 1918.115 26.465 ;
        RECT 2684.630 26.420 2684.950 26.480 ;
        RECT 1917.825 26.280 2684.950 26.420 ;
        RECT 1917.825 26.235 1918.115 26.280 ;
        RECT 2684.630 26.220 2684.950 26.280 ;
        RECT 1875.950 25.400 1876.270 25.460 ;
        RECT 1916.905 25.400 1917.195 25.445 ;
        RECT 1875.950 25.260 1917.195 25.400 ;
        RECT 1875.950 25.200 1876.270 25.260 ;
        RECT 1916.905 25.215 1917.195 25.260 ;
      LAYER via ;
        RECT 2684.660 26.220 2684.920 26.480 ;
        RECT 1875.980 25.200 1876.240 25.460 ;
      LAYER met2 ;
        RECT 1874.590 1700.410 1874.870 1704.000 ;
        RECT 1874.590 1700.270 1876.180 1700.410 ;
        RECT 1874.590 1700.000 1874.870 1700.270 ;
        RECT 1876.040 25.490 1876.180 1700.270 ;
        RECT 2684.660 26.190 2684.920 26.510 ;
        RECT 1875.980 25.170 1876.240 25.490 ;
        RECT 2684.720 2.400 2684.860 26.190 ;
=======
      LAYER met1 ;
        RECT 1877.790 1684.600 1878.110 1684.660 ;
        RECT 1883.310 1684.600 1883.630 1684.660 ;
        RECT 1877.790 1684.460 1883.630 1684.600 ;
        RECT 1877.790 1684.400 1878.110 1684.460 ;
        RECT 1883.310 1684.400 1883.630 1684.460 ;
        RECT 1883.310 23.360 1883.630 23.420 ;
        RECT 2684.630 23.360 2684.950 23.420 ;
        RECT 1883.310 23.220 2684.950 23.360 ;
        RECT 1883.310 23.160 1883.630 23.220 ;
        RECT 2684.630 23.160 2684.950 23.220 ;
      LAYER via ;
        RECT 1877.820 1684.400 1878.080 1684.660 ;
        RECT 1883.340 1684.400 1883.600 1684.660 ;
        RECT 1883.340 23.160 1883.600 23.420 ;
        RECT 2684.660 23.160 2684.920 23.420 ;
      LAYER met2 ;
        RECT 1877.810 1700.000 1878.090 1704.000 ;
        RECT 1877.880 1684.690 1878.020 1700.000 ;
        RECT 1877.820 1684.370 1878.080 1684.690 ;
        RECT 1883.340 1684.370 1883.600 1684.690 ;
        RECT 1883.400 23.450 1883.540 1684.370 ;
        RECT 1883.340 23.130 1883.600 23.450 ;
        RECT 2684.660 23.130 2684.920 23.450 ;
        RECT 2684.720 2.400 2684.860 23.130 ;
>>>>>>> re-updated local openlane
        RECT 2684.510 -4.800 2685.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1882.850 23.700 1883.170 23.760 ;
        RECT 2702.570 23.700 2702.890 23.760 ;
        RECT 1882.850 23.560 2702.890 23.700 ;
        RECT 1882.850 23.500 1883.170 23.560 ;
        RECT 2702.570 23.500 2702.890 23.560 ;
      LAYER via ;
        RECT 1882.880 23.500 1883.140 23.760 ;
        RECT 2702.600 23.500 2702.860 23.760 ;
      LAYER met2 ;
        RECT 1882.410 1700.410 1882.690 1704.000 ;
        RECT 1882.410 1700.270 1883.080 1700.410 ;
        RECT 1882.410 1700.000 1882.690 1700.270 ;
        RECT 1882.940 23.790 1883.080 1700.270 ;
        RECT 1882.880 23.470 1883.140 23.790 ;
        RECT 2702.600 23.470 2702.860 23.790 ;
        RECT 2702.660 2.400 2702.800 23.470 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 0.300 ;
=======
      LAYER li1 ;
        RECT 1916.505 25.075 1916.675 26.095 ;
        RECT 1917.425 25.585 1918.975 25.755 ;
        RECT 1917.425 25.075 1917.595 25.585 ;
        RECT 1916.505 24.905 1917.595 25.075 ;
      LAYER mcon ;
        RECT 1916.505 25.925 1916.675 26.095 ;
        RECT 1918.805 25.585 1918.975 25.755 ;
      LAYER met1 ;
        RECT 1884.230 1685.280 1884.550 1685.340 ;
        RECT 1890.210 1685.280 1890.530 1685.340 ;
        RECT 1884.230 1685.140 1890.530 1685.280 ;
        RECT 1884.230 1685.080 1884.550 1685.140 ;
        RECT 1890.210 1685.080 1890.530 1685.140 ;
        RECT 1890.210 26.080 1890.530 26.140 ;
        RECT 1916.445 26.080 1916.735 26.125 ;
        RECT 1890.210 25.940 1916.735 26.080 ;
        RECT 1890.210 25.880 1890.530 25.940 ;
        RECT 1916.445 25.895 1916.735 25.940 ;
        RECT 1918.745 25.740 1919.035 25.785 ;
        RECT 2720.510 25.740 2720.830 25.800 ;
        RECT 1918.745 25.600 2720.830 25.740 ;
        RECT 1918.745 25.555 1919.035 25.600 ;
        RECT 2720.510 25.540 2720.830 25.600 ;
      LAYER via ;
        RECT 1884.260 1685.080 1884.520 1685.340 ;
        RECT 1890.240 1685.080 1890.500 1685.340 ;
        RECT 1890.240 25.880 1890.500 26.140 ;
        RECT 2720.540 25.540 2720.800 25.800 ;
=======
      LAYER met1 ;
        RECT 1887.450 1683.920 1887.770 1683.980 ;
        RECT 1889.750 1683.920 1890.070 1683.980 ;
        RECT 1887.450 1683.780 1890.070 1683.920 ;
        RECT 1887.450 1683.720 1887.770 1683.780 ;
        RECT 1889.750 1683.720 1890.070 1683.780 ;
        RECT 1889.750 27.440 1890.070 27.500 ;
        RECT 2720.510 27.440 2720.830 27.500 ;
        RECT 1889.750 27.300 2720.830 27.440 ;
        RECT 1889.750 27.240 1890.070 27.300 ;
        RECT 2720.510 27.240 2720.830 27.300 ;
      LAYER via ;
        RECT 1887.480 1683.720 1887.740 1683.980 ;
        RECT 1889.780 1683.720 1890.040 1683.980 ;
        RECT 1889.780 27.240 1890.040 27.500 ;
        RECT 2720.540 27.240 2720.800 27.500 ;
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1887.470 1700.000 1887.750 1704.000 ;
        RECT 1887.540 1684.010 1887.680 1700.000 ;
        RECT 1887.480 1683.690 1887.740 1684.010 ;
        RECT 1889.780 1683.690 1890.040 1684.010 ;
        RECT 1889.840 27.530 1889.980 1683.690 ;
        RECT 1889.780 27.210 1890.040 27.530 ;
        RECT 2720.540 27.210 2720.800 27.530 ;
        RECT 2720.600 2.400 2720.740 27.210 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 0.300 ;
=======
      LAYER met1 ;
        RECT 1892.050 1684.600 1892.370 1684.660 ;
        RECT 1895.730 1684.600 1896.050 1684.660 ;
        RECT 1892.050 1684.460 1896.050 1684.600 ;
        RECT 1892.050 1684.400 1892.370 1684.460 ;
        RECT 1895.730 1684.400 1896.050 1684.460 ;
        RECT 1895.730 27.100 1896.050 27.160 ;
        RECT 2738.450 27.100 2738.770 27.160 ;
        RECT 1895.730 26.960 2738.770 27.100 ;
        RECT 1895.730 26.900 1896.050 26.960 ;
        RECT 2738.450 26.900 2738.770 26.960 ;
      LAYER via ;
        RECT 1892.080 1684.400 1892.340 1684.660 ;
        RECT 1895.760 1684.400 1896.020 1684.660 ;
        RECT 1895.760 26.900 1896.020 27.160 ;
        RECT 2738.480 26.900 2738.740 27.160 ;
      LAYER met2 ;
        RECT 1892.070 1700.000 1892.350 1704.000 ;
        RECT 1892.140 1684.690 1892.280 1700.000 ;
        RECT 1892.080 1684.370 1892.340 1684.690 ;
        RECT 1895.760 1684.370 1896.020 1684.690 ;
        RECT 1895.820 27.190 1895.960 1684.370 ;
        RECT 1895.760 26.870 1896.020 27.190 ;
        RECT 2738.480 26.870 2738.740 27.190 ;
        RECT 2738.540 2.400 2738.680 26.870 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1889.770 26.720 1890.050 27.000 ;
        RECT 2738.470 26.720 2738.750 27.000 ;
      LAYER met3 ;
        RECT 1889.745 27.010 1890.075 27.025 ;
        RECT 2738.445 27.010 2738.775 27.025 ;
        RECT 1889.745 26.710 2738.775 27.010 ;
        RECT 1889.745 26.695 1890.075 26.710 ;
        RECT 2738.445 26.695 2738.775 26.710 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 0.300 ;
=======
      LAYER met1 ;
        RECT 1896.190 26.760 1896.510 26.820 ;
        RECT 2755.930 26.760 2756.250 26.820 ;
        RECT 1896.190 26.620 2756.250 26.760 ;
        RECT 1896.190 26.560 1896.510 26.620 ;
        RECT 2755.930 26.560 2756.250 26.620 ;
      LAYER via ;
        RECT 1896.220 26.560 1896.480 26.820 ;
        RECT 2755.960 26.560 2756.220 26.820 ;
      LAYER met2 ;
        RECT 1897.130 1700.410 1897.410 1704.000 ;
        RECT 1896.280 1700.270 1897.410 1700.410 ;
        RECT 1896.280 26.850 1896.420 1700.270 ;
        RECT 1897.130 1700.000 1897.410 1700.270 ;
        RECT 1896.220 26.530 1896.480 26.850 ;
        RECT 2755.960 26.530 2756.220 26.850 ;
        RECT 2756.020 2.400 2756.160 26.530 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1897.130 26.040 1897.410 26.320 ;
        RECT 2755.950 26.040 2756.230 26.320 ;
      LAYER met3 ;
        RECT 1897.105 26.330 1897.435 26.345 ;
        RECT 2755.925 26.330 2756.255 26.345 ;
        RECT 1897.105 26.030 2756.255 26.330 ;
        RECT 1897.105 26.015 1897.435 26.030 ;
        RECT 2755.925 26.015 2756.255 26.030 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 0.300 ;
=======
      LAYER met1 ;
        RECT 834.510 1666.580 834.830 1666.640 ;
        RECT 1374.550 1666.580 1374.870 1666.640 ;
        RECT 834.510 1666.440 1374.870 1666.580 ;
        RECT 834.510 1666.380 834.830 1666.440 ;
        RECT 1374.550 1666.380 1374.870 1666.440 ;
        RECT 829.450 2.960 829.770 3.020 ;
        RECT 834.510 2.960 834.830 3.020 ;
        RECT 829.450 2.820 834.830 2.960 ;
        RECT 829.450 2.760 829.770 2.820 ;
        RECT 834.510 2.760 834.830 2.820 ;
      LAYER via ;
        RECT 834.540 1666.380 834.800 1666.640 ;
        RECT 1374.580 1666.380 1374.840 1666.640 ;
        RECT 829.480 2.760 829.740 3.020 ;
        RECT 834.540 2.760 834.800 3.020 ;
      LAYER met2 ;
        RECT 1374.570 1700.000 1374.850 1704.000 ;
        RECT 1374.640 1666.670 1374.780 1700.000 ;
        RECT 834.540 1666.350 834.800 1666.670 ;
        RECT 1374.580 1666.350 1374.840 1666.670 ;
        RECT 834.600 3.050 834.740 1666.350 ;
        RECT 829.480 2.730 829.740 3.050 ;
        RECT 834.540 2.730 834.800 3.050 ;
        RECT 829.540 2.400 829.680 2.730 ;
        RECT 829.330 -4.800 829.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1901.710 1684.260 1902.030 1684.320 ;
        RECT 1903.550 1684.260 1903.870 1684.320 ;
        RECT 1901.710 1684.120 1903.870 1684.260 ;
        RECT 1901.710 1684.060 1902.030 1684.120 ;
        RECT 1903.550 1684.060 1903.870 1684.120 ;
        RECT 1903.550 26.420 1903.870 26.480 ;
        RECT 2773.870 26.420 2774.190 26.480 ;
        RECT 1903.550 26.280 2774.190 26.420 ;
        RECT 1903.550 26.220 1903.870 26.280 ;
        RECT 2773.870 26.220 2774.190 26.280 ;
      LAYER via ;
        RECT 1901.740 1684.060 1902.000 1684.320 ;
        RECT 1903.580 1684.060 1903.840 1684.320 ;
        RECT 1903.580 26.220 1903.840 26.480 ;
        RECT 2773.900 26.220 2774.160 26.480 ;
      LAYER met2 ;
        RECT 1901.730 1700.000 1902.010 1704.000 ;
        RECT 1901.800 1684.350 1901.940 1700.000 ;
        RECT 1901.740 1684.030 1902.000 1684.350 ;
        RECT 1903.580 1684.030 1903.840 1684.350 ;
        RECT 1903.640 26.510 1903.780 1684.030 ;
        RECT 1903.580 26.190 1903.840 26.510 ;
        RECT 2773.900 26.190 2774.160 26.510 ;
        RECT 2773.960 2.400 2774.100 26.190 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1906.770 1683.920 1907.090 1683.980 ;
        RECT 1909.990 1683.920 1910.310 1683.980 ;
        RECT 1906.770 1683.780 1910.310 1683.920 ;
        RECT 1906.770 1683.720 1907.090 1683.780 ;
        RECT 1909.990 1683.720 1910.310 1683.780 ;
        RECT 1909.990 26.080 1910.310 26.140 ;
        RECT 2791.810 26.080 2792.130 26.140 ;
        RECT 1909.990 25.940 2792.130 26.080 ;
        RECT 1909.990 25.880 1910.310 25.940 ;
        RECT 2791.810 25.880 2792.130 25.940 ;
      LAYER via ;
        RECT 1906.800 1683.720 1907.060 1683.980 ;
        RECT 1910.020 1683.720 1910.280 1683.980 ;
        RECT 1910.020 25.880 1910.280 26.140 ;
        RECT 2791.840 25.880 2792.100 26.140 ;
      LAYER met2 ;
        RECT 1906.790 1700.000 1907.070 1704.000 ;
        RECT 1906.860 1684.010 1907.000 1700.000 ;
        RECT 1906.800 1683.690 1907.060 1684.010 ;
        RECT 1910.020 1683.690 1910.280 1684.010 ;
        RECT 1910.080 26.170 1910.220 1683.690 ;
        RECT 1910.020 25.850 1910.280 26.170 ;
        RECT 2791.840 25.850 2792.100 26.170 ;
        RECT 2791.900 2.400 2792.040 25.850 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1903.570 25.360 1903.850 25.640 ;
        RECT 2791.830 25.360 2792.110 25.640 ;
      LAYER met3 ;
        RECT 1903.545 25.650 1903.875 25.665 ;
        RECT 2791.805 25.650 2792.135 25.665 ;
        RECT 1903.545 25.350 2792.135 25.650 ;
        RECT 1903.545 25.335 1903.875 25.350 ;
        RECT 2791.805 25.335 2792.135 25.350 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1911.370 1684.940 1911.690 1685.000 ;
        RECT 1916.890 1684.940 1917.210 1685.000 ;
        RECT 1911.370 1684.800 1917.210 1684.940 ;
        RECT 1911.370 1684.740 1911.690 1684.800 ;
        RECT 1916.890 1684.740 1917.210 1684.800 ;
        RECT 1916.890 25.740 1917.210 25.800 ;
        RECT 2809.750 25.740 2810.070 25.800 ;
        RECT 1916.890 25.600 2810.070 25.740 ;
        RECT 1916.890 25.540 1917.210 25.600 ;
        RECT 2809.750 25.540 2810.070 25.600 ;
      LAYER via ;
        RECT 1911.400 1684.740 1911.660 1685.000 ;
        RECT 1916.920 1684.740 1917.180 1685.000 ;
        RECT 1916.920 25.540 1917.180 25.800 ;
        RECT 2809.780 25.540 2810.040 25.800 ;
      LAYER met2 ;
        RECT 1911.390 1700.000 1911.670 1704.000 ;
        RECT 1911.460 1685.030 1911.600 1700.000 ;
        RECT 1911.400 1684.710 1911.660 1685.030 ;
        RECT 1916.920 1684.710 1917.180 1685.030 ;
        RECT 1916.980 25.830 1917.120 1684.710 ;
        RECT 1916.920 25.510 1917.180 25.830 ;
        RECT 2809.780 25.510 2810.040 25.830 ;
        RECT 2809.840 2.400 2809.980 25.510 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 0.300 ;
=======
      LAYER li1 ;
        RECT 1941.805 24.735 1941.975 25.415 ;
        RECT 1941.805 24.565 1943.815 24.735 ;
      LAYER mcon ;
        RECT 1941.805 25.245 1941.975 25.415 ;
        RECT 1943.645 24.565 1943.815 24.735 ;
      LAYER met1 ;
        RECT 1913.210 1685.620 1913.530 1685.680 ;
        RECT 1917.810 1685.620 1918.130 1685.680 ;
        RECT 1913.210 1685.480 1918.130 1685.620 ;
        RECT 1913.210 1685.420 1913.530 1685.480 ;
        RECT 1917.810 1685.420 1918.130 1685.480 ;
        RECT 1917.810 25.400 1918.130 25.460 ;
        RECT 1941.745 25.400 1942.035 25.445 ;
        RECT 1917.810 25.260 1942.035 25.400 ;
        RECT 1917.810 25.200 1918.130 25.260 ;
        RECT 1941.745 25.215 1942.035 25.260 ;
        RECT 1943.585 24.720 1943.875 24.765 ;
        RECT 2827.690 24.720 2828.010 24.780 ;
        RECT 1943.585 24.580 2828.010 24.720 ;
        RECT 1943.585 24.535 1943.875 24.580 ;
        RECT 2827.690 24.520 2828.010 24.580 ;
      LAYER via ;
        RECT 1913.240 1685.420 1913.500 1685.680 ;
        RECT 1917.840 1685.420 1918.100 1685.680 ;
        RECT 1917.840 25.200 1918.100 25.460 ;
        RECT 2827.720 24.520 2827.980 24.780 ;
=======
      LAYER met1 ;
        RECT 1917.350 25.400 1917.670 25.460 ;
        RECT 2827.690 25.400 2828.010 25.460 ;
        RECT 1917.350 25.260 2828.010 25.400 ;
        RECT 1917.350 25.200 1917.670 25.260 ;
        RECT 2827.690 25.200 2828.010 25.260 ;
      LAYER via ;
        RECT 1917.380 25.200 1917.640 25.460 ;
        RECT 2827.720 25.200 2827.980 25.460 ;
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1916.450 1700.410 1916.730 1704.000 ;
        RECT 1916.450 1700.270 1917.580 1700.410 ;
        RECT 1916.450 1700.000 1916.730 1700.270 ;
        RECT 1917.440 25.490 1917.580 1700.270 ;
        RECT 1917.380 25.170 1917.640 25.490 ;
        RECT 2827.720 25.170 2827.980 25.490 ;
        RECT 2827.780 2.400 2827.920 25.170 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 0.300 ;
=======
      LAYER li1 ;
        RECT 1935.825 23.885 1935.995 24.735 ;
        RECT 1941.345 24.395 1941.515 24.735 ;
        RECT 1941.345 24.225 1943.355 24.395 ;
      LAYER mcon ;
        RECT 1935.825 24.565 1935.995 24.735 ;
        RECT 1941.345 24.565 1941.515 24.735 ;
        RECT 1943.185 24.225 1943.355 24.395 ;
      LAYER met1 ;
        RECT 1918.270 1686.300 1918.590 1686.360 ;
        RECT 1924.250 1686.300 1924.570 1686.360 ;
        RECT 1918.270 1686.160 1924.570 1686.300 ;
        RECT 1918.270 1686.100 1918.590 1686.160 ;
        RECT 1924.250 1686.100 1924.570 1686.160 ;
        RECT 1935.765 24.720 1936.055 24.765 ;
        RECT 1941.285 24.720 1941.575 24.765 ;
        RECT 1935.765 24.580 1941.575 24.720 ;
        RECT 1935.765 24.535 1936.055 24.580 ;
        RECT 1941.285 24.535 1941.575 24.580 ;
        RECT 1943.125 24.380 1943.415 24.425 ;
        RECT 2845.170 24.380 2845.490 24.440 ;
        RECT 1943.125 24.240 2845.490 24.380 ;
        RECT 1943.125 24.195 1943.415 24.240 ;
        RECT 2845.170 24.180 2845.490 24.240 ;
        RECT 1924.250 24.040 1924.570 24.100 ;
        RECT 1935.765 24.040 1936.055 24.085 ;
        RECT 1924.250 23.900 1936.055 24.040 ;
        RECT 1924.250 23.840 1924.570 23.900 ;
        RECT 1935.765 23.855 1936.055 23.900 ;
      LAYER via ;
        RECT 1918.300 1686.100 1918.560 1686.360 ;
        RECT 1924.280 1686.100 1924.540 1686.360 ;
        RECT 2845.200 24.180 2845.460 24.440 ;
        RECT 1924.280 23.840 1924.540 24.100 ;
      LAYER met2 ;
        RECT 1918.290 1700.000 1918.570 1704.000 ;
        RECT 1918.360 1686.390 1918.500 1700.000 ;
        RECT 1918.300 1686.070 1918.560 1686.390 ;
        RECT 1924.280 1686.070 1924.540 1686.390 ;
        RECT 1924.340 24.130 1924.480 1686.070 ;
        RECT 2845.200 24.150 2845.460 24.470 ;
        RECT 1924.280 23.810 1924.540 24.130 ;
        RECT 2845.260 2.400 2845.400 24.150 ;
=======
      LAYER met1 ;
        RECT 1921.030 1683.920 1921.350 1683.980 ;
        RECT 1923.790 1683.920 1924.110 1683.980 ;
        RECT 1921.030 1683.780 1924.110 1683.920 ;
        RECT 1921.030 1683.720 1921.350 1683.780 ;
        RECT 1923.790 1683.720 1924.110 1683.780 ;
        RECT 1923.790 25.060 1924.110 25.120 ;
        RECT 2845.170 25.060 2845.490 25.120 ;
        RECT 1923.790 24.920 2845.490 25.060 ;
        RECT 1923.790 24.860 1924.110 24.920 ;
        RECT 2845.170 24.860 2845.490 24.920 ;
      LAYER via ;
        RECT 1921.060 1683.720 1921.320 1683.980 ;
        RECT 1923.820 1683.720 1924.080 1683.980 ;
        RECT 1923.820 24.860 1924.080 25.120 ;
        RECT 2845.200 24.860 2845.460 25.120 ;
      LAYER met2 ;
        RECT 1921.050 1700.000 1921.330 1704.000 ;
        RECT 1921.120 1684.010 1921.260 1700.000 ;
        RECT 1921.060 1683.690 1921.320 1684.010 ;
        RECT 1923.820 1683.690 1924.080 1684.010 ;
        RECT 1923.880 25.150 1924.020 1683.690 ;
        RECT 1923.820 24.830 1924.080 25.150 ;
        RECT 2845.200 24.830 2845.460 25.150 ;
        RECT 2845.260 2.400 2845.400 24.830 ;
>>>>>>> re-updated local openlane
        RECT 2845.050 -4.800 2845.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1926.090 1684.260 1926.410 1684.320 ;
        RECT 1930.690 1684.260 1931.010 1684.320 ;
        RECT 1926.090 1684.120 1931.010 1684.260 ;
        RECT 1926.090 1684.060 1926.410 1684.120 ;
        RECT 1930.690 1684.060 1931.010 1684.120 ;
        RECT 1930.690 24.720 1931.010 24.780 ;
        RECT 2863.110 24.720 2863.430 24.780 ;
        RECT 1930.690 24.580 2863.430 24.720 ;
        RECT 1930.690 24.520 1931.010 24.580 ;
        RECT 2863.110 24.520 2863.430 24.580 ;
      LAYER via ;
        RECT 1926.120 1684.060 1926.380 1684.320 ;
        RECT 1930.720 1684.060 1930.980 1684.320 ;
        RECT 1930.720 24.520 1930.980 24.780 ;
        RECT 2863.140 24.520 2863.400 24.780 ;
      LAYER met2 ;
        RECT 1926.110 1700.000 1926.390 1704.000 ;
        RECT 1926.180 1684.350 1926.320 1700.000 ;
        RECT 1926.120 1684.030 1926.380 1684.350 ;
        RECT 1930.720 1684.030 1930.980 1684.350 ;
        RECT 1930.780 24.810 1930.920 1684.030 ;
        RECT 1930.720 24.490 1930.980 24.810 ;
        RECT 2863.140 24.490 2863.400 24.810 ;
        RECT 2863.200 2.400 2863.340 24.490 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1923.810 24.680 1924.090 24.960 ;
        RECT 2863.130 24.680 2863.410 24.960 ;
      LAYER met3 ;
        RECT 1923.785 24.970 1924.115 24.985 ;
        RECT 2863.105 24.970 2863.435 24.985 ;
        RECT 1923.785 24.670 2863.435 24.970 ;
        RECT 1923.785 24.655 1924.115 24.670 ;
        RECT 2863.105 24.655 2863.435 24.670 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1931.150 24.380 1931.470 24.440 ;
        RECT 2881.050 24.380 2881.370 24.440 ;
        RECT 1931.150 24.240 2881.370 24.380 ;
        RECT 1931.150 24.180 1931.470 24.240 ;
        RECT 2881.050 24.180 2881.370 24.240 ;
      LAYER via ;
        RECT 1931.180 24.180 1931.440 24.440 ;
        RECT 2881.080 24.180 2881.340 24.440 ;
      LAYER met2 ;
        RECT 1930.710 1700.410 1930.990 1704.000 ;
        RECT 1930.710 1700.270 1931.380 1700.410 ;
        RECT 1930.710 1700.000 1930.990 1700.270 ;
        RECT 1931.240 24.470 1931.380 1700.270 ;
        RECT 1931.180 24.150 1931.440 24.470 ;
        RECT 2881.080 24.150 2881.340 24.470 ;
        RECT 2881.140 2.400 2881.280 24.150 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1931.170 24.000 1931.450 24.280 ;
        RECT 2881.070 24.000 2881.350 24.280 ;
      LAYER met3 ;
        RECT 1931.145 24.290 1931.475 24.305 ;
        RECT 2881.045 24.290 2881.375 24.305 ;
        RECT 1931.145 23.990 2881.375 24.290 ;
        RECT 1931.145 23.975 1931.475 23.990 ;
        RECT 2881.045 23.975 2881.375 23.990 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1935.750 1683.920 1936.070 1683.980 ;
        RECT 1938.050 1683.920 1938.370 1683.980 ;
        RECT 1935.750 1683.780 1938.370 1683.920 ;
        RECT 1935.750 1683.720 1936.070 1683.780 ;
        RECT 1938.050 1683.720 1938.370 1683.780 ;
        RECT 1938.050 24.040 1938.370 24.100 ;
        RECT 2898.990 24.040 2899.310 24.100 ;
        RECT 1938.050 23.900 2899.310 24.040 ;
        RECT 1938.050 23.840 1938.370 23.900 ;
        RECT 2898.990 23.840 2899.310 23.900 ;
      LAYER via ;
        RECT 1935.780 1683.720 1936.040 1683.980 ;
        RECT 1938.080 1683.720 1938.340 1683.980 ;
        RECT 1938.080 23.840 1938.340 24.100 ;
        RECT 2899.020 23.840 2899.280 24.100 ;
      LAYER met2 ;
        RECT 1935.770 1700.000 1936.050 1704.000 ;
        RECT 1935.840 1684.010 1935.980 1700.000 ;
        RECT 1935.780 1683.690 1936.040 1684.010 ;
        RECT 1938.080 1683.690 1938.340 1684.010 ;
        RECT 1938.140 24.130 1938.280 1683.690 ;
        RECT 1938.080 23.810 1938.340 24.130 ;
        RECT 2899.020 23.810 2899.280 24.130 ;
        RECT 2899.080 2.400 2899.220 23.810 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 0.300 ;
=======
      LAYER met1 ;
        RECT 848.310 1659.780 848.630 1659.840 ;
        RECT 1379.150 1659.780 1379.470 1659.840 ;
        RECT 848.310 1659.640 1379.470 1659.780 ;
        RECT 848.310 1659.580 848.630 1659.640 ;
        RECT 1379.150 1659.580 1379.470 1659.640 ;
        RECT 846.930 2.960 847.250 3.020 ;
        RECT 848.310 2.960 848.630 3.020 ;
        RECT 846.930 2.820 848.630 2.960 ;
        RECT 846.930 2.760 847.250 2.820 ;
        RECT 848.310 2.760 848.630 2.820 ;
      LAYER via ;
        RECT 848.340 1659.580 848.600 1659.840 ;
        RECT 1379.180 1659.580 1379.440 1659.840 ;
        RECT 846.960 2.760 847.220 3.020 ;
        RECT 848.340 2.760 848.600 3.020 ;
      LAYER met2 ;
        RECT 1379.170 1700.000 1379.450 1704.000 ;
        RECT 1379.240 1659.870 1379.380 1700.000 ;
        RECT 848.340 1659.550 848.600 1659.870 ;
        RECT 1379.180 1659.550 1379.440 1659.870 ;
        RECT 848.400 3.050 848.540 1659.550 ;
        RECT 846.960 2.730 847.220 3.050 ;
        RECT 848.340 2.730 848.600 3.050 ;
        RECT 847.020 2.400 847.160 2.730 ;
        RECT 846.810 -4.800 847.370 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 846.950 26.040 847.230 26.320 ;
        RECT 1373.190 26.040 1373.470 26.320 ;
      LAYER met3 ;
        RECT 846.925 26.330 847.255 26.345 ;
        RECT 1373.165 26.330 1373.495 26.345 ;
        RECT 846.925 26.030 1373.495 26.330 ;
        RECT 846.925 26.015 847.255 26.030 ;
        RECT 1373.165 26.015 1373.495 26.030 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 864.750 -4.800 865.310 0.300 ;
=======
        RECT 1383.310 1700.410 1383.590 1704.000 ;
        RECT 1382.460 1700.270 1383.590 1700.410 ;
        RECT 1382.460 27.045 1382.600 1700.270 ;
        RECT 1383.310 1700.000 1383.590 1700.270 ;
        RECT 864.890 26.675 865.170 27.045 ;
        RECT 1382.390 26.675 1382.670 27.045 ;
        RECT 864.960 2.400 865.100 26.675 ;
        RECT 864.750 -4.800 865.310 2.400 ;
      LAYER via2 ;
        RECT 864.890 26.720 865.170 27.000 ;
        RECT 1382.390 26.720 1382.670 27.000 ;
      LAYER met3 ;
        RECT 864.865 27.010 865.195 27.025 ;
        RECT 1382.365 27.010 1382.695 27.025 ;
        RECT 864.865 26.710 1382.695 27.010 ;
        RECT 864.865 26.695 865.195 26.710 ;
        RECT 1382.365 26.695 1382.695 26.710 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1380.990 1678.140 1381.310 1678.200 ;
        RECT 1382.830 1678.140 1383.150 1678.200 ;
        RECT 1380.990 1678.000 1383.150 1678.140 ;
        RECT 1380.990 1677.940 1381.310 1678.000 ;
        RECT 1382.830 1677.940 1383.150 1678.000 ;
        RECT 869.010 1645.840 869.330 1645.900 ;
        RECT 1380.990 1645.840 1381.310 1645.900 ;
        RECT 869.010 1645.700 1381.310 1645.840 ;
        RECT 869.010 1645.640 869.330 1645.700 ;
        RECT 1380.990 1645.640 1381.310 1645.700 ;
        RECT 864.870 2.960 865.190 3.020 ;
        RECT 869.010 2.960 869.330 3.020 ;
        RECT 864.870 2.820 869.330 2.960 ;
        RECT 864.870 2.760 865.190 2.820 ;
        RECT 869.010 2.760 869.330 2.820 ;
      LAYER via ;
        RECT 1381.020 1677.940 1381.280 1678.200 ;
        RECT 1382.860 1677.940 1383.120 1678.200 ;
        RECT 869.040 1645.640 869.300 1645.900 ;
        RECT 1381.020 1645.640 1381.280 1645.900 ;
        RECT 864.900 2.760 865.160 3.020 ;
        RECT 869.040 2.760 869.300 3.020 ;
      LAYER met2 ;
        RECT 1384.230 1700.410 1384.510 1704.000 ;
        RECT 1382.920 1700.270 1384.510 1700.410 ;
        RECT 1382.920 1678.230 1383.060 1700.270 ;
        RECT 1384.230 1700.000 1384.510 1700.270 ;
        RECT 1381.020 1677.910 1381.280 1678.230 ;
        RECT 1382.860 1677.910 1383.120 1678.230 ;
        RECT 1381.080 1645.930 1381.220 1677.910 ;
        RECT 869.040 1645.610 869.300 1645.930 ;
        RECT 1381.020 1645.610 1381.280 1645.930 ;
        RECT 869.100 3.050 869.240 1645.610 ;
        RECT 864.900 2.730 865.160 3.050 ;
        RECT 869.040 2.730 869.300 3.050 ;
        RECT 864.960 2.400 865.100 2.730 ;
        RECT 864.750 -4.800 865.310 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 882.690 -4.800 883.250 0.300 ;
=======
        RECT 1387.910 1700.410 1388.190 1704.000 ;
        RECT 1387.060 1700.270 1388.190 1700.410 ;
        RECT 1387.060 27.725 1387.200 1700.270 ;
        RECT 1387.910 1700.000 1388.190 1700.270 ;
        RECT 882.830 27.355 883.110 27.725 ;
        RECT 1386.990 27.355 1387.270 27.725 ;
        RECT 882.900 2.400 883.040 27.355 ;
        RECT 882.690 -4.800 883.250 2.400 ;
      LAYER via2 ;
        RECT 882.830 27.400 883.110 27.680 ;
        RECT 1386.990 27.400 1387.270 27.680 ;
      LAYER met3 ;
        RECT 882.805 27.690 883.135 27.705 ;
        RECT 1386.965 27.690 1387.295 27.705 ;
        RECT 882.805 27.390 1387.295 27.690 ;
        RECT 882.805 27.375 883.135 27.390 ;
        RECT 1386.965 27.375 1387.295 27.390 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1386.510 1683.920 1386.830 1683.980 ;
        RECT 1388.810 1683.920 1389.130 1683.980 ;
        RECT 1386.510 1683.780 1389.130 1683.920 ;
        RECT 1386.510 1683.720 1386.830 1683.780 ;
        RECT 1388.810 1683.720 1389.130 1683.780 ;
        RECT 882.810 1652.980 883.130 1653.040 ;
        RECT 1386.510 1652.980 1386.830 1653.040 ;
        RECT 882.810 1652.840 1386.830 1652.980 ;
        RECT 882.810 1652.780 883.130 1652.840 ;
        RECT 1386.510 1652.780 1386.830 1652.840 ;
      LAYER via ;
        RECT 1386.540 1683.720 1386.800 1683.980 ;
        RECT 1388.840 1683.720 1389.100 1683.980 ;
        RECT 882.840 1652.780 883.100 1653.040 ;
        RECT 1386.540 1652.780 1386.800 1653.040 ;
      LAYER met2 ;
        RECT 1388.830 1700.000 1389.110 1704.000 ;
        RECT 1388.900 1684.010 1389.040 1700.000 ;
        RECT 1386.540 1683.690 1386.800 1684.010 ;
        RECT 1388.840 1683.690 1389.100 1684.010 ;
        RECT 1386.600 1653.070 1386.740 1683.690 ;
        RECT 882.840 1652.750 883.100 1653.070 ;
        RECT 1386.540 1652.750 1386.800 1653.070 ;
        RECT 882.900 2.400 883.040 1652.750 ;
        RECT 882.690 -4.800 883.250 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 0.300 ;
=======
      LAYER met1 ;
        RECT 903.510 1680.520 903.830 1680.580 ;
        RECT 1393.870 1680.520 1394.190 1680.580 ;
        RECT 903.510 1680.380 1394.190 1680.520 ;
        RECT 903.510 1680.320 903.830 1680.380 ;
        RECT 1393.870 1680.320 1394.190 1680.380 ;
        RECT 900.750 2.960 901.070 3.020 ;
        RECT 903.510 2.960 903.830 3.020 ;
        RECT 900.750 2.820 903.830 2.960 ;
        RECT 900.750 2.760 901.070 2.820 ;
        RECT 903.510 2.760 903.830 2.820 ;
      LAYER via ;
        RECT 903.540 1680.320 903.800 1680.580 ;
        RECT 1393.900 1680.320 1394.160 1680.580 ;
        RECT 900.780 2.760 901.040 3.020 ;
        RECT 903.540 2.760 903.800 3.020 ;
      LAYER met2 ;
        RECT 1393.890 1700.000 1394.170 1704.000 ;
        RECT 1393.960 1680.610 1394.100 1700.000 ;
        RECT 903.540 1680.290 903.800 1680.610 ;
        RECT 1393.900 1680.290 1394.160 1680.610 ;
        RECT 903.600 3.050 903.740 1680.290 ;
        RECT 900.780 2.730 901.040 3.050 ;
        RECT 903.540 2.730 903.800 3.050 ;
        RECT 900.840 2.400 900.980 2.730 ;
        RECT 900.630 -4.800 901.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 0.300 ;
=======
      LAYER met1 ;
        RECT 924.210 1632.240 924.530 1632.300 ;
        RECT 1396.630 1632.240 1396.950 1632.300 ;
        RECT 924.210 1632.100 1396.950 1632.240 ;
        RECT 924.210 1632.040 924.530 1632.100 ;
        RECT 1396.630 1632.040 1396.950 1632.100 ;
      LAYER via ;
        RECT 924.240 1632.040 924.500 1632.300 ;
        RECT 1396.660 1632.040 1396.920 1632.300 ;
      LAYER met2 ;
        RECT 1398.490 1700.410 1398.770 1704.000 ;
        RECT 1397.640 1700.270 1398.770 1700.410 ;
        RECT 1397.640 1678.140 1397.780 1700.270 ;
        RECT 1398.490 1700.000 1398.770 1700.270 ;
        RECT 1396.720 1678.000 1397.780 1678.140 ;
        RECT 1396.720 1632.330 1396.860 1678.000 ;
        RECT 924.240 1632.010 924.500 1632.330 ;
        RECT 1396.660 1632.010 1396.920 1632.330 ;
        RECT 924.300 58.890 924.440 1632.010 ;
        RECT 918.780 58.750 924.440 58.890 ;
        RECT 918.780 2.400 918.920 58.750 ;
        RECT 918.570 -4.800 919.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1400.770 1700.920 1401.090 1700.980 ;
        RECT 1402.150 1700.920 1402.470 1700.980 ;
        RECT 1400.770 1700.780 1402.470 1700.920 ;
        RECT 1400.770 1700.720 1401.090 1700.780 ;
        RECT 1402.150 1700.720 1402.470 1700.780 ;
      LAYER via ;
        RECT 1400.800 1700.720 1401.060 1700.980 ;
        RECT 1402.180 1700.720 1402.440 1700.980 ;
      LAYER met2 ;
        RECT 1403.550 1701.090 1403.830 1704.000 ;
        RECT 1402.240 1701.010 1403.830 1701.090 ;
        RECT 1400.800 1700.690 1401.060 1701.010 ;
        RECT 1402.180 1700.950 1403.830 1701.010 ;
        RECT 1402.180 1700.690 1402.440 1700.950 ;
        RECT 1400.860 24.325 1401.000 1700.690 ;
        RECT 1403.550 1700.000 1403.830 1700.950 ;
        RECT 936.190 23.955 936.470 24.325 ;
        RECT 1400.790 23.955 1401.070 24.325 ;
        RECT 936.260 2.400 936.400 23.955 ;
        RECT 936.050 -4.800 936.610 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 936.190 24.000 936.470 24.280 ;
        RECT 1400.790 24.000 1401.070 24.280 ;
      LAYER met3 ;
        RECT 936.165 24.290 936.495 24.305 ;
        RECT 1400.765 24.290 1401.095 24.305 ;
        RECT 936.165 23.990 1401.095 24.290 ;
        RECT 936.165 23.975 936.495 23.990 ;
        RECT 1400.765 23.975 1401.095 23.990 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 0.300 ;
=======
      LAYER li1 ;
        RECT 1403.605 1490.645 1403.775 1568.675 ;
        RECT 1404.065 1248.905 1404.235 1297.015 ;
        RECT 1403.145 1048.985 1403.315 1097.095 ;
        RECT 1403.145 993.565 1403.315 1041.675 ;
        RECT 1403.605 234.685 1403.775 255.935 ;
      LAYER mcon ;
        RECT 1403.605 1568.505 1403.775 1568.675 ;
        RECT 1404.065 1296.845 1404.235 1297.015 ;
        RECT 1403.145 1096.925 1403.315 1097.095 ;
        RECT 1403.145 1041.505 1403.315 1041.675 ;
        RECT 1403.605 255.765 1403.775 255.935 ;
      LAYER met1 ;
        RECT 1403.530 1686.640 1403.850 1686.700 ;
        RECT 1407.210 1686.640 1407.530 1686.700 ;
        RECT 1403.530 1686.500 1407.530 1686.640 ;
        RECT 1403.530 1686.440 1403.850 1686.500 ;
        RECT 1407.210 1686.440 1407.530 1686.500 ;
        RECT 1403.070 1593.820 1403.390 1593.880 ;
        RECT 1403.530 1593.820 1403.850 1593.880 ;
        RECT 1403.070 1593.680 1403.850 1593.820 ;
        RECT 1403.070 1593.620 1403.390 1593.680 ;
        RECT 1403.530 1593.620 1403.850 1593.680 ;
        RECT 1403.070 1568.660 1403.390 1568.720 ;
        RECT 1403.545 1568.660 1403.835 1568.705 ;
        RECT 1403.070 1568.520 1403.835 1568.660 ;
        RECT 1403.070 1568.460 1403.390 1568.520 ;
        RECT 1403.545 1568.475 1403.835 1568.520 ;
        RECT 1403.530 1490.800 1403.850 1490.860 ;
        RECT 1403.335 1490.660 1403.850 1490.800 ;
        RECT 1403.530 1490.600 1403.850 1490.660 ;
        RECT 1403.530 1463.060 1403.850 1463.320 ;
        RECT 1403.620 1462.640 1403.760 1463.060 ;
        RECT 1403.530 1462.380 1403.850 1462.640 ;
        RECT 1403.530 1327.600 1403.850 1327.660 ;
        RECT 1403.990 1327.600 1404.310 1327.660 ;
        RECT 1403.530 1327.460 1404.310 1327.600 ;
        RECT 1403.530 1327.400 1403.850 1327.460 ;
        RECT 1403.990 1327.400 1404.310 1327.460 ;
        RECT 1403.990 1297.000 1404.310 1297.060 ;
        RECT 1403.795 1296.860 1404.310 1297.000 ;
        RECT 1403.990 1296.800 1404.310 1296.860 ;
        RECT 1404.005 1249.060 1404.295 1249.105 ;
        RECT 1404.450 1249.060 1404.770 1249.120 ;
        RECT 1404.005 1248.920 1404.770 1249.060 ;
        RECT 1404.005 1248.875 1404.295 1248.920 ;
        RECT 1404.450 1248.860 1404.770 1248.920 ;
        RECT 1403.530 1159.100 1403.850 1159.360 ;
        RECT 1403.620 1158.680 1403.760 1159.100 ;
        RECT 1403.530 1158.420 1403.850 1158.680 ;
        RECT 1403.530 1135.300 1403.850 1135.560 ;
        RECT 1403.620 1134.880 1403.760 1135.300 ;
        RECT 1403.530 1134.620 1403.850 1134.880 ;
        RECT 1403.085 1097.080 1403.375 1097.125 ;
        RECT 1403.530 1097.080 1403.850 1097.140 ;
        RECT 1403.085 1096.940 1403.850 1097.080 ;
        RECT 1403.085 1096.895 1403.375 1096.940 ;
        RECT 1403.530 1096.880 1403.850 1096.940 ;
        RECT 1403.070 1049.140 1403.390 1049.200 ;
        RECT 1402.875 1049.000 1403.390 1049.140 ;
        RECT 1403.070 1048.940 1403.390 1049.000 ;
        RECT 1403.070 1041.660 1403.390 1041.720 ;
        RECT 1402.875 1041.520 1403.390 1041.660 ;
        RECT 1403.070 1041.460 1403.390 1041.520 ;
        RECT 1403.085 993.720 1403.375 993.765 ;
        RECT 1403.530 993.720 1403.850 993.780 ;
        RECT 1403.085 993.580 1403.850 993.720 ;
        RECT 1403.085 993.535 1403.375 993.580 ;
        RECT 1403.530 993.520 1403.850 993.580 ;
        RECT 1403.530 966.520 1403.850 966.580 ;
        RECT 1403.160 966.380 1403.850 966.520 ;
        RECT 1403.160 965.900 1403.300 966.380 ;
        RECT 1403.530 966.320 1403.850 966.380 ;
        RECT 1403.070 965.640 1403.390 965.900 ;
        RECT 1403.070 917.900 1403.390 917.960 ;
        RECT 1403.530 917.900 1403.850 917.960 ;
        RECT 1403.070 917.760 1403.850 917.900 ;
        RECT 1403.070 917.700 1403.390 917.760 ;
        RECT 1403.530 917.700 1403.850 917.760 ;
        RECT 1403.070 724.440 1403.390 724.500 ;
        RECT 1403.990 724.440 1404.310 724.500 ;
        RECT 1403.070 724.300 1404.310 724.440 ;
        RECT 1403.070 724.240 1403.390 724.300 ;
        RECT 1403.990 724.240 1404.310 724.300 ;
        RECT 1403.070 579.600 1403.390 579.660 ;
        RECT 1403.990 579.600 1404.310 579.660 ;
        RECT 1403.070 579.460 1404.310 579.600 ;
        RECT 1403.070 579.400 1403.390 579.460 ;
        RECT 1403.990 579.400 1404.310 579.460 ;
        RECT 1403.530 255.920 1403.850 255.980 ;
        RECT 1403.335 255.780 1403.850 255.920 ;
        RECT 1403.530 255.720 1403.850 255.780 ;
        RECT 1403.530 234.840 1403.850 234.900 ;
        RECT 1403.335 234.700 1403.850 234.840 ;
        RECT 1403.530 234.640 1403.850 234.700 ;
        RECT 1403.530 137.740 1403.850 138.000 ;
        RECT 1403.620 137.320 1403.760 137.740 ;
        RECT 1403.530 137.060 1403.850 137.320 ;
=======
      LAYER met1 ;
>>>>>>> re-updated local openlane
        RECT 954.110 27.100 954.430 27.160 ;
        RECT 1407.670 27.100 1407.990 27.160 ;
        RECT 954.110 26.960 1407.990 27.100 ;
        RECT 954.110 26.900 954.430 26.960 ;
        RECT 1407.670 26.900 1407.990 26.960 ;
      LAYER via ;
        RECT 954.140 26.900 954.400 27.160 ;
        RECT 1407.700 26.900 1407.960 27.160 ;
      LAYER met2 ;
        RECT 1408.150 1700.410 1408.430 1704.000 ;
        RECT 1407.760 1700.270 1408.430 1700.410 ;
        RECT 1407.760 27.190 1407.900 1700.270 ;
        RECT 1408.150 1700.000 1408.430 1700.270 ;
        RECT 954.140 26.870 954.400 27.190 ;
        RECT 1407.700 26.870 1407.960 27.190 ;
        RECT 954.200 2.400 954.340 26.870 ;
        RECT 953.990 -4.800 954.550 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1403.090 724.400 1403.370 724.680 ;
        RECT 1404.010 724.400 1404.290 724.680 ;
        RECT 1403.550 580.240 1403.830 580.520 ;
        RECT 1403.090 579.560 1403.370 579.840 ;
      LAYER met3 ;
        RECT 1403.065 724.690 1403.395 724.705 ;
        RECT 1403.985 724.690 1404.315 724.705 ;
        RECT 1403.065 724.390 1404.315 724.690 ;
        RECT 1403.065 724.375 1403.395 724.390 ;
        RECT 1403.985 724.375 1404.315 724.390 ;
        RECT 1403.525 580.530 1403.855 580.545 ;
        RECT 1402.390 580.230 1403.855 580.530 ;
        RECT 1402.390 579.850 1402.690 580.230 ;
        RECT 1403.525 580.215 1403.855 580.230 ;
        RECT 1403.065 579.850 1403.395 579.865 ;
        RECT 1402.390 579.550 1403.395 579.850 ;
        RECT 1403.065 579.535 1403.395 579.550 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1407.670 1678.480 1407.990 1678.540 ;
        RECT 1410.890 1678.480 1411.210 1678.540 ;
        RECT 1407.670 1678.340 1411.210 1678.480 ;
        RECT 1407.670 1678.280 1407.990 1678.340 ;
        RECT 1410.890 1678.280 1411.210 1678.340 ;
=======
      LAYER li1 ;
        RECT 1409.585 324.445 1409.755 372.215 ;
        RECT 1410.505 228.225 1410.675 275.995 ;
        RECT 1410.045 179.605 1410.215 227.715 ;
        RECT 1410.045 27.285 1410.215 41.395 ;
      LAYER mcon ;
        RECT 1409.585 372.045 1409.755 372.215 ;
        RECT 1410.505 275.825 1410.675 275.995 ;
        RECT 1410.045 227.545 1410.215 227.715 ;
        RECT 1410.045 41.225 1410.215 41.395 ;
      LAYER met1 ;
        RECT 1409.510 1580.220 1409.830 1580.280 ;
        RECT 1409.970 1580.220 1410.290 1580.280 ;
        RECT 1409.510 1580.080 1410.290 1580.220 ;
        RECT 1409.510 1580.020 1409.830 1580.080 ;
        RECT 1409.970 1580.020 1410.290 1580.080 ;
        RECT 1409.970 1497.400 1410.290 1497.660 ;
        RECT 1410.060 1496.920 1410.200 1497.400 ;
        RECT 1410.430 1496.920 1410.750 1496.980 ;
        RECT 1410.060 1496.780 1410.750 1496.920 ;
        RECT 1410.430 1496.720 1410.750 1496.780 ;
        RECT 1409.510 1435.380 1409.830 1435.440 ;
        RECT 1409.970 1435.380 1410.290 1435.440 ;
        RECT 1409.510 1435.240 1410.290 1435.380 ;
        RECT 1409.510 1435.180 1409.830 1435.240 ;
        RECT 1409.970 1435.180 1410.290 1435.240 ;
        RECT 1409.970 1290.540 1410.290 1290.600 ;
        RECT 1410.430 1290.540 1410.750 1290.600 ;
        RECT 1409.970 1290.400 1410.750 1290.540 ;
        RECT 1409.970 1290.340 1410.290 1290.400 ;
        RECT 1410.430 1290.340 1410.750 1290.400 ;
        RECT 1409.510 1256.200 1409.830 1256.260 ;
        RECT 1409.970 1256.200 1410.290 1256.260 ;
        RECT 1409.510 1256.060 1410.290 1256.200 ;
        RECT 1409.510 1256.000 1409.830 1256.060 ;
        RECT 1409.970 1256.000 1410.290 1256.060 ;
        RECT 1409.510 1097.080 1409.830 1097.140 ;
        RECT 1409.970 1097.080 1410.290 1097.140 ;
        RECT 1409.510 1096.940 1410.290 1097.080 ;
        RECT 1409.510 1096.880 1409.830 1096.940 ;
        RECT 1409.970 1096.880 1410.290 1096.940 ;
        RECT 1409.970 993.380 1410.290 993.440 ;
        RECT 1410.890 993.380 1411.210 993.440 ;
        RECT 1409.970 993.240 1411.210 993.380 ;
        RECT 1409.970 993.180 1410.290 993.240 ;
        RECT 1410.890 993.180 1411.210 993.240 ;
        RECT 1411.350 904.300 1411.670 904.360 ;
        RECT 1410.980 904.160 1411.670 904.300 ;
        RECT 1410.980 904.020 1411.120 904.160 ;
        RECT 1411.350 904.100 1411.670 904.160 ;
        RECT 1410.890 903.760 1411.210 904.020 ;
        RECT 1410.430 524.520 1410.750 524.580 ;
        RECT 1410.890 524.520 1411.210 524.580 ;
        RECT 1410.430 524.380 1411.210 524.520 ;
        RECT 1410.430 524.320 1410.750 524.380 ;
        RECT 1410.890 524.320 1411.210 524.380 ;
        RECT 1409.970 449.380 1410.290 449.440 ;
        RECT 1409.600 449.240 1410.290 449.380 ;
        RECT 1409.600 448.420 1409.740 449.240 ;
        RECT 1409.970 449.180 1410.290 449.240 ;
        RECT 1409.510 448.160 1409.830 448.420 ;
        RECT 1409.510 386.620 1409.830 386.880 ;
        RECT 1409.600 386.480 1409.740 386.620 ;
        RECT 1409.970 386.480 1410.290 386.540 ;
        RECT 1409.600 386.340 1410.290 386.480 ;
        RECT 1409.970 386.280 1410.290 386.340 ;
        RECT 1409.970 372.340 1410.290 372.600 ;
        RECT 1409.525 372.200 1409.815 372.245 ;
        RECT 1410.060 372.200 1410.200 372.340 ;
        RECT 1409.525 372.060 1410.200 372.200 ;
        RECT 1409.525 372.015 1409.815 372.060 ;
        RECT 1409.510 324.600 1409.830 324.660 ;
        RECT 1409.315 324.460 1409.830 324.600 ;
        RECT 1409.510 324.400 1409.830 324.460 ;
        RECT 1409.510 282.780 1409.830 282.840 ;
        RECT 1410.890 282.780 1411.210 282.840 ;
        RECT 1409.510 282.640 1411.210 282.780 ;
        RECT 1409.510 282.580 1409.830 282.640 ;
        RECT 1410.890 282.580 1411.210 282.640 ;
        RECT 1410.445 275.980 1410.735 276.025 ;
        RECT 1410.890 275.980 1411.210 276.040 ;
        RECT 1410.445 275.840 1411.210 275.980 ;
        RECT 1410.445 275.795 1410.735 275.840 ;
        RECT 1410.890 275.780 1411.210 275.840 ;
        RECT 1410.430 228.380 1410.750 228.440 ;
        RECT 1410.235 228.240 1410.750 228.380 ;
        RECT 1410.430 228.180 1410.750 228.240 ;
        RECT 1409.985 227.700 1410.275 227.745 ;
        RECT 1410.430 227.700 1410.750 227.760 ;
        RECT 1409.985 227.560 1410.750 227.700 ;
        RECT 1409.985 227.515 1410.275 227.560 ;
        RECT 1410.430 227.500 1410.750 227.560 ;
        RECT 1409.970 179.760 1410.290 179.820 ;
        RECT 1409.775 179.620 1410.290 179.760 ;
        RECT 1409.970 179.560 1410.290 179.620 ;
        RECT 1409.510 137.940 1409.830 138.000 ;
        RECT 1410.430 137.940 1410.750 138.000 ;
        RECT 1409.510 137.800 1410.750 137.940 ;
        RECT 1409.510 137.740 1409.830 137.800 ;
        RECT 1410.430 137.740 1410.750 137.800 ;
        RECT 1409.970 41.380 1410.290 41.440 ;
        RECT 1409.775 41.240 1410.290 41.380 ;
        RECT 1409.970 41.180 1410.290 41.240 ;
>>>>>>> re-updated local openlane
        RECT 972.050 27.440 972.370 27.500 ;
        RECT 1409.985 27.440 1410.275 27.485 ;
        RECT 972.050 27.300 1410.275 27.440 ;
        RECT 972.050 27.240 972.370 27.300 ;
        RECT 1409.985 27.255 1410.275 27.300 ;
      LAYER via ;
        RECT 1409.540 1580.020 1409.800 1580.280 ;
        RECT 1410.000 1580.020 1410.260 1580.280 ;
        RECT 1410.000 1497.400 1410.260 1497.660 ;
        RECT 1410.460 1496.720 1410.720 1496.980 ;
        RECT 1409.540 1435.180 1409.800 1435.440 ;
        RECT 1410.000 1435.180 1410.260 1435.440 ;
        RECT 1410.000 1290.340 1410.260 1290.600 ;
        RECT 1410.460 1290.340 1410.720 1290.600 ;
        RECT 1409.540 1256.000 1409.800 1256.260 ;
        RECT 1410.000 1256.000 1410.260 1256.260 ;
        RECT 1409.540 1096.880 1409.800 1097.140 ;
        RECT 1410.000 1096.880 1410.260 1097.140 ;
        RECT 1410.000 993.180 1410.260 993.440 ;
        RECT 1410.920 993.180 1411.180 993.440 ;
        RECT 1411.380 904.100 1411.640 904.360 ;
        RECT 1410.920 903.760 1411.180 904.020 ;
        RECT 1410.460 524.320 1410.720 524.580 ;
        RECT 1410.920 524.320 1411.180 524.580 ;
        RECT 1410.000 449.180 1410.260 449.440 ;
        RECT 1409.540 448.160 1409.800 448.420 ;
        RECT 1409.540 386.620 1409.800 386.880 ;
        RECT 1410.000 386.280 1410.260 386.540 ;
        RECT 1410.000 372.340 1410.260 372.600 ;
        RECT 1409.540 324.400 1409.800 324.660 ;
        RECT 1409.540 282.580 1409.800 282.840 ;
        RECT 1410.920 282.580 1411.180 282.840 ;
        RECT 1410.920 275.780 1411.180 276.040 ;
        RECT 1410.460 228.180 1410.720 228.440 ;
        RECT 1410.460 227.500 1410.720 227.760 ;
        RECT 1410.000 179.560 1410.260 179.820 ;
        RECT 1409.540 137.740 1409.800 138.000 ;
        RECT 1410.460 137.740 1410.720 138.000 ;
        RECT 1410.000 41.180 1410.260 41.440 ;
        RECT 972.080 27.240 972.340 27.500 ;
      LAYER met2 ;
        RECT 1413.210 1700.410 1413.490 1704.000 ;
        RECT 1411.900 1700.270 1413.490 1700.410 ;
        RECT 1411.900 1677.290 1412.040 1700.270 ;
        RECT 1413.210 1700.000 1413.490 1700.270 ;
        RECT 1409.600 1677.150 1412.040 1677.290 ;
        RECT 1409.600 1580.310 1409.740 1677.150 ;
        RECT 1409.540 1579.990 1409.800 1580.310 ;
        RECT 1410.000 1579.990 1410.260 1580.310 ;
        RECT 1410.060 1497.690 1410.200 1579.990 ;
        RECT 1410.000 1497.370 1410.260 1497.690 ;
        RECT 1410.460 1496.690 1410.720 1497.010 ;
        RECT 1410.520 1460.370 1410.660 1496.690 ;
        RECT 1410.060 1460.230 1410.660 1460.370 ;
        RECT 1410.060 1435.470 1410.200 1460.230 ;
        RECT 1409.540 1435.150 1409.800 1435.470 ;
        RECT 1410.000 1435.150 1410.260 1435.470 ;
        RECT 1409.600 1411.410 1409.740 1435.150 ;
        RECT 1409.600 1411.270 1410.200 1411.410 ;
        RECT 1410.060 1338.650 1410.200 1411.270 ;
        RECT 1410.060 1338.510 1410.660 1338.650 ;
        RECT 1410.520 1290.630 1410.660 1338.510 ;
        RECT 1410.000 1290.310 1410.260 1290.630 ;
        RECT 1410.460 1290.310 1410.720 1290.630 ;
        RECT 1410.060 1256.290 1410.200 1290.310 ;
        RECT 1409.540 1255.970 1409.800 1256.290 ;
        RECT 1410.000 1255.970 1410.260 1256.290 ;
        RECT 1409.600 1217.610 1409.740 1255.970 ;
        RECT 1409.600 1217.470 1410.200 1217.610 ;
        RECT 1410.060 1097.170 1410.200 1217.470 ;
        RECT 1409.540 1096.850 1409.800 1097.170 ;
        RECT 1410.000 1096.850 1410.260 1097.170 ;
        RECT 1409.600 1014.405 1409.740 1096.850 ;
        RECT 1409.530 1014.035 1409.810 1014.405 ;
        RECT 1409.990 1013.355 1410.270 1013.725 ;
        RECT 1410.060 993.470 1410.200 1013.355 ;
        RECT 1410.000 993.150 1410.260 993.470 ;
        RECT 1410.920 993.150 1411.180 993.470 ;
        RECT 1410.980 968.730 1411.120 993.150 ;
        RECT 1410.980 968.590 1411.580 968.730 ;
        RECT 1411.440 904.390 1411.580 968.590 ;
        RECT 1411.380 904.070 1411.640 904.390 ;
        RECT 1410.920 903.730 1411.180 904.050 ;
        RECT 1410.980 751.810 1411.120 903.730 ;
        RECT 1410.520 751.670 1411.120 751.810 ;
        RECT 1410.520 596.770 1410.660 751.670 ;
        RECT 1410.520 596.630 1411.120 596.770 ;
        RECT 1410.980 524.610 1411.120 596.630 ;
        RECT 1410.460 524.290 1410.720 524.610 ;
        RECT 1410.920 524.290 1411.180 524.610 ;
        RECT 1410.520 499.530 1410.660 524.290 ;
        RECT 1410.060 499.390 1410.660 499.530 ;
        RECT 1410.060 449.470 1410.200 499.390 ;
        RECT 1410.000 449.150 1410.260 449.470 ;
        RECT 1409.540 448.130 1409.800 448.450 ;
        RECT 1409.600 386.910 1409.740 448.130 ;
        RECT 1409.540 386.590 1409.800 386.910 ;
        RECT 1410.000 386.250 1410.260 386.570 ;
        RECT 1410.060 372.630 1410.200 386.250 ;
        RECT 1410.000 372.310 1410.260 372.630 ;
        RECT 1409.540 324.370 1409.800 324.690 ;
        RECT 1409.600 282.870 1409.740 324.370 ;
        RECT 1409.540 282.550 1409.800 282.870 ;
        RECT 1410.920 282.550 1411.180 282.870 ;
        RECT 1410.980 276.070 1411.120 282.550 ;
        RECT 1410.920 275.750 1411.180 276.070 ;
        RECT 1410.460 228.150 1410.720 228.470 ;
        RECT 1410.520 227.790 1410.660 228.150 ;
        RECT 1410.460 227.470 1410.720 227.790 ;
        RECT 1410.000 179.530 1410.260 179.850 ;
        RECT 1410.060 162.250 1410.200 179.530 ;
        RECT 1409.600 162.110 1410.200 162.250 ;
        RECT 1409.600 138.030 1409.740 162.110 ;
        RECT 1409.540 137.710 1409.800 138.030 ;
        RECT 1410.460 137.710 1410.720 138.030 ;
        RECT 1410.520 107.170 1410.660 137.710 ;
        RECT 1409.600 107.030 1410.660 107.170 ;
        RECT 1409.600 89.490 1409.740 107.030 ;
        RECT 1409.600 89.350 1410.200 89.490 ;
        RECT 1410.060 41.470 1410.200 89.350 ;
        RECT 1410.000 41.150 1410.260 41.470 ;
        RECT 972.080 27.210 972.340 27.530 ;
        RECT 972.140 2.400 972.280 27.210 ;
        RECT 971.930 -4.800 972.490 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 1409.530 1014.080 1409.810 1014.360 ;
        RECT 1409.990 1013.400 1410.270 1013.680 ;
      LAYER met3 ;
        RECT 1409.505 1014.370 1409.835 1014.385 ;
        RECT 1409.505 1014.055 1410.050 1014.370 ;
        RECT 1409.750 1013.705 1410.050 1014.055 ;
        RECT 1409.750 1013.390 1410.295 1013.705 ;
        RECT 1409.965 1013.375 1410.295 1013.390 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 650.970 26.420 651.290 26.480 ;
        RECT 1325.330 26.420 1325.650 26.480 ;
        RECT 650.970 26.280 1325.650 26.420 ;
        RECT 650.970 26.220 651.290 26.280 ;
        RECT 1325.330 26.220 1325.650 26.280 ;
      LAYER via ;
        RECT 651.000 26.220 651.260 26.480 ;
        RECT 1325.360 26.220 1325.620 26.480 ;
      LAYER met2 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 650.850 -4.800 651.410 0.300 ;
=======
        RECT 1325.350 1700.410 1325.630 1704.000 ;
        RECT 1324.960 1700.270 1325.630 1700.410 ;
        RECT 1324.960 25.685 1325.100 1700.270 ;
        RECT 1325.350 1700.000 1325.630 1700.270 ;
        RECT 650.990 25.315 651.270 25.685 ;
        RECT 1324.890 25.315 1325.170 25.685 ;
        RECT 651.060 2.400 651.200 25.315 ;
        RECT 650.850 -4.800 651.410 2.400 ;
      LAYER via2 ;
        RECT 650.990 25.360 651.270 25.640 ;
        RECT 1324.890 25.360 1325.170 25.640 ;
      LAYER met3 ;
        RECT 650.965 25.650 651.295 25.665 ;
        RECT 1324.865 25.650 1325.195 25.665 ;
        RECT 650.965 25.350 1325.195 25.650 ;
        RECT 650.965 25.335 651.295 25.350 ;
        RECT 1324.865 25.335 1325.195 25.350 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1326.270 1700.410 1326.550 1704.000 ;
        RECT 1325.420 1700.270 1326.550 1700.410 ;
        RECT 1325.420 26.510 1325.560 1700.270 ;
        RECT 1326.270 1700.000 1326.550 1700.270 ;
        RECT 651.000 26.190 651.260 26.510 ;
        RECT 1325.360 26.190 1325.620 26.510 ;
        RECT 651.060 2.400 651.200 26.190 ;
        RECT 650.850 -4.800 651.410 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 0.300 ;
=======
      LAYER met1 ;
        RECT 989.990 23.700 990.310 23.760 ;
        RECT 1416.870 23.700 1417.190 23.760 ;
        RECT 989.990 23.560 1417.190 23.700 ;
        RECT 989.990 23.500 990.310 23.560 ;
        RECT 1416.870 23.500 1417.190 23.560 ;
      LAYER via ;
        RECT 990.020 23.500 990.280 23.760 ;
        RECT 1416.900 23.500 1417.160 23.760 ;
      LAYER met2 ;
        RECT 1418.270 1700.410 1418.550 1704.000 ;
        RECT 1416.960 1700.270 1418.550 1700.410 ;
        RECT 1416.960 23.790 1417.100 1700.270 ;
        RECT 1418.270 1700.000 1418.550 1700.270 ;
        RECT 990.020 23.470 990.280 23.790 ;
        RECT 1416.900 23.470 1417.160 23.790 ;
        RECT 990.080 2.400 990.220 23.470 ;
        RECT 989.870 -4.800 990.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1007.470 23.360 1007.790 23.420 ;
        RECT 1421.930 23.360 1422.250 23.420 ;
        RECT 1007.470 23.220 1422.250 23.360 ;
        RECT 1007.470 23.160 1007.790 23.220 ;
        RECT 1421.930 23.160 1422.250 23.220 ;
      LAYER via ;
        RECT 1007.500 23.160 1007.760 23.420 ;
        RECT 1421.960 23.160 1422.220 23.420 ;
      LAYER met2 ;
        RECT 1422.870 1700.410 1423.150 1704.000 ;
        RECT 1422.020 1700.270 1423.150 1700.410 ;
        RECT 1422.020 23.450 1422.160 1700.270 ;
        RECT 1422.870 1700.000 1423.150 1700.270 ;
        RECT 1007.500 23.130 1007.760 23.450 ;
        RECT 1421.960 23.130 1422.220 23.450 ;
        RECT 1007.560 2.400 1007.700 23.130 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1423.310 1659.100 1423.630 1659.160 ;
        RECT 1426.530 1659.100 1426.850 1659.160 ;
        RECT 1423.310 1658.960 1426.850 1659.100 ;
        RECT 1423.310 1658.900 1423.630 1658.960 ;
        RECT 1426.530 1658.900 1426.850 1658.960 ;
        RECT 1025.410 23.020 1025.730 23.080 ;
        RECT 1423.310 23.020 1423.630 23.080 ;
        RECT 1025.410 22.880 1423.630 23.020 ;
        RECT 1025.410 22.820 1025.730 22.880 ;
        RECT 1423.310 22.820 1423.630 22.880 ;
      LAYER via ;
        RECT 1423.340 1658.900 1423.600 1659.160 ;
        RECT 1426.560 1658.900 1426.820 1659.160 ;
        RECT 1025.440 22.820 1025.700 23.080 ;
        RECT 1423.340 22.820 1423.600 23.080 ;
      LAYER met2 ;
        RECT 1427.930 1700.410 1428.210 1704.000 ;
        RECT 1426.620 1700.270 1428.210 1700.410 ;
        RECT 1426.620 1659.190 1426.760 1700.270 ;
        RECT 1427.930 1700.000 1428.210 1700.270 ;
        RECT 1423.340 1658.870 1423.600 1659.190 ;
        RECT 1426.560 1658.870 1426.820 1659.190 ;
        RECT 1423.400 23.110 1423.540 1658.870 ;
        RECT 1025.440 22.790 1025.700 23.110 ;
        RECT 1423.340 22.790 1423.600 23.110 ;
        RECT 1025.500 2.400 1025.640 22.790 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 0.300 ;
=======
      LAYER met1 ;
        RECT 1043.350 22.680 1043.670 22.740 ;
        RECT 1429.750 22.680 1430.070 22.740 ;
        RECT 1043.350 22.540 1430.070 22.680 ;
        RECT 1043.350 22.480 1043.670 22.540 ;
        RECT 1429.750 22.480 1430.070 22.540 ;
      LAYER via ;
        RECT 1043.380 22.480 1043.640 22.740 ;
        RECT 1429.780 22.480 1430.040 22.740 ;
      LAYER met2 ;
        RECT 1432.530 1700.410 1432.810 1704.000 ;
        RECT 1431.680 1700.270 1432.810 1700.410 ;
        RECT 1431.680 1659.610 1431.820 1700.270 ;
        RECT 1432.530 1700.000 1432.810 1700.270 ;
        RECT 1429.840 1659.470 1431.820 1659.610 ;
        RECT 1429.840 22.770 1429.980 1659.470 ;
        RECT 1043.380 22.450 1043.640 22.770 ;
        RECT 1429.780 22.450 1430.040 22.770 ;
        RECT 1043.440 2.400 1043.580 22.450 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1061.290 22.340 1061.610 22.400 ;
        RECT 1436.650 22.340 1436.970 22.400 ;
        RECT 1061.290 22.200 1436.970 22.340 ;
        RECT 1061.290 22.140 1061.610 22.200 ;
        RECT 1436.650 22.140 1436.970 22.200 ;
      LAYER via ;
        RECT 1061.320 22.140 1061.580 22.400 ;
        RECT 1436.680 22.140 1436.940 22.400 ;
      LAYER met2 ;
        RECT 1437.590 1700.410 1437.870 1704.000 ;
        RECT 1436.740 1700.270 1437.870 1700.410 ;
        RECT 1436.740 22.430 1436.880 1700.270 ;
        RECT 1437.590 1700.000 1437.870 1700.270 ;
        RECT 1061.320 22.110 1061.580 22.430 ;
        RECT 1436.680 22.110 1436.940 22.430 ;
        RECT 1061.380 2.400 1061.520 22.110 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1442.170 1689.360 1442.490 1689.420 ;
        RECT 1444.470 1689.360 1444.790 1689.420 ;
        RECT 1442.170 1689.220 1444.790 1689.360 ;
        RECT 1442.170 1689.160 1442.490 1689.220 ;
        RECT 1444.470 1689.160 1444.790 1689.220 ;
        RECT 1079.230 22.000 1079.550 22.060 ;
        RECT 1444.470 22.000 1444.790 22.060 ;
        RECT 1079.230 21.860 1444.790 22.000 ;
        RECT 1079.230 21.800 1079.550 21.860 ;
        RECT 1444.470 21.800 1444.790 21.860 ;
      LAYER via ;
        RECT 1442.200 1689.160 1442.460 1689.420 ;
        RECT 1444.500 1689.160 1444.760 1689.420 ;
        RECT 1079.260 21.800 1079.520 22.060 ;
        RECT 1444.500 21.800 1444.760 22.060 ;
      LAYER met2 ;
        RECT 1442.190 1700.000 1442.470 1704.000 ;
        RECT 1442.260 1689.450 1442.400 1700.000 ;
        RECT 1442.200 1689.130 1442.460 1689.450 ;
        RECT 1444.500 1689.130 1444.760 1689.450 ;
        RECT 1444.560 22.090 1444.700 1689.130 ;
        RECT 1079.260 21.770 1079.520 22.090 ;
        RECT 1444.500 21.770 1444.760 22.090 ;
        RECT 1079.320 2.400 1079.460 21.770 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 0.300 ;
=======
      LAYER met1 ;
        RECT 1443.550 1674.060 1443.870 1674.120 ;
        RECT 1445.850 1674.060 1446.170 1674.120 ;
        RECT 1443.550 1673.920 1446.170 1674.060 ;
        RECT 1443.550 1673.860 1443.870 1673.920 ;
        RECT 1445.850 1673.860 1446.170 1673.920 ;
        RECT 1096.710 21.660 1097.030 21.720 ;
        RECT 1443.550 21.660 1443.870 21.720 ;
        RECT 1096.710 21.520 1443.870 21.660 ;
        RECT 1096.710 21.460 1097.030 21.520 ;
        RECT 1443.550 21.460 1443.870 21.520 ;
      LAYER via ;
        RECT 1443.580 1673.860 1443.840 1674.120 ;
        RECT 1445.880 1673.860 1446.140 1674.120 ;
        RECT 1096.740 21.460 1097.000 21.720 ;
        RECT 1443.580 21.460 1443.840 21.720 ;
      LAYER met2 ;
        RECT 1447.250 1700.410 1447.530 1704.000 ;
        RECT 1445.940 1700.270 1447.530 1700.410 ;
        RECT 1445.940 1674.150 1446.080 1700.270 ;
        RECT 1447.250 1700.000 1447.530 1700.270 ;
        RECT 1443.580 1673.830 1443.840 1674.150 ;
        RECT 1445.880 1673.830 1446.140 1674.150 ;
        RECT 1443.640 21.750 1443.780 1673.830 ;
        RECT 1096.740 21.430 1097.000 21.750 ;
        RECT 1443.580 21.430 1443.840 21.750 ;
        RECT 1096.800 2.400 1096.940 21.430 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1449.070 1678.140 1449.390 1678.200 ;
        RECT 1450.910 1678.140 1451.230 1678.200 ;
        RECT 1449.070 1678.000 1451.230 1678.140 ;
        RECT 1449.070 1677.940 1449.390 1678.000 ;
        RECT 1450.910 1677.940 1451.230 1678.000 ;
        RECT 1114.650 21.320 1114.970 21.380 ;
        RECT 1449.070 21.320 1449.390 21.380 ;
        RECT 1114.650 21.180 1449.390 21.320 ;
        RECT 1114.650 21.120 1114.970 21.180 ;
        RECT 1449.070 21.120 1449.390 21.180 ;
      LAYER via ;
        RECT 1449.100 1677.940 1449.360 1678.200 ;
        RECT 1450.940 1677.940 1451.200 1678.200 ;
        RECT 1114.680 21.120 1114.940 21.380 ;
        RECT 1449.100 21.120 1449.360 21.380 ;
      LAYER met2 ;
        RECT 1451.850 1700.410 1452.130 1704.000 ;
        RECT 1451.000 1700.270 1452.130 1700.410 ;
        RECT 1451.000 1678.230 1451.140 1700.270 ;
        RECT 1451.850 1700.000 1452.130 1700.270 ;
        RECT 1449.100 1677.910 1449.360 1678.230 ;
        RECT 1450.940 1677.910 1451.200 1678.230 ;
        RECT 1449.160 21.410 1449.300 1677.910 ;
        RECT 1114.680 21.090 1114.940 21.410 ;
        RECT 1449.100 21.090 1449.360 21.410 ;
        RECT 1114.740 2.400 1114.880 21.090 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 0.300 ;
=======
      LAYER li1 ;
        RECT 1451.445 964.665 1451.615 966.535 ;
      LAYER mcon ;
        RECT 1451.445 966.365 1451.615 966.535 ;
      LAYER met1 ;
        RECT 1451.370 1678.140 1451.690 1678.200 ;
        RECT 1454.130 1678.140 1454.450 1678.200 ;
        RECT 1451.370 1678.000 1454.450 1678.140 ;
        RECT 1451.370 1677.940 1451.690 1678.000 ;
        RECT 1454.130 1677.940 1454.450 1678.000 ;
        RECT 1451.370 1153.320 1451.690 1153.580 ;
        RECT 1451.460 1152.560 1451.600 1153.320 ;
        RECT 1451.370 1152.300 1451.690 1152.560 ;
        RECT 1451.370 966.520 1451.690 966.580 ;
        RECT 1451.175 966.380 1451.690 966.520 ;
        RECT 1451.370 966.320 1451.690 966.380 ;
        RECT 1451.370 964.820 1451.690 964.880 ;
        RECT 1451.175 964.680 1451.690 964.820 ;
        RECT 1451.370 964.620 1451.690 964.680 ;
=======
      LAYER met1 ;
>>>>>>> re-updated local openlane
        RECT 1132.590 20.980 1132.910 21.040 ;
        RECT 1455.970 20.980 1456.290 21.040 ;
        RECT 1132.590 20.840 1456.290 20.980 ;
        RECT 1132.590 20.780 1132.910 20.840 ;
        RECT 1455.970 20.780 1456.290 20.840 ;
      LAYER via ;
        RECT 1132.620 20.780 1132.880 21.040 ;
        RECT 1456.000 20.780 1456.260 21.040 ;
      LAYER met2 ;
        RECT 1456.910 1700.410 1457.190 1704.000 ;
        RECT 1456.060 1700.270 1457.190 1700.410 ;
        RECT 1456.060 21.070 1456.200 1700.270 ;
        RECT 1456.910 1700.000 1457.190 1700.270 ;
        RECT 1132.620 20.750 1132.880 21.070 ;
        RECT 1456.000 20.750 1456.260 21.070 ;
        RECT 1132.680 2.400 1132.820 20.750 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 0.300 ;
=======
      LAYER met1 ;
        RECT 1456.430 1678.140 1456.750 1678.200 ;
        RECT 1460.570 1678.140 1460.890 1678.200 ;
        RECT 1456.430 1678.000 1460.890 1678.140 ;
        RECT 1456.430 1677.940 1456.750 1678.000 ;
        RECT 1460.570 1677.940 1460.890 1678.000 ;
        RECT 1150.530 24.040 1150.850 24.100 ;
        RECT 1456.430 24.040 1456.750 24.100 ;
        RECT 1150.530 23.900 1456.750 24.040 ;
        RECT 1150.530 23.840 1150.850 23.900 ;
        RECT 1456.430 23.840 1456.750 23.900 ;
      LAYER via ;
        RECT 1456.460 1677.940 1456.720 1678.200 ;
        RECT 1460.600 1677.940 1460.860 1678.200 ;
        RECT 1150.560 23.840 1150.820 24.100 ;
        RECT 1456.460 23.840 1456.720 24.100 ;
      LAYER met2 ;
        RECT 1461.510 1700.410 1461.790 1704.000 ;
        RECT 1460.660 1700.270 1461.790 1700.410 ;
        RECT 1460.660 1678.230 1460.800 1700.270 ;
        RECT 1461.510 1700.000 1461.790 1700.270 ;
        RECT 1456.460 1677.910 1456.720 1678.230 ;
        RECT 1460.600 1677.910 1460.860 1678.230 ;
        RECT 1456.520 24.130 1456.660 1677.910 ;
        RECT 1150.560 23.810 1150.820 24.130 ;
        RECT 1456.460 23.810 1456.720 24.130 ;
        RECT 1150.620 2.400 1150.760 23.810 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 0.300 ;
=======
      LAYER li1 ;
        RECT 1326.785 1345.125 1326.955 1368.075 ;
        RECT 1326.785 642.345 1326.955 710.515 ;
        RECT 1327.245 559.045 1327.415 607.155 ;
        RECT 1327.705 475.745 1327.875 537.115 ;
      LAYER mcon ;
        RECT 1326.785 1367.905 1326.955 1368.075 ;
        RECT 1326.785 710.345 1326.955 710.515 ;
        RECT 1327.245 606.985 1327.415 607.155 ;
        RECT 1327.705 536.945 1327.875 537.115 ;
      LAYER met1 ;
        RECT 1326.710 1642.440 1327.030 1642.500 ;
        RECT 1329.470 1642.440 1329.790 1642.500 ;
        RECT 1326.710 1642.300 1329.790 1642.440 ;
        RECT 1326.710 1642.240 1327.030 1642.300 ;
        RECT 1329.470 1642.240 1329.790 1642.300 ;
        RECT 1326.710 1545.880 1327.030 1545.940 ;
        RECT 1327.170 1545.880 1327.490 1545.940 ;
        RECT 1326.710 1545.740 1327.490 1545.880 ;
        RECT 1326.710 1545.680 1327.030 1545.740 ;
        RECT 1327.170 1545.680 1327.490 1545.740 ;
        RECT 1327.630 1401.380 1327.950 1401.440 ;
        RECT 1326.800 1401.240 1327.950 1401.380 ;
        RECT 1326.800 1401.100 1326.940 1401.240 ;
        RECT 1327.630 1401.180 1327.950 1401.240 ;
        RECT 1326.710 1400.840 1327.030 1401.100 ;
        RECT 1326.710 1368.060 1327.030 1368.120 ;
        RECT 1326.515 1367.920 1327.030 1368.060 ;
        RECT 1326.710 1367.860 1327.030 1367.920 ;
        RECT 1326.725 1345.280 1327.015 1345.325 ;
        RECT 1327.630 1345.280 1327.950 1345.340 ;
        RECT 1326.725 1345.140 1327.950 1345.280 ;
        RECT 1326.725 1345.095 1327.015 1345.140 ;
        RECT 1327.630 1345.080 1327.950 1345.140 ;
        RECT 1327.170 1297.340 1327.490 1297.400 ;
        RECT 1327.630 1297.340 1327.950 1297.400 ;
        RECT 1327.170 1297.200 1327.950 1297.340 ;
        RECT 1327.170 1297.140 1327.490 1297.200 ;
        RECT 1327.630 1297.140 1327.950 1297.200 ;
        RECT 1326.710 1249.060 1327.030 1249.120 ;
        RECT 1327.170 1249.060 1327.490 1249.120 ;
        RECT 1326.710 1248.920 1327.490 1249.060 ;
        RECT 1326.710 1248.860 1327.030 1248.920 ;
        RECT 1327.170 1248.860 1327.490 1248.920 ;
        RECT 1327.170 814.540 1327.490 814.600 ;
        RECT 1326.800 814.400 1327.490 814.540 ;
        RECT 1326.800 814.260 1326.940 814.400 ;
        RECT 1327.170 814.340 1327.490 814.400 ;
        RECT 1326.710 814.000 1327.030 814.260 ;
        RECT 1326.710 710.500 1327.030 710.560 ;
        RECT 1326.515 710.360 1327.030 710.500 ;
        RECT 1326.710 710.300 1327.030 710.360 ;
        RECT 1326.725 642.500 1327.015 642.545 ;
        RECT 1327.170 642.500 1327.490 642.560 ;
        RECT 1326.725 642.360 1327.490 642.500 ;
        RECT 1326.725 642.315 1327.015 642.360 ;
        RECT 1327.170 642.300 1327.490 642.360 ;
        RECT 1327.170 607.140 1327.490 607.200 ;
        RECT 1326.975 607.000 1327.490 607.140 ;
        RECT 1327.170 606.940 1327.490 607.000 ;
        RECT 1326.710 559.200 1327.030 559.260 ;
        RECT 1327.185 559.200 1327.475 559.245 ;
        RECT 1326.710 559.060 1327.475 559.200 ;
        RECT 1326.710 559.000 1327.030 559.060 ;
        RECT 1327.185 559.015 1327.475 559.060 ;
        RECT 1326.710 537.100 1327.030 537.160 ;
        RECT 1327.645 537.100 1327.935 537.145 ;
        RECT 1326.710 536.960 1327.935 537.100 ;
        RECT 1326.710 536.900 1327.030 536.960 ;
        RECT 1327.645 536.915 1327.935 536.960 ;
        RECT 1327.630 475.900 1327.950 475.960 ;
        RECT 1327.435 475.760 1327.950 475.900 ;
        RECT 1327.630 475.700 1327.950 475.760 ;
        RECT 1327.170 427.960 1327.490 428.020 ;
        RECT 1327.630 427.960 1327.950 428.020 ;
        RECT 1327.170 427.820 1327.950 427.960 ;
        RECT 1327.170 427.760 1327.490 427.820 ;
        RECT 1327.630 427.760 1327.950 427.820 ;
        RECT 1326.710 379.680 1327.030 379.740 ;
        RECT 1327.170 379.680 1327.490 379.740 ;
        RECT 1326.710 379.540 1327.490 379.680 ;
        RECT 1326.710 379.480 1327.030 379.540 ;
        RECT 1327.170 379.480 1327.490 379.540 ;
        RECT 1326.710 331.060 1327.030 331.120 ;
        RECT 1327.170 331.060 1327.490 331.120 ;
        RECT 1326.710 330.920 1327.490 331.060 ;
        RECT 1326.710 330.860 1327.030 330.920 ;
        RECT 1327.170 330.860 1327.490 330.920 ;
        RECT 1327.170 186.900 1327.490 186.960 ;
        RECT 1326.800 186.760 1327.490 186.900 ;
        RECT 1326.800 186.620 1326.940 186.760 ;
        RECT 1327.170 186.700 1327.490 186.760 ;
        RECT 1326.710 186.360 1327.030 186.620 ;
        RECT 1326.710 110.540 1327.030 110.800 ;
        RECT 1326.800 110.060 1326.940 110.540 ;
        RECT 1327.170 110.060 1327.490 110.120 ;
        RECT 1326.800 109.920 1327.490 110.060 ;
        RECT 1327.170 109.860 1327.490 109.920 ;
        RECT 668.910 25.740 669.230 25.800 ;
        RECT 1326.710 25.740 1327.030 25.800 ;
        RECT 668.910 25.600 1327.030 25.740 ;
        RECT 668.910 25.540 669.230 25.600 ;
        RECT 1326.710 25.540 1327.030 25.600 ;
      LAYER via ;
        RECT 1326.740 1642.240 1327.000 1642.500 ;
        RECT 1329.500 1642.240 1329.760 1642.500 ;
        RECT 1326.740 1545.680 1327.000 1545.940 ;
        RECT 1327.200 1545.680 1327.460 1545.940 ;
        RECT 1327.660 1401.180 1327.920 1401.440 ;
        RECT 1326.740 1400.840 1327.000 1401.100 ;
        RECT 1326.740 1367.860 1327.000 1368.120 ;
        RECT 1327.660 1345.080 1327.920 1345.340 ;
        RECT 1327.200 1297.140 1327.460 1297.400 ;
        RECT 1327.660 1297.140 1327.920 1297.400 ;
        RECT 1326.740 1248.860 1327.000 1249.120 ;
        RECT 1327.200 1248.860 1327.460 1249.120 ;
        RECT 1327.200 814.340 1327.460 814.600 ;
        RECT 1326.740 814.000 1327.000 814.260 ;
        RECT 1326.740 710.300 1327.000 710.560 ;
        RECT 1327.200 642.300 1327.460 642.560 ;
        RECT 1327.200 606.940 1327.460 607.200 ;
        RECT 1326.740 559.000 1327.000 559.260 ;
        RECT 1326.740 536.900 1327.000 537.160 ;
        RECT 1327.660 475.700 1327.920 475.960 ;
        RECT 1327.200 427.760 1327.460 428.020 ;
        RECT 1327.660 427.760 1327.920 428.020 ;
        RECT 1326.740 379.480 1327.000 379.740 ;
        RECT 1327.200 379.480 1327.460 379.740 ;
        RECT 1326.740 330.860 1327.000 331.120 ;
        RECT 1327.200 330.860 1327.460 331.120 ;
        RECT 1327.200 186.700 1327.460 186.960 ;
        RECT 1326.740 186.360 1327.000 186.620 ;
        RECT 1326.740 110.540 1327.000 110.800 ;
        RECT 1327.200 109.860 1327.460 110.120 ;
        RECT 668.940 25.540 669.200 25.800 ;
        RECT 1326.740 25.540 1327.000 25.800 ;
      LAYER met2 ;
        RECT 1330.410 1700.410 1330.690 1704.000 ;
        RECT 1329.560 1700.270 1330.690 1700.410 ;
        RECT 1329.560 1642.530 1329.700 1700.270 ;
        RECT 1330.410 1700.000 1330.690 1700.270 ;
        RECT 1326.740 1642.210 1327.000 1642.530 ;
        RECT 1329.500 1642.210 1329.760 1642.530 ;
        RECT 1326.800 1545.970 1326.940 1642.210 ;
        RECT 1326.740 1545.650 1327.000 1545.970 ;
        RECT 1327.200 1545.650 1327.460 1545.970 ;
        RECT 1327.260 1425.010 1327.400 1545.650 ;
        RECT 1327.260 1424.870 1327.860 1425.010 ;
        RECT 1327.720 1401.470 1327.860 1424.870 ;
        RECT 1327.660 1401.150 1327.920 1401.470 ;
        RECT 1326.740 1400.810 1327.000 1401.130 ;
        RECT 1326.800 1368.150 1326.940 1400.810 ;
        RECT 1326.740 1367.830 1327.000 1368.150 ;
        RECT 1327.660 1345.050 1327.920 1345.370 ;
        RECT 1327.720 1297.430 1327.860 1345.050 ;
        RECT 1327.200 1297.110 1327.460 1297.430 ;
        RECT 1327.660 1297.110 1327.920 1297.430 ;
        RECT 1327.260 1249.150 1327.400 1297.110 ;
        RECT 1326.740 1248.830 1327.000 1249.150 ;
        RECT 1327.200 1248.830 1327.460 1249.150 ;
        RECT 1326.800 1110.965 1326.940 1248.830 ;
        RECT 1326.730 1110.595 1327.010 1110.965 ;
        RECT 1327.190 1109.915 1327.470 1110.285 ;
        RECT 1327.260 814.630 1327.400 1109.915 ;
        RECT 1327.200 814.310 1327.460 814.630 ;
        RECT 1326.740 813.970 1327.000 814.290 ;
        RECT 1326.800 710.590 1326.940 813.970 ;
        RECT 1326.740 710.270 1327.000 710.590 ;
        RECT 1327.200 642.270 1327.460 642.590 ;
        RECT 1327.260 607.230 1327.400 642.270 ;
        RECT 1327.200 606.910 1327.460 607.230 ;
        RECT 1326.740 558.970 1327.000 559.290 ;
        RECT 1326.800 537.190 1326.940 558.970 ;
        RECT 1326.740 536.870 1327.000 537.190 ;
        RECT 1327.660 475.670 1327.920 475.990 ;
        RECT 1327.720 428.050 1327.860 475.670 ;
        RECT 1327.200 427.730 1327.460 428.050 ;
        RECT 1327.660 427.730 1327.920 428.050 ;
        RECT 1327.260 379.770 1327.400 427.730 ;
        RECT 1326.740 379.450 1327.000 379.770 ;
        RECT 1327.200 379.450 1327.460 379.770 ;
        RECT 1326.800 331.150 1326.940 379.450 ;
        RECT 1326.740 330.830 1327.000 331.150 ;
        RECT 1327.200 330.830 1327.460 331.150 ;
        RECT 1327.260 186.990 1327.400 330.830 ;
        RECT 1327.200 186.670 1327.460 186.990 ;
        RECT 1326.740 186.330 1327.000 186.650 ;
        RECT 1326.800 110.830 1326.940 186.330 ;
        RECT 1326.740 110.510 1327.000 110.830 ;
        RECT 1327.200 109.830 1327.460 110.150 ;
        RECT 1327.260 41.210 1327.400 109.830 ;
        RECT 1326.800 41.070 1327.400 41.210 ;
        RECT 1326.800 25.830 1326.940 41.070 ;
        RECT 668.940 25.510 669.200 25.830 ;
        RECT 1326.740 25.510 1327.000 25.830 ;
        RECT 669.000 2.400 669.140 25.510 ;
        RECT 668.790 -4.800 669.350 2.400 ;
      LAYER via2 ;
        RECT 1326.730 1110.640 1327.010 1110.920 ;
        RECT 1327.190 1109.960 1327.470 1110.240 ;
      LAYER met3 ;
        RECT 1326.705 1110.930 1327.035 1110.945 ;
        RECT 1326.705 1110.615 1327.250 1110.930 ;
        RECT 1326.950 1110.265 1327.250 1110.615 ;
        RECT 1326.950 1109.950 1327.495 1110.265 ;
        RECT 1327.165 1109.935 1327.495 1109.950 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1324.870 1678.140 1325.190 1678.200 ;
        RECT 1329.930 1678.140 1330.250 1678.200 ;
        RECT 1324.870 1678.000 1330.250 1678.140 ;
        RECT 1324.870 1677.940 1325.190 1678.000 ;
        RECT 1329.930 1677.940 1330.250 1678.000 ;
        RECT 668.910 26.760 669.230 26.820 ;
        RECT 1324.870 26.760 1325.190 26.820 ;
        RECT 668.910 26.620 1325.190 26.760 ;
        RECT 668.910 26.560 669.230 26.620 ;
        RECT 1324.870 26.560 1325.190 26.620 ;
      LAYER via ;
        RECT 1324.900 1677.940 1325.160 1678.200 ;
        RECT 1329.960 1677.940 1330.220 1678.200 ;
        RECT 668.940 26.560 669.200 26.820 ;
        RECT 1324.900 26.560 1325.160 26.820 ;
      LAYER met2 ;
        RECT 1330.870 1700.410 1331.150 1704.000 ;
        RECT 1330.020 1700.270 1331.150 1700.410 ;
        RECT 1330.020 1678.230 1330.160 1700.270 ;
        RECT 1330.870 1700.000 1331.150 1700.270 ;
        RECT 1324.900 1677.910 1325.160 1678.230 ;
        RECT 1329.960 1677.910 1330.220 1678.230 ;
        RECT 1324.960 26.850 1325.100 1677.910 ;
        RECT 668.940 26.530 669.200 26.850 ;
        RECT 1324.900 26.530 1325.160 26.850 ;
        RECT 669.000 2.400 669.140 26.530 ;
        RECT 668.790 -4.800 669.350 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1464.250 1692.760 1464.570 1692.820 ;
        RECT 1466.550 1692.760 1466.870 1692.820 ;
        RECT 1464.250 1692.620 1466.870 1692.760 ;
        RECT 1464.250 1692.560 1464.570 1692.620 ;
        RECT 1466.550 1692.560 1466.870 1692.620 ;
        RECT 1168.470 24.380 1168.790 24.440 ;
        RECT 1464.250 24.380 1464.570 24.440 ;
        RECT 1168.470 24.240 1464.570 24.380 ;
        RECT 1168.470 24.180 1168.790 24.240 ;
        RECT 1464.250 24.180 1464.570 24.240 ;
      LAYER via ;
        RECT 1464.280 1692.560 1464.540 1692.820 ;
        RECT 1466.580 1692.560 1466.840 1692.820 ;
        RECT 1168.500 24.180 1168.760 24.440 ;
        RECT 1464.280 24.180 1464.540 24.440 ;
      LAYER met2 ;
        RECT 1466.570 1700.000 1466.850 1704.000 ;
        RECT 1466.640 1692.850 1466.780 1700.000 ;
        RECT 1464.280 1692.530 1464.540 1692.850 ;
        RECT 1466.580 1692.530 1466.840 1692.850 ;
        RECT 1464.340 24.470 1464.480 1692.530 ;
        RECT 1168.500 24.150 1168.760 24.470 ;
        RECT 1464.280 24.150 1464.540 24.470 ;
        RECT 1168.560 2.400 1168.700 24.150 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1185.830 -4.800 1186.390 0.300 ;
=======
        RECT 1469.790 1700.000 1470.070 1704.000 ;
        RECT 1469.860 16.845 1470.000 1700.000 ;
        RECT 1185.970 16.475 1186.250 16.845 ;
        RECT 1469.790 16.475 1470.070 16.845 ;
        RECT 1186.040 2.400 1186.180 16.475 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
      LAYER via2 ;
        RECT 1185.970 16.520 1186.250 16.800 ;
        RECT 1469.790 16.520 1470.070 16.800 ;
      LAYER met3 ;
        RECT 1185.945 16.810 1186.275 16.825 ;
        RECT 1469.765 16.810 1470.095 16.825 ;
        RECT 1185.945 16.510 1470.095 16.810 ;
        RECT 1185.945 16.495 1186.275 16.510 ;
        RECT 1469.765 16.495 1470.095 16.510 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1472.145 1635.485 1472.315 1683.595 ;
      LAYER mcon ;
        RECT 1472.145 1683.425 1472.315 1683.595 ;
      LAYER met1 ;
        RECT 1472.070 1683.580 1472.390 1683.640 ;
        RECT 1471.875 1683.440 1472.390 1683.580 ;
        RECT 1472.070 1683.380 1472.390 1683.440 ;
        RECT 1472.085 1635.640 1472.375 1635.685 ;
        RECT 1472.530 1635.640 1472.850 1635.700 ;
        RECT 1472.085 1635.500 1472.850 1635.640 ;
        RECT 1472.085 1635.455 1472.375 1635.500 ;
        RECT 1472.530 1635.440 1472.850 1635.500 ;
        RECT 1472.070 1545.880 1472.390 1545.940 ;
        RECT 1472.530 1545.880 1472.850 1545.940 ;
        RECT 1472.070 1545.740 1472.850 1545.880 ;
        RECT 1472.070 1545.680 1472.390 1545.740 ;
        RECT 1472.530 1545.680 1472.850 1545.740 ;
        RECT 1472.070 1418.040 1472.390 1418.100 ;
        RECT 1472.990 1418.040 1473.310 1418.100 ;
        RECT 1472.070 1417.900 1473.310 1418.040 ;
        RECT 1472.070 1417.840 1472.390 1417.900 ;
        RECT 1472.990 1417.840 1473.310 1417.900 ;
        RECT 1471.150 1389.140 1471.470 1389.200 ;
        RECT 1472.070 1389.140 1472.390 1389.200 ;
        RECT 1471.150 1389.000 1472.390 1389.140 ;
        RECT 1471.150 1388.940 1471.470 1389.000 ;
        RECT 1472.070 1388.940 1472.390 1389.000 ;
        RECT 1471.150 1318.080 1471.470 1318.140 ;
        RECT 1472.070 1318.080 1472.390 1318.140 ;
        RECT 1471.150 1317.940 1472.390 1318.080 ;
        RECT 1471.150 1317.880 1471.470 1317.940 ;
        RECT 1472.070 1317.880 1472.390 1317.940 ;
        RECT 1472.070 1269.800 1472.390 1269.860 ;
        RECT 1472.990 1269.800 1473.310 1269.860 ;
        RECT 1472.070 1269.660 1473.310 1269.800 ;
        RECT 1472.070 1269.600 1472.390 1269.660 ;
        RECT 1472.990 1269.600 1473.310 1269.660 ;
        RECT 1472.070 1221.520 1472.390 1221.580 ;
        RECT 1472.990 1221.520 1473.310 1221.580 ;
        RECT 1472.070 1221.380 1473.310 1221.520 ;
        RECT 1472.070 1221.320 1472.390 1221.380 ;
        RECT 1472.990 1221.320 1473.310 1221.380 ;
        RECT 1471.150 1197.380 1471.470 1197.440 ;
        RECT 1472.070 1197.380 1472.390 1197.440 ;
        RECT 1471.150 1197.240 1472.390 1197.380 ;
        RECT 1471.150 1197.180 1471.470 1197.240 ;
        RECT 1472.070 1197.180 1472.390 1197.240 ;
        RECT 1471.150 1124.960 1471.470 1125.020 ;
        RECT 1472.070 1124.960 1472.390 1125.020 ;
        RECT 1471.150 1124.820 1472.390 1124.960 ;
        RECT 1471.150 1124.760 1471.470 1124.820 ;
        RECT 1472.070 1124.760 1472.390 1124.820 ;
        RECT 1472.070 1076.680 1472.390 1076.740 ;
        RECT 1472.990 1076.680 1473.310 1076.740 ;
        RECT 1472.070 1076.540 1473.310 1076.680 ;
        RECT 1472.070 1076.480 1472.390 1076.540 ;
        RECT 1472.990 1076.480 1473.310 1076.540 ;
        RECT 1472.070 1028.400 1472.390 1028.460 ;
        RECT 1472.990 1028.400 1473.310 1028.460 ;
        RECT 1472.070 1028.260 1473.310 1028.400 ;
        RECT 1472.070 1028.200 1472.390 1028.260 ;
        RECT 1472.990 1028.200 1473.310 1028.260 ;
        RECT 1471.150 979.780 1471.470 979.840 ;
        RECT 1472.070 979.780 1472.390 979.840 ;
        RECT 1471.150 979.640 1472.390 979.780 ;
        RECT 1471.150 979.580 1471.470 979.640 ;
        RECT 1472.070 979.580 1472.390 979.640 ;
        RECT 1471.150 931.840 1471.470 931.900 ;
        RECT 1472.070 931.840 1472.390 931.900 ;
        RECT 1471.150 931.700 1472.390 931.840 ;
        RECT 1471.150 931.640 1471.470 931.700 ;
        RECT 1472.070 931.640 1472.390 931.700 ;
        RECT 1471.150 883.220 1471.470 883.280 ;
        RECT 1472.070 883.220 1472.390 883.280 ;
        RECT 1471.150 883.080 1472.390 883.220 ;
        RECT 1471.150 883.020 1471.470 883.080 ;
        RECT 1472.070 883.020 1472.390 883.080 ;
        RECT 1471.150 835.280 1471.470 835.340 ;
        RECT 1472.070 835.280 1472.390 835.340 ;
        RECT 1471.150 835.140 1472.390 835.280 ;
        RECT 1471.150 835.080 1471.470 835.140 ;
        RECT 1472.070 835.080 1472.390 835.140 ;
        RECT 1472.070 786.660 1472.390 786.720 ;
        RECT 1472.990 786.660 1473.310 786.720 ;
        RECT 1472.070 786.520 1473.310 786.660 ;
        RECT 1472.070 786.460 1472.390 786.520 ;
        RECT 1472.990 786.460 1473.310 786.520 ;
        RECT 1472.070 738.380 1472.390 738.440 ;
        RECT 1472.990 738.380 1473.310 738.440 ;
        RECT 1472.070 738.240 1473.310 738.380 ;
        RECT 1472.070 738.180 1472.390 738.240 ;
        RECT 1472.990 738.180 1473.310 738.240 ;
        RECT 1471.150 712.540 1471.470 712.600 ;
        RECT 1472.070 712.540 1472.390 712.600 ;
        RECT 1471.150 712.400 1472.390 712.540 ;
        RECT 1471.150 712.340 1471.470 712.400 ;
        RECT 1472.070 712.340 1472.390 712.400 ;
        RECT 1471.150 641.820 1471.470 641.880 ;
        RECT 1472.070 641.820 1472.390 641.880 ;
        RECT 1471.150 641.680 1472.390 641.820 ;
        RECT 1471.150 641.620 1471.470 641.680 ;
        RECT 1472.070 641.620 1472.390 641.680 ;
        RECT 1472.070 593.880 1472.390 593.940 ;
        RECT 1472.990 593.880 1473.310 593.940 ;
        RECT 1472.070 593.740 1473.310 593.880 ;
        RECT 1472.070 593.680 1472.390 593.740 ;
        RECT 1472.990 593.680 1473.310 593.740 ;
        RECT 1472.070 545.260 1472.390 545.320 ;
        RECT 1472.990 545.260 1473.310 545.320 ;
        RECT 1472.070 545.120 1473.310 545.260 ;
        RECT 1472.070 545.060 1472.390 545.120 ;
        RECT 1472.990 545.060 1473.310 545.120 ;
        RECT 1471.150 521.120 1471.470 521.180 ;
        RECT 1472.070 521.120 1472.390 521.180 ;
        RECT 1471.150 520.980 1472.390 521.120 ;
        RECT 1471.150 520.920 1471.470 520.980 ;
        RECT 1472.070 520.920 1472.390 520.980 ;
        RECT 1471.150 448.020 1471.470 448.080 ;
        RECT 1473.450 448.020 1473.770 448.080 ;
        RECT 1471.150 447.880 1473.770 448.020 ;
        RECT 1471.150 447.820 1471.470 447.880 ;
        RECT 1473.450 447.820 1473.770 447.880 ;
        RECT 1472.070 352.140 1472.390 352.200 ;
        RECT 1472.990 352.140 1473.310 352.200 ;
        RECT 1472.070 352.000 1473.310 352.140 ;
        RECT 1472.070 351.940 1472.390 352.000 ;
        RECT 1472.990 351.940 1473.310 352.000 ;
        RECT 1472.070 326.980 1472.390 327.040 ;
        RECT 1472.990 326.980 1473.310 327.040 ;
        RECT 1472.070 326.840 1473.310 326.980 ;
        RECT 1472.070 326.780 1472.390 326.840 ;
        RECT 1472.990 326.780 1473.310 326.840 ;
        RECT 1472.070 255.580 1472.390 255.640 ;
        RECT 1472.990 255.580 1473.310 255.640 ;
        RECT 1472.070 255.440 1473.310 255.580 ;
        RECT 1472.070 255.380 1472.390 255.440 ;
        RECT 1472.990 255.380 1473.310 255.440 ;
        RECT 1472.070 206.960 1472.390 207.020 ;
        RECT 1472.990 206.960 1473.310 207.020 ;
        RECT 1472.070 206.820 1473.310 206.960 ;
        RECT 1472.070 206.760 1472.390 206.820 ;
        RECT 1472.990 206.760 1473.310 206.820 ;
        RECT 1472.070 164.800 1472.390 164.860 ;
        RECT 1472.990 164.800 1473.310 164.860 ;
        RECT 1472.070 164.660 1473.310 164.800 ;
        RECT 1472.070 164.600 1472.390 164.660 ;
        RECT 1472.990 164.600 1473.310 164.660 ;
        RECT 1471.150 96.800 1471.470 96.860 ;
        RECT 1472.070 96.800 1472.390 96.860 ;
        RECT 1471.150 96.660 1472.390 96.800 ;
        RECT 1471.150 96.600 1471.470 96.660 ;
        RECT 1472.070 96.600 1472.390 96.660 ;
        RECT 1185.950 24.720 1186.270 24.780 ;
        RECT 1471.150 24.720 1471.470 24.780 ;
        RECT 1185.950 24.580 1471.470 24.720 ;
        RECT 1185.950 24.520 1186.270 24.580 ;
        RECT 1471.150 24.520 1471.470 24.580 ;
      LAYER via ;
        RECT 1472.100 1683.380 1472.360 1683.640 ;
        RECT 1472.560 1635.440 1472.820 1635.700 ;
        RECT 1472.100 1545.680 1472.360 1545.940 ;
        RECT 1472.560 1545.680 1472.820 1545.940 ;
        RECT 1472.100 1417.840 1472.360 1418.100 ;
        RECT 1473.020 1417.840 1473.280 1418.100 ;
        RECT 1471.180 1388.940 1471.440 1389.200 ;
        RECT 1472.100 1388.940 1472.360 1389.200 ;
        RECT 1471.180 1317.880 1471.440 1318.140 ;
        RECT 1472.100 1317.880 1472.360 1318.140 ;
        RECT 1472.100 1269.600 1472.360 1269.860 ;
        RECT 1473.020 1269.600 1473.280 1269.860 ;
        RECT 1472.100 1221.320 1472.360 1221.580 ;
        RECT 1473.020 1221.320 1473.280 1221.580 ;
        RECT 1471.180 1197.180 1471.440 1197.440 ;
        RECT 1472.100 1197.180 1472.360 1197.440 ;
        RECT 1471.180 1124.760 1471.440 1125.020 ;
        RECT 1472.100 1124.760 1472.360 1125.020 ;
        RECT 1472.100 1076.480 1472.360 1076.740 ;
        RECT 1473.020 1076.480 1473.280 1076.740 ;
        RECT 1472.100 1028.200 1472.360 1028.460 ;
        RECT 1473.020 1028.200 1473.280 1028.460 ;
        RECT 1471.180 979.580 1471.440 979.840 ;
        RECT 1472.100 979.580 1472.360 979.840 ;
        RECT 1471.180 931.640 1471.440 931.900 ;
        RECT 1472.100 931.640 1472.360 931.900 ;
        RECT 1471.180 883.020 1471.440 883.280 ;
        RECT 1472.100 883.020 1472.360 883.280 ;
        RECT 1471.180 835.080 1471.440 835.340 ;
        RECT 1472.100 835.080 1472.360 835.340 ;
        RECT 1472.100 786.460 1472.360 786.720 ;
        RECT 1473.020 786.460 1473.280 786.720 ;
        RECT 1472.100 738.180 1472.360 738.440 ;
        RECT 1473.020 738.180 1473.280 738.440 ;
        RECT 1471.180 712.340 1471.440 712.600 ;
        RECT 1472.100 712.340 1472.360 712.600 ;
        RECT 1471.180 641.620 1471.440 641.880 ;
        RECT 1472.100 641.620 1472.360 641.880 ;
        RECT 1472.100 593.680 1472.360 593.940 ;
        RECT 1473.020 593.680 1473.280 593.940 ;
        RECT 1472.100 545.060 1472.360 545.320 ;
        RECT 1473.020 545.060 1473.280 545.320 ;
        RECT 1471.180 520.920 1471.440 521.180 ;
        RECT 1472.100 520.920 1472.360 521.180 ;
        RECT 1471.180 447.820 1471.440 448.080 ;
        RECT 1473.480 447.820 1473.740 448.080 ;
        RECT 1472.100 351.940 1472.360 352.200 ;
        RECT 1473.020 351.940 1473.280 352.200 ;
        RECT 1472.100 326.780 1472.360 327.040 ;
        RECT 1473.020 326.780 1473.280 327.040 ;
        RECT 1472.100 255.380 1472.360 255.640 ;
        RECT 1473.020 255.380 1473.280 255.640 ;
        RECT 1472.100 206.760 1472.360 207.020 ;
        RECT 1473.020 206.760 1473.280 207.020 ;
        RECT 1472.100 164.600 1472.360 164.860 ;
        RECT 1473.020 164.600 1473.280 164.860 ;
        RECT 1471.180 96.600 1471.440 96.860 ;
        RECT 1472.100 96.600 1472.360 96.860 ;
        RECT 1185.980 24.520 1186.240 24.780 ;
        RECT 1471.180 24.520 1471.440 24.780 ;
      LAYER met2 ;
        RECT 1471.170 1700.410 1471.450 1704.000 ;
        RECT 1471.170 1700.270 1471.840 1700.410 ;
        RECT 1471.170 1700.000 1471.450 1700.270 ;
        RECT 1471.700 1695.650 1471.840 1700.270 ;
        RECT 1471.700 1695.510 1472.300 1695.650 ;
        RECT 1472.160 1683.670 1472.300 1695.510 ;
        RECT 1472.100 1683.350 1472.360 1683.670 ;
        RECT 1472.560 1635.410 1472.820 1635.730 ;
        RECT 1472.620 1618.130 1472.760 1635.410 ;
        RECT 1472.160 1617.990 1472.760 1618.130 ;
        RECT 1472.160 1545.970 1472.300 1617.990 ;
        RECT 1472.100 1545.650 1472.360 1545.970 ;
        RECT 1472.560 1545.650 1472.820 1545.970 ;
        RECT 1472.620 1545.370 1472.760 1545.650 ;
        RECT 1472.620 1545.230 1473.220 1545.370 ;
        RECT 1473.080 1418.130 1473.220 1545.230 ;
        RECT 1472.100 1417.810 1472.360 1418.130 ;
        RECT 1473.020 1417.810 1473.280 1418.130 ;
        RECT 1472.160 1389.230 1472.300 1417.810 ;
        RECT 1471.180 1388.910 1471.440 1389.230 ;
        RECT 1472.100 1388.910 1472.360 1389.230 ;
        RECT 1471.240 1318.170 1471.380 1388.910 ;
        RECT 1471.180 1317.850 1471.440 1318.170 ;
        RECT 1472.100 1317.850 1472.360 1318.170 ;
        RECT 1472.160 1269.890 1472.300 1317.850 ;
        RECT 1472.100 1269.570 1472.360 1269.890 ;
        RECT 1473.020 1269.570 1473.280 1269.890 ;
        RECT 1473.080 1221.610 1473.220 1269.570 ;
        RECT 1472.100 1221.290 1472.360 1221.610 ;
        RECT 1473.020 1221.290 1473.280 1221.610 ;
        RECT 1472.160 1197.470 1472.300 1221.290 ;
        RECT 1471.180 1197.150 1471.440 1197.470 ;
        RECT 1472.100 1197.150 1472.360 1197.470 ;
        RECT 1471.240 1125.050 1471.380 1197.150 ;
        RECT 1471.180 1124.730 1471.440 1125.050 ;
        RECT 1472.100 1124.730 1472.360 1125.050 ;
        RECT 1472.160 1076.770 1472.300 1124.730 ;
        RECT 1472.100 1076.450 1472.360 1076.770 ;
        RECT 1473.020 1076.450 1473.280 1076.770 ;
        RECT 1473.080 1028.490 1473.220 1076.450 ;
        RECT 1472.100 1028.170 1472.360 1028.490 ;
        RECT 1473.020 1028.170 1473.280 1028.490 ;
        RECT 1472.160 979.870 1472.300 1028.170 ;
        RECT 1471.180 979.550 1471.440 979.870 ;
        RECT 1472.100 979.550 1472.360 979.870 ;
        RECT 1471.240 931.930 1471.380 979.550 ;
        RECT 1471.180 931.610 1471.440 931.930 ;
        RECT 1472.100 931.610 1472.360 931.930 ;
        RECT 1472.160 883.310 1472.300 931.610 ;
        RECT 1471.180 882.990 1471.440 883.310 ;
        RECT 1472.100 882.990 1472.360 883.310 ;
        RECT 1471.240 835.370 1471.380 882.990 ;
        RECT 1471.180 835.050 1471.440 835.370 ;
        RECT 1472.100 835.050 1472.360 835.370 ;
        RECT 1472.160 786.750 1472.300 835.050 ;
        RECT 1472.100 786.430 1472.360 786.750 ;
        RECT 1473.020 786.430 1473.280 786.750 ;
        RECT 1473.080 738.470 1473.220 786.430 ;
        RECT 1472.100 738.150 1472.360 738.470 ;
        RECT 1473.020 738.150 1473.280 738.470 ;
        RECT 1472.160 712.630 1472.300 738.150 ;
        RECT 1471.180 712.310 1471.440 712.630 ;
        RECT 1472.100 712.310 1472.360 712.630 ;
        RECT 1471.240 641.910 1471.380 712.310 ;
        RECT 1471.180 641.590 1471.440 641.910 ;
        RECT 1472.100 641.590 1472.360 641.910 ;
        RECT 1472.160 593.970 1472.300 641.590 ;
        RECT 1472.100 593.650 1472.360 593.970 ;
        RECT 1473.020 593.650 1473.280 593.970 ;
        RECT 1473.080 545.350 1473.220 593.650 ;
        RECT 1472.100 545.030 1472.360 545.350 ;
        RECT 1473.020 545.030 1473.280 545.350 ;
        RECT 1472.160 521.210 1472.300 545.030 ;
        RECT 1471.180 520.890 1471.440 521.210 ;
        RECT 1472.100 520.890 1472.360 521.210 ;
        RECT 1471.240 448.110 1471.380 520.890 ;
        RECT 1471.180 447.790 1471.440 448.110 ;
        RECT 1473.480 447.790 1473.740 448.110 ;
        RECT 1473.540 400.930 1473.680 447.790 ;
        RECT 1473.080 400.790 1473.680 400.930 ;
        RECT 1473.080 352.230 1473.220 400.790 ;
        RECT 1472.100 351.910 1472.360 352.230 ;
        RECT 1473.020 351.910 1473.280 352.230 ;
        RECT 1472.160 327.070 1472.300 351.910 ;
        RECT 1472.100 326.750 1472.360 327.070 ;
        RECT 1473.020 326.750 1473.280 327.070 ;
        RECT 1473.080 255.670 1473.220 326.750 ;
        RECT 1472.100 255.350 1472.360 255.670 ;
        RECT 1473.020 255.350 1473.280 255.670 ;
        RECT 1472.160 207.050 1472.300 255.350 ;
        RECT 1472.100 206.730 1472.360 207.050 ;
        RECT 1473.020 206.730 1473.280 207.050 ;
        RECT 1473.080 164.890 1473.220 206.730 ;
        RECT 1472.100 164.570 1472.360 164.890 ;
        RECT 1473.020 164.570 1473.280 164.890 ;
        RECT 1472.160 96.890 1472.300 164.570 ;
        RECT 1471.180 96.570 1471.440 96.890 ;
        RECT 1472.100 96.570 1472.360 96.890 ;
        RECT 1471.240 24.810 1471.380 96.570 ;
        RECT 1185.980 24.490 1186.240 24.810 ;
        RECT 1471.180 24.490 1471.440 24.810 ;
        RECT 1186.040 2.400 1186.180 24.490 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1470.230 1678.140 1470.550 1678.200 ;
        RECT 1474.830 1678.140 1475.150 1678.200 ;
        RECT 1470.230 1678.000 1475.150 1678.140 ;
        RECT 1470.230 1677.940 1470.550 1678.000 ;
        RECT 1474.830 1677.940 1475.150 1678.000 ;
        RECT 1203.890 25.060 1204.210 25.120 ;
        RECT 1470.230 25.060 1470.550 25.120 ;
        RECT 1203.890 24.920 1470.550 25.060 ;
        RECT 1203.890 24.860 1204.210 24.920 ;
        RECT 1470.230 24.860 1470.550 24.920 ;
      LAYER via ;
        RECT 1470.260 1677.940 1470.520 1678.200 ;
        RECT 1474.860 1677.940 1475.120 1678.200 ;
        RECT 1203.920 24.860 1204.180 25.120 ;
        RECT 1470.260 24.860 1470.520 25.120 ;
      LAYER met2 ;
        RECT 1476.230 1700.410 1476.510 1704.000 ;
        RECT 1474.920 1700.270 1476.510 1700.410 ;
        RECT 1474.920 1678.230 1475.060 1700.270 ;
        RECT 1476.230 1700.000 1476.510 1700.270 ;
        RECT 1470.260 1677.910 1470.520 1678.230 ;
        RECT 1474.860 1677.910 1475.120 1678.230 ;
        RECT 1470.320 25.150 1470.460 1677.910 ;
        RECT 1203.920 24.830 1204.180 25.150 ;
        RECT 1470.260 24.830 1470.520 25.150 ;
        RECT 1203.980 2.400 1204.120 24.830 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1203.910 19.240 1204.190 19.520 ;
        RECT 1470.710 19.240 1470.990 19.520 ;
      LAYER met3 ;
        RECT 1203.885 19.530 1204.215 19.545 ;
        RECT 1470.685 19.530 1471.015 19.545 ;
        RECT 1203.885 19.230 1471.015 19.530 ;
        RECT 1203.885 19.215 1204.215 19.230 ;
        RECT 1470.685 19.215 1471.015 19.230 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 0.300 ;
=======
      LAYER li1 ;
        RECT 1422.925 14.025 1423.095 17.935 ;
      LAYER mcon ;
        RECT 1422.925 17.765 1423.095 17.935 ;
      LAYER met1 ;
        RECT 1477.590 1666.240 1477.910 1666.300 ;
        RECT 1478.510 1666.240 1478.830 1666.300 ;
        RECT 1477.590 1666.100 1478.830 1666.240 ;
        RECT 1477.590 1666.040 1477.910 1666.100 ;
        RECT 1478.510 1666.040 1478.830 1666.100 ;
        RECT 1221.830 17.920 1222.150 17.980 ;
        RECT 1422.865 17.920 1423.155 17.965 ;
        RECT 1221.830 17.780 1423.155 17.920 ;
        RECT 1221.830 17.720 1222.150 17.780 ;
        RECT 1422.865 17.735 1423.155 17.780 ;
        RECT 1422.865 14.180 1423.155 14.225 ;
        RECT 1422.865 14.040 1471.380 14.180 ;
        RECT 1422.865 13.995 1423.155 14.040 ;
        RECT 1471.240 13.840 1471.380 14.040 ;
        RECT 1478.050 13.840 1478.370 13.900 ;
        RECT 1471.240 13.700 1478.370 13.840 ;
        RECT 1478.050 13.640 1478.370 13.700 ;
      LAYER via ;
        RECT 1477.620 1666.040 1477.880 1666.300 ;
        RECT 1478.540 1666.040 1478.800 1666.300 ;
        RECT 1221.860 17.720 1222.120 17.980 ;
        RECT 1478.080 13.640 1478.340 13.900 ;
      LAYER met2 ;
        RECT 1479.450 1700.410 1479.730 1704.000 ;
        RECT 1478.600 1700.270 1479.730 1700.410 ;
        RECT 1478.600 1666.330 1478.740 1700.270 ;
        RECT 1479.450 1700.000 1479.730 1700.270 ;
        RECT 1477.620 1666.010 1477.880 1666.330 ;
        RECT 1478.540 1666.010 1478.800 1666.330 ;
        RECT 1477.680 37.810 1477.820 1666.010 ;
        RECT 1477.680 37.670 1478.280 37.810 ;
        RECT 1221.860 17.690 1222.120 18.010 ;
        RECT 1221.920 2.400 1222.060 17.690 ;
        RECT 1478.140 13.930 1478.280 37.670 ;
        RECT 1478.080 13.610 1478.340 13.930 ;
=======
      LAYER met1 ;
        RECT 1221.830 25.400 1222.150 25.460 ;
        RECT 1478.050 25.400 1478.370 25.460 ;
        RECT 1221.830 25.260 1478.370 25.400 ;
        RECT 1221.830 25.200 1222.150 25.260 ;
        RECT 1478.050 25.200 1478.370 25.260 ;
      LAYER via ;
        RECT 1221.860 25.200 1222.120 25.460 ;
        RECT 1478.080 25.200 1478.340 25.460 ;
      LAYER met2 ;
        RECT 1480.830 1700.410 1481.110 1704.000 ;
        RECT 1480.440 1700.270 1481.110 1700.410 ;
        RECT 1480.440 1677.290 1480.580 1700.270 ;
        RECT 1480.830 1700.000 1481.110 1700.270 ;
        RECT 1478.140 1677.150 1480.580 1677.290 ;
        RECT 1478.140 25.490 1478.280 1677.150 ;
        RECT 1221.860 25.170 1222.120 25.490 ;
        RECT 1478.080 25.170 1478.340 25.490 ;
        RECT 1221.920 2.400 1222.060 25.170 ;
>>>>>>> re-updated local openlane
        RECT 1221.710 -4.800 1222.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 0.300 ;
=======
      LAYER li1 ;
        RECT 1463.865 18.445 1464.955 18.615 ;
      LAYER mcon ;
        RECT 1464.785 18.445 1464.955 18.615 ;
      LAYER met1 ;
        RECT 1239.770 18.600 1240.090 18.660 ;
        RECT 1463.805 18.600 1464.095 18.645 ;
        RECT 1239.770 18.460 1464.095 18.600 ;
        RECT 1239.770 18.400 1240.090 18.460 ;
        RECT 1463.805 18.415 1464.095 18.460 ;
        RECT 1464.725 18.600 1465.015 18.645 ;
        RECT 1484.950 18.600 1485.270 18.660 ;
        RECT 1464.725 18.460 1485.270 18.600 ;
        RECT 1464.725 18.415 1465.015 18.460 ;
        RECT 1484.950 18.400 1485.270 18.460 ;
      LAYER via ;
        RECT 1239.800 18.400 1240.060 18.660 ;
        RECT 1484.980 18.400 1485.240 18.660 ;
      LAYER met2 ;
        RECT 1484.510 1700.410 1484.790 1704.000 ;
        RECT 1484.510 1700.270 1485.180 1700.410 ;
        RECT 1484.510 1700.000 1484.790 1700.270 ;
        RECT 1485.040 18.690 1485.180 1700.270 ;
        RECT 1239.800 18.370 1240.060 18.690 ;
        RECT 1484.980 18.370 1485.240 18.690 ;
        RECT 1239.860 2.400 1240.000 18.370 ;
=======
      LAYER met1 ;
        RECT 1239.770 25.740 1240.090 25.800 ;
        RECT 1485.410 25.740 1485.730 25.800 ;
        RECT 1239.770 25.600 1485.730 25.740 ;
        RECT 1239.770 25.540 1240.090 25.600 ;
        RECT 1485.410 25.540 1485.730 25.600 ;
      LAYER via ;
        RECT 1239.800 25.540 1240.060 25.800 ;
        RECT 1485.440 25.540 1485.700 25.800 ;
      LAYER met2 ;
        RECT 1485.890 1700.410 1486.170 1704.000 ;
        RECT 1485.500 1700.270 1486.170 1700.410 ;
        RECT 1485.500 25.830 1485.640 1700.270 ;
        RECT 1485.890 1700.000 1486.170 1700.270 ;
        RECT 1239.800 25.510 1240.060 25.830 ;
        RECT 1485.440 25.510 1485.700 25.830 ;
        RECT 1239.860 2.400 1240.000 25.510 ;
>>>>>>> re-updated local openlane
        RECT 1239.650 -4.800 1240.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1257.250 26.080 1257.570 26.140 ;
        RECT 1490.930 26.080 1491.250 26.140 ;
        RECT 1257.250 25.940 1491.250 26.080 ;
        RECT 1257.250 25.880 1257.570 25.940 ;
        RECT 1490.930 25.880 1491.250 25.940 ;
      LAYER via ;
        RECT 1257.280 25.880 1257.540 26.140 ;
        RECT 1490.960 25.880 1491.220 26.140 ;
      LAYER met2 ;
        RECT 1490.490 1700.410 1490.770 1704.000 ;
        RECT 1490.490 1700.270 1491.160 1700.410 ;
        RECT 1490.490 1700.000 1490.770 1700.270 ;
        RECT 1491.020 26.170 1491.160 1700.270 ;
        RECT 1257.280 25.850 1257.540 26.170 ;
        RECT 1490.960 25.850 1491.220 26.170 ;
        RECT 1257.340 2.400 1257.480 25.850 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 0.300 ;
=======
      LAYER li1 ;
        RECT 1494.225 531.505 1494.395 620.755 ;
        RECT 1493.765 96.645 1493.935 110.755 ;
      LAYER mcon ;
        RECT 1494.225 620.585 1494.395 620.755 ;
        RECT 1493.765 110.585 1493.935 110.755 ;
      LAYER met1 ;
        RECT 1493.690 1062.740 1494.010 1062.800 ;
        RECT 1494.610 1062.740 1494.930 1062.800 ;
        RECT 1493.690 1062.600 1494.930 1062.740 ;
        RECT 1493.690 1062.540 1494.010 1062.600 ;
        RECT 1494.610 1062.540 1494.930 1062.600 ;
        RECT 1493.690 979.580 1494.010 979.840 ;
        RECT 1493.780 979.160 1493.920 979.580 ;
        RECT 1493.690 978.900 1494.010 979.160 ;
        RECT 1493.690 641.620 1494.010 641.880 ;
        RECT 1493.780 641.480 1493.920 641.620 ;
        RECT 1494.150 641.480 1494.470 641.540 ;
        RECT 1493.780 641.340 1494.470 641.480 ;
        RECT 1494.150 641.280 1494.470 641.340 ;
        RECT 1494.150 627.880 1494.470 627.940 ;
        RECT 1495.070 627.880 1495.390 627.940 ;
        RECT 1494.150 627.740 1495.390 627.880 ;
        RECT 1494.150 627.680 1494.470 627.740 ;
        RECT 1495.070 627.680 1495.390 627.740 ;
        RECT 1494.165 620.740 1494.455 620.785 ;
        RECT 1495.070 620.740 1495.390 620.800 ;
        RECT 1494.165 620.600 1495.390 620.740 ;
        RECT 1494.165 620.555 1494.455 620.600 ;
        RECT 1495.070 620.540 1495.390 620.600 ;
        RECT 1494.150 531.660 1494.470 531.720 ;
        RECT 1493.955 531.520 1494.470 531.660 ;
        RECT 1494.150 531.460 1494.470 531.520 ;
        RECT 1494.150 304.200 1494.470 304.260 ;
        RECT 1493.780 304.060 1494.470 304.200 ;
        RECT 1493.780 303.920 1493.920 304.060 ;
        RECT 1494.150 304.000 1494.470 304.060 ;
        RECT 1493.690 303.660 1494.010 303.920 ;
        RECT 1493.705 110.740 1493.995 110.785 ;
        RECT 1494.150 110.740 1494.470 110.800 ;
        RECT 1493.705 110.600 1494.470 110.740 ;
        RECT 1493.705 110.555 1493.995 110.600 ;
        RECT 1494.150 110.540 1494.470 110.600 ;
        RECT 1493.690 96.800 1494.010 96.860 ;
        RECT 1493.495 96.660 1494.010 96.800 ;
        RECT 1493.690 96.600 1494.010 96.660 ;
        RECT 1276.110 59.400 1276.430 59.460 ;
        RECT 1493.690 59.400 1494.010 59.460 ;
        RECT 1276.110 59.260 1494.010 59.400 ;
        RECT 1276.110 59.200 1276.430 59.260 ;
        RECT 1493.690 59.200 1494.010 59.260 ;
      LAYER via ;
        RECT 1493.720 1062.540 1493.980 1062.800 ;
        RECT 1494.640 1062.540 1494.900 1062.800 ;
        RECT 1493.720 979.580 1493.980 979.840 ;
        RECT 1493.720 978.900 1493.980 979.160 ;
        RECT 1493.720 641.620 1493.980 641.880 ;
        RECT 1494.180 641.280 1494.440 641.540 ;
        RECT 1494.180 627.680 1494.440 627.940 ;
        RECT 1495.100 627.680 1495.360 627.940 ;
        RECT 1495.100 620.540 1495.360 620.800 ;
        RECT 1494.180 531.460 1494.440 531.720 ;
        RECT 1494.180 304.000 1494.440 304.260 ;
        RECT 1493.720 303.660 1493.980 303.920 ;
        RECT 1494.180 110.540 1494.440 110.800 ;
        RECT 1493.720 96.600 1493.980 96.860 ;
        RECT 1276.140 59.200 1276.400 59.460 ;
        RECT 1493.720 59.200 1493.980 59.460 ;
      LAYER met2 ;
        RECT 1495.550 1700.410 1495.830 1704.000 ;
        RECT 1494.700 1700.270 1495.830 1700.410 ;
        RECT 1494.700 1678.140 1494.840 1700.270 ;
        RECT 1495.550 1700.000 1495.830 1700.270 ;
        RECT 1493.780 1678.000 1494.840 1678.140 ;
        RECT 1493.780 1618.130 1493.920 1678.000 ;
        RECT 1493.780 1617.990 1494.380 1618.130 ;
        RECT 1494.240 1463.090 1494.380 1617.990 ;
        RECT 1493.320 1462.950 1494.380 1463.090 ;
        RECT 1493.320 1462.410 1493.460 1462.950 ;
        RECT 1493.320 1462.270 1494.380 1462.410 ;
        RECT 1494.240 1365.850 1494.380 1462.270 ;
        RECT 1493.780 1365.710 1494.380 1365.850 ;
        RECT 1493.780 1318.250 1493.920 1365.710 ;
        RECT 1493.320 1318.110 1493.920 1318.250 ;
        RECT 1493.320 1317.570 1493.460 1318.110 ;
        RECT 1493.320 1317.430 1494.380 1317.570 ;
        RECT 1494.240 1173.410 1494.380 1317.430 ;
        RECT 1493.320 1173.270 1494.380 1173.410 ;
        RECT 1493.320 1172.730 1493.460 1173.270 ;
        RECT 1493.320 1172.590 1493.920 1172.730 ;
        RECT 1493.780 1110.965 1493.920 1172.590 ;
        RECT 1493.710 1110.595 1493.990 1110.965 ;
        RECT 1494.630 1110.595 1494.910 1110.965 ;
        RECT 1494.700 1062.830 1494.840 1110.595 ;
        RECT 1493.720 1062.510 1493.980 1062.830 ;
        RECT 1494.640 1062.510 1494.900 1062.830 ;
        RECT 1493.780 979.870 1493.920 1062.510 ;
        RECT 1493.720 979.550 1493.980 979.870 ;
        RECT 1493.720 978.870 1493.980 979.190 ;
        RECT 1493.780 845.650 1493.920 978.870 ;
        RECT 1493.320 845.510 1493.920 845.650 ;
        RECT 1493.320 821.285 1493.460 845.510 ;
        RECT 1493.250 820.915 1493.530 821.285 ;
        RECT 1494.630 820.915 1494.910 821.285 ;
        RECT 1494.700 773.005 1494.840 820.915 ;
        RECT 1493.710 772.635 1493.990 773.005 ;
        RECT 1494.630 772.635 1494.910 773.005 ;
        RECT 1493.780 690.610 1493.920 772.635 ;
        RECT 1493.320 690.470 1493.920 690.610 ;
        RECT 1493.320 689.930 1493.460 690.470 ;
        RECT 1493.320 689.790 1493.920 689.930 ;
        RECT 1493.780 641.910 1493.920 689.790 ;
        RECT 1493.720 641.590 1493.980 641.910 ;
        RECT 1494.180 641.250 1494.440 641.570 ;
        RECT 1494.240 627.970 1494.380 641.250 ;
        RECT 1494.180 627.650 1494.440 627.970 ;
        RECT 1495.100 627.650 1495.360 627.970 ;
        RECT 1495.160 620.830 1495.300 627.650 ;
        RECT 1495.100 620.510 1495.360 620.830 ;
        RECT 1494.180 531.430 1494.440 531.750 ;
        RECT 1494.240 304.290 1494.380 531.430 ;
        RECT 1494.180 303.970 1494.440 304.290 ;
        RECT 1493.720 303.630 1493.980 303.950 ;
        RECT 1493.780 303.010 1493.920 303.630 ;
        RECT 1493.780 302.870 1494.380 303.010 ;
        RECT 1494.240 110.830 1494.380 302.870 ;
        RECT 1494.180 110.510 1494.440 110.830 ;
        RECT 1493.720 96.570 1493.980 96.890 ;
        RECT 1493.780 59.490 1493.920 96.570 ;
        RECT 1276.140 59.170 1276.400 59.490 ;
        RECT 1493.720 59.170 1493.980 59.490 ;
        RECT 1276.200 5.850 1276.340 59.170 ;
        RECT 1275.280 5.710 1276.340 5.850 ;
        RECT 1275.280 2.400 1275.420 5.710 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
      LAYER via2 ;
        RECT 1493.710 1110.640 1493.990 1110.920 ;
        RECT 1494.630 1110.640 1494.910 1110.920 ;
        RECT 1493.250 820.960 1493.530 821.240 ;
        RECT 1494.630 820.960 1494.910 821.240 ;
        RECT 1493.710 772.680 1493.990 772.960 ;
        RECT 1494.630 772.680 1494.910 772.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1492.305 531.570 1492.635 531.585 ;
        RECT 1492.305 531.255 1492.850 531.570 ;
        RECT 1492.550 530.890 1492.850 531.255 ;
        RECT 1493.225 530.890 1493.555 530.905 ;
        RECT 1492.550 530.590 1493.555 530.890 ;
        RECT 1493.225 530.575 1493.555 530.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1493.685 1110.930 1494.015 1110.945 ;
        RECT 1494.605 1110.930 1494.935 1110.945 ;
        RECT 1493.685 1110.630 1494.935 1110.930 ;
        RECT 1493.685 1110.615 1494.015 1110.630 ;
        RECT 1494.605 1110.615 1494.935 1110.630 ;
        RECT 1493.225 821.250 1493.555 821.265 ;
        RECT 1494.605 821.250 1494.935 821.265 ;
        RECT 1493.225 820.950 1494.935 821.250 ;
        RECT 1493.225 820.935 1493.555 820.950 ;
        RECT 1494.605 820.935 1494.935 820.950 ;
        RECT 1493.685 772.970 1494.015 772.985 ;
        RECT 1494.605 772.970 1494.935 772.985 ;
        RECT 1493.685 772.670 1494.935 772.970 ;
        RECT 1493.685 772.655 1494.015 772.670 ;
        RECT 1494.605 772.655 1494.935 772.670 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 0.300 ;
=======
      LAYER li1 ;
        RECT 1463.405 18.275 1463.575 19.295 ;
        RECT 1463.405 18.105 1465.875 18.275 ;
        RECT 1465.705 17.085 1465.875 18.105 ;
      LAYER mcon ;
        RECT 1463.405 19.125 1463.575 19.295 ;
      LAYER met1 ;
        RECT 1293.130 19.280 1293.450 19.340 ;
        RECT 1463.345 19.280 1463.635 19.325 ;
        RECT 1293.130 19.140 1463.635 19.280 ;
        RECT 1293.130 19.080 1293.450 19.140 ;
        RECT 1463.345 19.095 1463.635 19.140 ;
        RECT 1487.250 18.260 1487.570 18.320 ;
        RECT 1498.750 18.260 1499.070 18.320 ;
        RECT 1487.250 18.120 1499.070 18.260 ;
        RECT 1487.250 18.060 1487.570 18.120 ;
        RECT 1498.750 18.060 1499.070 18.120 ;
        RECT 1465.645 17.240 1465.935 17.285 ;
        RECT 1484.030 17.240 1484.350 17.300 ;
        RECT 1465.645 17.100 1484.350 17.240 ;
        RECT 1465.645 17.055 1465.935 17.100 ;
        RECT 1484.030 17.040 1484.350 17.100 ;
      LAYER via ;
        RECT 1293.160 19.080 1293.420 19.340 ;
        RECT 1487.280 18.060 1487.540 18.320 ;
        RECT 1498.780 18.060 1499.040 18.320 ;
        RECT 1484.060 17.040 1484.320 17.300 ;
      LAYER met2 ;
        RECT 1498.770 1700.000 1499.050 1704.000 ;
        RECT 1293.160 19.050 1293.420 19.370 ;
        RECT 1293.220 2.400 1293.360 19.050 ;
        RECT 1498.840 18.350 1498.980 1700.000 ;
        RECT 1484.120 17.950 1485.180 18.090 ;
        RECT 1487.280 18.030 1487.540 18.350 ;
        RECT 1498.780 18.030 1499.040 18.350 ;
        RECT 1484.120 17.330 1484.260 17.950 ;
        RECT 1485.040 17.410 1485.180 17.950 ;
        RECT 1487.340 17.410 1487.480 18.030 ;
        RECT 1484.060 17.010 1484.320 17.330 ;
        RECT 1485.040 17.270 1487.480 17.410 ;
=======
      LAYER met1 ;
        RECT 1296.810 1638.700 1297.130 1638.760 ;
        RECT 1497.830 1638.700 1498.150 1638.760 ;
        RECT 1296.810 1638.560 1498.150 1638.700 ;
        RECT 1296.810 1638.500 1297.130 1638.560 ;
        RECT 1497.830 1638.500 1498.150 1638.560 ;
        RECT 1293.130 20.640 1293.450 20.700 ;
        RECT 1296.810 20.640 1297.130 20.700 ;
        RECT 1293.130 20.500 1297.130 20.640 ;
        RECT 1293.130 20.440 1293.450 20.500 ;
        RECT 1296.810 20.440 1297.130 20.500 ;
      LAYER via ;
        RECT 1296.840 1638.500 1297.100 1638.760 ;
        RECT 1497.860 1638.500 1498.120 1638.760 ;
        RECT 1293.160 20.440 1293.420 20.700 ;
        RECT 1296.840 20.440 1297.100 20.700 ;
      LAYER met2 ;
        RECT 1500.150 1700.410 1500.430 1704.000 ;
        RECT 1499.300 1700.270 1500.430 1700.410 ;
        RECT 1499.300 1676.610 1499.440 1700.270 ;
        RECT 1500.150 1700.000 1500.430 1700.270 ;
        RECT 1497.920 1676.470 1499.440 1676.610 ;
        RECT 1497.920 1638.790 1498.060 1676.470 ;
        RECT 1296.840 1638.470 1297.100 1638.790 ;
        RECT 1497.860 1638.470 1498.120 1638.790 ;
        RECT 1296.900 20.730 1297.040 1638.470 ;
        RECT 1293.160 20.410 1293.420 20.730 ;
        RECT 1296.840 20.410 1297.100 20.730 ;
        RECT 1293.220 2.400 1293.360 20.410 ;
>>>>>>> re-updated local openlane
        RECT 1293.010 -4.800 1293.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 0.300 ;
=======
      LAYER met1 ;
        RECT 1311.530 51.580 1311.850 51.640 ;
        RECT 1505.190 51.580 1505.510 51.640 ;
        RECT 1311.530 51.440 1505.510 51.580 ;
        RECT 1311.530 51.380 1311.850 51.440 ;
        RECT 1505.190 51.380 1505.510 51.440 ;
      LAYER via ;
        RECT 1311.560 51.380 1311.820 51.640 ;
        RECT 1505.220 51.380 1505.480 51.640 ;
      LAYER met2 ;
        RECT 1505.210 1700.000 1505.490 1704.000 ;
        RECT 1505.280 51.670 1505.420 1700.000 ;
        RECT 1311.560 51.350 1311.820 51.670 ;
        RECT 1505.220 51.350 1505.480 51.670 ;
        RECT 1311.620 33.050 1311.760 51.350 ;
        RECT 1311.160 32.910 1311.760 33.050 ;
        RECT 1311.160 2.400 1311.300 32.910 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 0.300 ;
=======
      LAYER li1 ;
        RECT 1505.725 1338.665 1505.895 1366.035 ;
        RECT 1505.725 766.105 1505.895 814.215 ;
      LAYER mcon ;
        RECT 1505.725 1365.865 1505.895 1366.035 ;
        RECT 1505.725 814.045 1505.895 814.215 ;
      LAYER met1 ;
        RECT 1505.650 1642.440 1505.970 1642.500 ;
        RECT 1507.030 1642.440 1507.350 1642.500 ;
        RECT 1505.650 1642.300 1507.350 1642.440 ;
        RECT 1505.650 1642.240 1505.970 1642.300 ;
        RECT 1507.030 1642.240 1507.350 1642.300 ;
        RECT 1505.650 1366.020 1505.970 1366.080 ;
        RECT 1505.455 1365.880 1505.970 1366.020 ;
        RECT 1505.650 1365.820 1505.970 1365.880 ;
        RECT 1505.650 1338.820 1505.970 1338.880 ;
        RECT 1505.455 1338.680 1505.970 1338.820 ;
        RECT 1505.650 1338.620 1505.970 1338.680 ;
        RECT 1505.650 1257.700 1505.970 1257.960 ;
        RECT 1505.740 1257.280 1505.880 1257.700 ;
        RECT 1505.650 1257.020 1505.970 1257.280 ;
        RECT 1504.730 886.620 1505.050 886.680 ;
        RECT 1505.650 886.620 1505.970 886.680 ;
        RECT 1504.730 886.480 1505.970 886.620 ;
        RECT 1504.730 886.420 1505.050 886.480 ;
        RECT 1505.650 886.420 1505.970 886.480 ;
        RECT 1505.650 814.200 1505.970 814.260 ;
        RECT 1505.455 814.060 1505.970 814.200 ;
        RECT 1505.650 814.000 1505.970 814.060 ;
        RECT 1505.650 766.260 1505.970 766.320 ;
        RECT 1505.455 766.120 1505.970 766.260 ;
        RECT 1505.650 766.060 1505.970 766.120 ;
        RECT 1506.110 676.300 1506.430 676.560 ;
        RECT 1506.200 675.820 1506.340 676.300 ;
        RECT 1506.570 675.820 1506.890 675.880 ;
        RECT 1506.200 675.680 1506.890 675.820 ;
        RECT 1506.570 675.620 1506.890 675.680 ;
        RECT 1505.650 593.340 1505.970 593.600 ;
        RECT 1505.740 592.920 1505.880 593.340 ;
        RECT 1505.650 592.660 1505.970 592.920 ;
        RECT 1505.190 62.460 1505.510 62.520 ;
        RECT 1504.820 62.320 1505.510 62.460 ;
        RECT 1504.820 62.180 1504.960 62.320 ;
        RECT 1505.190 62.260 1505.510 62.320 ;
        RECT 1504.730 61.920 1505.050 62.180 ;
        RECT 1329.010 25.740 1329.330 25.800 ;
        RECT 1504.730 25.740 1505.050 25.800 ;
        RECT 1329.010 25.600 1505.050 25.740 ;
        RECT 1329.010 25.540 1329.330 25.600 ;
        RECT 1504.730 25.540 1505.050 25.600 ;
      LAYER via ;
        RECT 1505.680 1642.240 1505.940 1642.500 ;
        RECT 1507.060 1642.240 1507.320 1642.500 ;
        RECT 1505.680 1365.820 1505.940 1366.080 ;
        RECT 1505.680 1338.620 1505.940 1338.880 ;
        RECT 1505.680 1257.700 1505.940 1257.960 ;
        RECT 1505.680 1257.020 1505.940 1257.280 ;
        RECT 1504.760 886.420 1505.020 886.680 ;
        RECT 1505.680 886.420 1505.940 886.680 ;
        RECT 1505.680 814.000 1505.940 814.260 ;
        RECT 1505.680 766.060 1505.940 766.320 ;
        RECT 1506.140 676.300 1506.400 676.560 ;
        RECT 1506.600 675.620 1506.860 675.880 ;
        RECT 1505.680 593.340 1505.940 593.600 ;
        RECT 1505.680 592.660 1505.940 592.920 ;
        RECT 1505.220 62.260 1505.480 62.520 ;
        RECT 1504.760 61.920 1505.020 62.180 ;
        RECT 1329.040 25.540 1329.300 25.800 ;
        RECT 1504.760 25.540 1505.020 25.800 ;
      LAYER met2 ;
        RECT 1508.430 1700.410 1508.710 1704.000 ;
        RECT 1507.580 1700.270 1508.710 1700.410 ;
        RECT 1507.580 1672.530 1507.720 1700.270 ;
        RECT 1508.430 1700.000 1508.710 1700.270 ;
        RECT 1507.120 1672.390 1507.720 1672.530 ;
        RECT 1507.120 1642.530 1507.260 1672.390 ;
        RECT 1505.680 1642.210 1505.940 1642.530 ;
        RECT 1507.060 1642.210 1507.320 1642.530 ;
        RECT 1505.740 1366.110 1505.880 1642.210 ;
        RECT 1505.680 1365.790 1505.940 1366.110 ;
        RECT 1505.680 1338.590 1505.940 1338.910 ;
        RECT 1505.740 1257.990 1505.880 1338.590 ;
        RECT 1505.680 1257.670 1505.940 1257.990 ;
        RECT 1505.680 1256.990 1505.940 1257.310 ;
        RECT 1505.740 1076.850 1505.880 1256.990 ;
        RECT 1505.280 1076.710 1505.880 1076.850 ;
        RECT 1505.280 1076.170 1505.420 1076.710 ;
        RECT 1505.280 1076.030 1505.880 1076.170 ;
        RECT 1505.740 886.710 1505.880 1076.030 ;
        RECT 1504.760 886.390 1505.020 886.710 ;
        RECT 1505.680 886.390 1505.940 886.710 ;
        RECT 1504.820 862.765 1504.960 886.390 ;
        RECT 1504.750 862.395 1505.030 862.765 ;
        RECT 1505.670 862.395 1505.950 862.765 ;
        RECT 1505.740 814.290 1505.880 862.395 ;
        RECT 1505.680 813.970 1505.940 814.290 ;
        RECT 1505.680 766.030 1505.940 766.350 ;
        RECT 1505.740 749.090 1505.880 766.030 ;
        RECT 1505.740 748.950 1506.800 749.090 ;
        RECT 1506.660 724.610 1506.800 748.950 ;
        RECT 1506.200 724.470 1506.800 724.610 ;
        RECT 1506.200 676.590 1506.340 724.470 ;
        RECT 1506.140 676.270 1506.400 676.590 ;
        RECT 1506.600 675.590 1506.860 675.910 ;
        RECT 1506.660 628.165 1506.800 675.590 ;
        RECT 1505.670 627.795 1505.950 628.165 ;
        RECT 1506.590 627.795 1506.870 628.165 ;
        RECT 1505.740 593.630 1505.880 627.795 ;
        RECT 1505.680 593.310 1505.940 593.630 ;
        RECT 1505.680 592.630 1505.940 592.950 ;
        RECT 1505.740 303.690 1505.880 592.630 ;
        RECT 1505.280 303.550 1505.880 303.690 ;
        RECT 1505.280 303.010 1505.420 303.550 ;
        RECT 1505.280 302.870 1505.880 303.010 ;
        RECT 1505.740 207.130 1505.880 302.870 ;
        RECT 1505.280 206.990 1505.880 207.130 ;
        RECT 1505.280 206.450 1505.420 206.990 ;
        RECT 1505.280 206.310 1505.880 206.450 ;
        RECT 1505.740 110.570 1505.880 206.310 ;
        RECT 1505.280 110.430 1505.880 110.570 ;
        RECT 1505.280 62.550 1505.420 110.430 ;
        RECT 1505.220 62.230 1505.480 62.550 ;
        RECT 1504.760 61.890 1505.020 62.210 ;
        RECT 1504.820 25.830 1504.960 61.890 ;
        RECT 1329.040 25.510 1329.300 25.830 ;
        RECT 1504.760 25.510 1505.020 25.830 ;
        RECT 1329.100 2.400 1329.240 25.510 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
      LAYER via2 ;
        RECT 1504.750 862.440 1505.030 862.720 ;
        RECT 1505.670 862.440 1505.950 862.720 ;
        RECT 1505.670 627.840 1505.950 628.120 ;
        RECT 1506.590 627.840 1506.870 628.120 ;
      LAYER met3 ;
        RECT 1504.725 862.730 1505.055 862.745 ;
        RECT 1505.645 862.730 1505.975 862.745 ;
        RECT 1504.725 862.430 1505.975 862.730 ;
        RECT 1504.725 862.415 1505.055 862.430 ;
        RECT 1505.645 862.415 1505.975 862.430 ;
        RECT 1505.645 628.130 1505.975 628.145 ;
        RECT 1506.565 628.130 1506.895 628.145 ;
        RECT 1505.645 627.830 1506.895 628.130 ;
        RECT 1505.645 627.815 1505.975 627.830 ;
        RECT 1506.565 627.815 1506.895 627.830 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1504.730 1678.140 1505.050 1678.200 ;
        RECT 1508.870 1678.140 1509.190 1678.200 ;
        RECT 1504.730 1678.000 1509.190 1678.140 ;
        RECT 1504.730 1677.940 1505.050 1678.000 ;
        RECT 1508.870 1677.940 1509.190 1678.000 ;
        RECT 1329.010 26.420 1329.330 26.480 ;
        RECT 1504.730 26.420 1505.050 26.480 ;
        RECT 1329.010 26.280 1505.050 26.420 ;
        RECT 1329.010 26.220 1329.330 26.280 ;
        RECT 1504.730 26.220 1505.050 26.280 ;
      LAYER via ;
        RECT 1504.760 1677.940 1505.020 1678.200 ;
        RECT 1508.900 1677.940 1509.160 1678.200 ;
        RECT 1329.040 26.220 1329.300 26.480 ;
        RECT 1504.760 26.220 1505.020 26.480 ;
      LAYER met2 ;
        RECT 1509.810 1700.410 1510.090 1704.000 ;
        RECT 1508.960 1700.270 1510.090 1700.410 ;
        RECT 1508.960 1678.230 1509.100 1700.270 ;
        RECT 1509.810 1700.000 1510.090 1700.270 ;
        RECT 1504.760 1677.910 1505.020 1678.230 ;
        RECT 1508.900 1677.910 1509.160 1678.230 ;
        RECT 1504.820 26.510 1504.960 1677.910 ;
        RECT 1329.040 26.190 1329.300 26.510 ;
        RECT 1504.760 26.190 1505.020 26.510 ;
        RECT 1329.100 2.400 1329.240 26.190 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 0.300 ;
=======
      LAYER met1 ;
        RECT 689.610 1625.100 689.930 1625.160 ;
        RECT 1333.150 1625.100 1333.470 1625.160 ;
        RECT 689.610 1624.960 1333.470 1625.100 ;
        RECT 689.610 1624.900 689.930 1624.960 ;
        RECT 1333.150 1624.900 1333.470 1624.960 ;
        RECT 686.390 2.960 686.710 3.020 ;
        RECT 689.610 2.960 689.930 3.020 ;
        RECT 686.390 2.820 689.930 2.960 ;
        RECT 686.390 2.760 686.710 2.820 ;
        RECT 689.610 2.760 689.930 2.820 ;
      LAYER via ;
        RECT 689.640 1624.900 689.900 1625.160 ;
        RECT 1333.180 1624.900 1333.440 1625.160 ;
        RECT 686.420 2.760 686.680 3.020 ;
        RECT 689.640 2.760 689.900 3.020 ;
      LAYER met2 ;
        RECT 1335.930 1700.410 1336.210 1704.000 ;
        RECT 1334.620 1700.270 1336.210 1700.410 ;
        RECT 1334.620 1677.290 1334.760 1700.270 ;
        RECT 1335.930 1700.000 1336.210 1700.270 ;
        RECT 1333.240 1677.150 1334.760 1677.290 ;
        RECT 1333.240 1625.190 1333.380 1677.150 ;
        RECT 689.640 1624.870 689.900 1625.190 ;
        RECT 1333.180 1624.870 1333.440 1625.190 ;
        RECT 689.700 3.050 689.840 1624.870 ;
        RECT 686.420 2.730 686.680 3.050 ;
        RECT 689.640 2.730 689.900 3.050 ;
        RECT 686.480 2.400 686.620 2.730 ;
        RECT 686.270 -4.800 686.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1346.490 26.760 1346.810 26.820 ;
        RECT 1513.470 26.760 1513.790 26.820 ;
        RECT 1346.490 26.620 1513.790 26.760 ;
        RECT 1346.490 26.560 1346.810 26.620 ;
        RECT 1513.470 26.560 1513.790 26.620 ;
      LAYER via ;
        RECT 1346.520 26.560 1346.780 26.820 ;
        RECT 1513.500 26.560 1513.760 26.820 ;
      LAYER met2 ;
        RECT 1514.870 1700.410 1515.150 1704.000 ;
        RECT 1513.560 1700.270 1515.150 1700.410 ;
        RECT 1513.560 26.850 1513.700 1700.270 ;
        RECT 1514.870 1700.000 1515.150 1700.270 ;
        RECT 1346.520 26.530 1346.780 26.850 ;
        RECT 1513.500 26.530 1513.760 26.850 ;
        RECT 1346.580 2.400 1346.720 26.530 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 0.300 ;
=======
      LAYER li1 ;
        RECT 1486.865 1686.825 1487.035 1690.395 ;
      LAYER mcon ;
        RECT 1486.865 1690.225 1487.035 1690.395 ;
      LAYER met1 ;
        RECT 1369.490 1690.380 1369.810 1690.440 ;
        RECT 1486.805 1690.380 1487.095 1690.425 ;
        RECT 1369.490 1690.240 1487.095 1690.380 ;
        RECT 1369.490 1690.180 1369.810 1690.240 ;
        RECT 1486.805 1690.195 1487.095 1690.240 ;
        RECT 1486.805 1686.980 1487.095 1687.025 ;
        RECT 1518.070 1686.980 1518.390 1687.040 ;
        RECT 1486.805 1686.840 1518.390 1686.980 ;
        RECT 1486.805 1686.795 1487.095 1686.840 ;
        RECT 1518.070 1686.780 1518.390 1686.840 ;
=======
      LAYER met1 ;
        RECT 1370.410 1688.340 1370.730 1688.400 ;
        RECT 1519.450 1688.340 1519.770 1688.400 ;
        RECT 1370.410 1688.200 1519.770 1688.340 ;
        RECT 1370.410 1688.140 1370.730 1688.200 ;
        RECT 1519.450 1688.140 1519.770 1688.200 ;
>>>>>>> re-updated local openlane
        RECT 1364.430 16.900 1364.750 16.960 ;
        RECT 1369.490 16.900 1369.810 16.960 ;
        RECT 1364.430 16.760 1369.810 16.900 ;
        RECT 1364.430 16.700 1364.750 16.760 ;
        RECT 1369.490 16.700 1369.810 16.760 ;
      LAYER via ;
        RECT 1370.440 1688.140 1370.700 1688.400 ;
        RECT 1519.480 1688.140 1519.740 1688.400 ;
        RECT 1364.460 16.700 1364.720 16.960 ;
        RECT 1369.520 16.700 1369.780 16.960 ;
      LAYER met2 ;
        RECT 1519.470 1700.000 1519.750 1704.000 ;
        RECT 1519.540 1688.430 1519.680 1700.000 ;
        RECT 1370.440 1688.110 1370.700 1688.430 ;
        RECT 1519.480 1688.110 1519.740 1688.430 ;
        RECT 1370.500 1672.530 1370.640 1688.110 ;
        RECT 1369.580 1672.390 1370.640 1672.530 ;
        RECT 1369.580 16.990 1369.720 1672.390 ;
        RECT 1364.460 16.670 1364.720 16.990 ;
        RECT 1369.520 16.670 1369.780 16.990 ;
        RECT 1364.520 2.400 1364.660 16.670 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 0.300 ;
=======
      LAYER li1 ;
        RECT 1438.565 1684.785 1438.735 1686.655 ;
      LAYER mcon ;
        RECT 1438.565 1686.485 1438.735 1686.655 ;
=======
>>>>>>> re-updated local openlane
      LAYER met1 ;
        RECT 1514.850 1683.920 1515.170 1683.980 ;
        RECT 1524.510 1683.920 1524.830 1683.980 ;
        RECT 1514.850 1683.780 1524.830 1683.920 ;
        RECT 1514.850 1683.720 1515.170 1683.780 ;
        RECT 1524.510 1683.720 1524.830 1683.780 ;
        RECT 1386.510 72.320 1386.830 72.380 ;
        RECT 1514.850 72.320 1515.170 72.380 ;
        RECT 1386.510 72.180 1515.170 72.320 ;
        RECT 1386.510 72.120 1386.830 72.180 ;
        RECT 1514.850 72.120 1515.170 72.180 ;
        RECT 1382.370 16.560 1382.690 16.620 ;
        RECT 1386.510 16.560 1386.830 16.620 ;
        RECT 1382.370 16.420 1386.830 16.560 ;
        RECT 1382.370 16.360 1382.690 16.420 ;
        RECT 1386.510 16.360 1386.830 16.420 ;
      LAYER via ;
        RECT 1514.880 1683.720 1515.140 1683.980 ;
        RECT 1524.540 1683.720 1524.800 1683.980 ;
        RECT 1386.540 72.120 1386.800 72.380 ;
        RECT 1514.880 72.120 1515.140 72.380 ;
        RECT 1382.400 16.360 1382.660 16.620 ;
        RECT 1386.540 16.360 1386.800 16.620 ;
      LAYER met2 ;
        RECT 1524.530 1700.000 1524.810 1704.000 ;
        RECT 1524.600 1684.010 1524.740 1700.000 ;
        RECT 1514.880 1683.690 1515.140 1684.010 ;
        RECT 1524.540 1683.690 1524.800 1684.010 ;
        RECT 1514.940 72.410 1515.080 1683.690 ;
        RECT 1386.540 72.090 1386.800 72.410 ;
        RECT 1514.880 72.090 1515.140 72.410 ;
        RECT 1386.600 16.650 1386.740 72.090 ;
        RECT 1382.400 16.330 1382.660 16.650 ;
        RECT 1386.540 16.330 1386.800 16.650 ;
        RECT 1382.460 2.400 1382.600 16.330 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 0.300 ;
=======
      LAYER li1 ;
        RECT 1459.265 16.065 1462.655 16.235 ;
        RECT 1465.245 16.065 1465.415 17.935 ;
        RECT 1508.025 17.765 1508.195 19.635 ;
        RECT 1437.645 14.535 1437.815 15.555 ;
        RECT 1437.645 14.365 1439.655 14.535 ;
        RECT 1459.265 14.365 1459.435 16.065 ;
      LAYER mcon ;
        RECT 1508.025 19.465 1508.195 19.635 ;
        RECT 1465.245 17.765 1465.415 17.935 ;
        RECT 1462.485 16.065 1462.655 16.235 ;
        RECT 1437.645 15.385 1437.815 15.555 ;
        RECT 1439.485 14.365 1439.655 14.535 ;
      LAYER met1 ;
        RECT 1526.810 19.960 1527.130 20.020 ;
        RECT 1518.620 19.820 1527.130 19.960 ;
        RECT 1507.965 19.620 1508.255 19.665 ;
        RECT 1518.620 19.620 1518.760 19.820 ;
        RECT 1526.810 19.760 1527.130 19.820 ;
        RECT 1507.965 19.480 1518.760 19.620 ;
        RECT 1507.965 19.435 1508.255 19.480 ;
        RECT 1465.185 17.920 1465.475 17.965 ;
        RECT 1507.965 17.920 1508.255 17.965 ;
        RECT 1465.185 17.780 1508.255 17.920 ;
        RECT 1465.185 17.735 1465.475 17.780 ;
        RECT 1507.965 17.735 1508.255 17.780 ;
        RECT 1462.425 16.220 1462.715 16.265 ;
        RECT 1465.185 16.220 1465.475 16.265 ;
        RECT 1462.425 16.080 1465.475 16.220 ;
        RECT 1462.425 16.035 1462.715 16.080 ;
        RECT 1465.185 16.035 1465.475 16.080 ;
        RECT 1400.310 15.540 1400.630 15.600 ;
        RECT 1437.585 15.540 1437.875 15.585 ;
        RECT 1400.310 15.400 1437.875 15.540 ;
        RECT 1400.310 15.340 1400.630 15.400 ;
        RECT 1437.585 15.355 1437.875 15.400 ;
        RECT 1439.425 14.520 1439.715 14.565 ;
        RECT 1459.205 14.520 1459.495 14.565 ;
        RECT 1439.425 14.380 1459.495 14.520 ;
        RECT 1439.425 14.335 1439.715 14.380 ;
        RECT 1459.205 14.335 1459.495 14.380 ;
      LAYER via ;
        RECT 1526.840 19.760 1527.100 20.020 ;
        RECT 1400.340 15.340 1400.600 15.600 ;
      LAYER met2 ;
        RECT 1527.750 1700.410 1528.030 1704.000 ;
        RECT 1526.900 1700.270 1528.030 1700.410 ;
        RECT 1526.900 20.050 1527.040 1700.270 ;
        RECT 1527.750 1700.000 1528.030 1700.270 ;
        RECT 1526.840 19.730 1527.100 20.050 ;
        RECT 1400.340 15.310 1400.600 15.630 ;
        RECT 1400.400 2.400 1400.540 15.310 ;
=======
      LAYER met1 ;
        RECT 1399.850 65.520 1400.170 65.580 ;
        RECT 1525.430 65.520 1525.750 65.580 ;
        RECT 1399.850 65.380 1525.750 65.520 ;
        RECT 1399.850 65.320 1400.170 65.380 ;
        RECT 1525.430 65.320 1525.750 65.380 ;
      LAYER via ;
        RECT 1399.880 65.320 1400.140 65.580 ;
        RECT 1525.460 65.320 1525.720 65.580 ;
      LAYER met2 ;
        RECT 1529.130 1700.410 1529.410 1704.000 ;
        RECT 1528.280 1700.270 1529.410 1700.410 ;
        RECT 1528.280 1679.330 1528.420 1700.270 ;
        RECT 1529.130 1700.000 1529.410 1700.270 ;
        RECT 1525.520 1679.190 1528.420 1679.330 ;
        RECT 1525.520 65.610 1525.660 1679.190 ;
        RECT 1399.880 65.290 1400.140 65.610 ;
        RECT 1525.460 65.290 1525.720 65.610 ;
        RECT 1399.940 20.130 1400.080 65.290 ;
        RECT 1399.940 19.990 1400.540 20.130 ;
        RECT 1400.400 2.400 1400.540 19.990 ;
>>>>>>> re-updated local openlane
        RECT 1400.190 -4.800 1400.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1452.750 1686.640 1453.070 1686.700 ;
        RECT 1534.170 1686.640 1534.490 1686.700 ;
        RECT 1452.750 1686.500 1534.490 1686.640 ;
        RECT 1452.750 1686.440 1453.070 1686.500 ;
        RECT 1534.170 1686.440 1534.490 1686.500 ;
        RECT 1418.250 20.640 1418.570 20.700 ;
        RECT 1452.290 20.640 1452.610 20.700 ;
        RECT 1418.250 20.500 1452.610 20.640 ;
        RECT 1418.250 20.440 1418.570 20.500 ;
        RECT 1452.290 20.440 1452.610 20.500 ;
      LAYER via ;
        RECT 1452.780 1686.440 1453.040 1686.700 ;
        RECT 1534.200 1686.440 1534.460 1686.700 ;
        RECT 1418.280 20.440 1418.540 20.700 ;
        RECT 1452.320 20.440 1452.580 20.700 ;
      LAYER met2 ;
        RECT 1534.190 1700.000 1534.470 1704.000 ;
        RECT 1534.260 1686.730 1534.400 1700.000 ;
        RECT 1452.780 1686.410 1453.040 1686.730 ;
        RECT 1534.200 1686.410 1534.460 1686.730 ;
        RECT 1452.840 1671.170 1452.980 1686.410 ;
        RECT 1452.380 1671.030 1452.980 1671.170 ;
        RECT 1452.380 20.730 1452.520 1671.030 ;
        RECT 1418.280 20.410 1418.540 20.730 ;
        RECT 1452.320 20.410 1452.580 20.730 ;
        RECT 1418.340 2.400 1418.480 20.410 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1486.790 1689.360 1487.110 1689.420 ;
        RECT 1538.770 1689.360 1539.090 1689.420 ;
        RECT 1486.790 1689.220 1539.090 1689.360 ;
        RECT 1486.790 1689.160 1487.110 1689.220 ;
        RECT 1538.770 1689.160 1539.090 1689.220 ;
        RECT 1435.730 14.860 1436.050 14.920 ;
        RECT 1435.730 14.720 1471.380 14.860 ;
        RECT 1435.730 14.660 1436.050 14.720 ;
        RECT 1471.240 14.520 1471.380 14.720 ;
        RECT 1484.950 14.520 1485.270 14.580 ;
        RECT 1471.240 14.380 1485.270 14.520 ;
        RECT 1484.950 14.320 1485.270 14.380 ;
      LAYER via ;
        RECT 1486.820 1689.160 1487.080 1689.420 ;
        RECT 1538.800 1689.160 1539.060 1689.420 ;
        RECT 1435.760 14.660 1436.020 14.920 ;
        RECT 1484.980 14.320 1485.240 14.580 ;
      LAYER met2 ;
        RECT 1538.790 1700.000 1539.070 1704.000 ;
        RECT 1538.860 1689.450 1539.000 1700.000 ;
        RECT 1486.820 1689.130 1487.080 1689.450 ;
        RECT 1538.800 1689.130 1539.060 1689.450 ;
        RECT 1486.880 24.890 1487.020 1689.130 ;
        RECT 1485.040 24.750 1487.020 24.890 ;
        RECT 1435.760 14.630 1436.020 14.950 ;
        RECT 1435.820 2.400 1435.960 14.630 ;
        RECT 1485.040 14.610 1485.180 24.750 ;
        RECT 1484.980 14.290 1485.240 14.610 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1539.690 1678.140 1540.010 1678.200 ;
        RECT 1542.450 1678.140 1542.770 1678.200 ;
        RECT 1539.690 1678.000 1542.770 1678.140 ;
        RECT 1539.690 1677.940 1540.010 1678.000 ;
        RECT 1542.450 1677.940 1542.770 1678.000 ;
        RECT 1539.690 16.560 1540.010 16.620 ;
        RECT 1486.880 16.420 1540.010 16.560 ;
        RECT 1453.670 16.220 1453.990 16.280 ;
        RECT 1486.880 16.220 1487.020 16.420 ;
        RECT 1539.690 16.360 1540.010 16.420 ;
        RECT 1453.670 16.080 1487.020 16.220 ;
        RECT 1453.670 16.020 1453.990 16.080 ;
      LAYER via ;
        RECT 1539.720 1677.940 1539.980 1678.200 ;
        RECT 1542.480 1677.940 1542.740 1678.200 ;
        RECT 1453.700 16.020 1453.960 16.280 ;
        RECT 1539.720 16.360 1539.980 16.620 ;
      LAYER met2 ;
        RECT 1543.850 1700.410 1544.130 1704.000 ;
        RECT 1542.540 1700.270 1544.130 1700.410 ;
        RECT 1542.540 1678.230 1542.680 1700.270 ;
        RECT 1543.850 1700.000 1544.130 1700.270 ;
        RECT 1539.720 1677.910 1539.980 1678.230 ;
        RECT 1542.480 1677.910 1542.740 1678.230 ;
        RECT 1539.780 16.650 1539.920 1677.910 ;
        RECT 1539.720 16.330 1539.980 16.650 ;
        RECT 1453.700 15.990 1453.960 16.310 ;
        RECT 1453.760 2.400 1453.900 15.990 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1507.950 1687.320 1508.270 1687.380 ;
        RECT 1547.050 1687.320 1547.370 1687.380 ;
        RECT 1507.950 1687.180 1547.370 1687.320 ;
        RECT 1507.950 1687.120 1508.270 1687.180 ;
        RECT 1547.050 1687.120 1547.370 1687.180 ;
        RECT 1471.610 19.620 1471.930 19.680 ;
        RECT 1507.490 19.620 1507.810 19.680 ;
        RECT 1471.610 19.480 1507.810 19.620 ;
        RECT 1471.610 19.420 1471.930 19.480 ;
        RECT 1507.490 19.420 1507.810 19.480 ;
      LAYER via ;
        RECT 1507.980 1687.120 1508.240 1687.380 ;
        RECT 1547.080 1687.120 1547.340 1687.380 ;
        RECT 1471.640 19.420 1471.900 19.680 ;
        RECT 1507.520 19.420 1507.780 19.680 ;
=======
      LAYER li1 ;
        RECT 1487.325 14.705 1487.495 16.235 ;
      LAYER mcon ;
        RECT 1487.325 16.065 1487.495 16.235 ;
      LAYER met1 ;
        RECT 1514.390 1684.940 1514.710 1685.000 ;
        RECT 1548.430 1684.940 1548.750 1685.000 ;
        RECT 1514.390 1684.800 1548.750 1684.940 ;
        RECT 1514.390 1684.740 1514.710 1684.800 ;
        RECT 1548.430 1684.740 1548.750 1684.800 ;
        RECT 1487.265 16.220 1487.555 16.265 ;
        RECT 1514.390 16.220 1514.710 16.280 ;
        RECT 1487.265 16.080 1514.710 16.220 ;
        RECT 1487.265 16.035 1487.555 16.080 ;
        RECT 1514.390 16.020 1514.710 16.080 ;
        RECT 1471.610 14.860 1471.930 14.920 ;
        RECT 1487.265 14.860 1487.555 14.905 ;
        RECT 1471.610 14.720 1487.555 14.860 ;
        RECT 1471.610 14.660 1471.930 14.720 ;
        RECT 1487.265 14.675 1487.555 14.720 ;
      LAYER via ;
        RECT 1514.420 1684.740 1514.680 1685.000 ;
        RECT 1548.460 1684.740 1548.720 1685.000 ;
        RECT 1514.420 16.020 1514.680 16.280 ;
        RECT 1471.640 14.660 1471.900 14.920 ;
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1548.450 1700.000 1548.730 1704.000 ;
        RECT 1548.520 1685.030 1548.660 1700.000 ;
        RECT 1514.420 1684.710 1514.680 1685.030 ;
        RECT 1548.460 1684.710 1548.720 1685.030 ;
        RECT 1514.480 16.310 1514.620 1684.710 ;
        RECT 1514.420 15.990 1514.680 16.310 ;
        RECT 1471.640 14.630 1471.900 14.950 ;
        RECT 1471.700 2.400 1471.840 14.630 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1521.290 1684.260 1521.610 1684.320 ;
        RECT 1553.490 1684.260 1553.810 1684.320 ;
        RECT 1521.290 1684.120 1553.810 1684.260 ;
        RECT 1521.290 1684.060 1521.610 1684.120 ;
        RECT 1553.490 1684.060 1553.810 1684.120 ;
        RECT 1489.550 14.520 1489.870 14.580 ;
        RECT 1521.290 14.520 1521.610 14.580 ;
        RECT 1489.550 14.380 1521.610 14.520 ;
        RECT 1489.550 14.320 1489.870 14.380 ;
        RECT 1521.290 14.320 1521.610 14.380 ;
      LAYER via ;
        RECT 1521.320 1684.060 1521.580 1684.320 ;
        RECT 1553.520 1684.060 1553.780 1684.320 ;
        RECT 1489.580 14.320 1489.840 14.580 ;
        RECT 1521.320 14.320 1521.580 14.580 ;
      LAYER met2 ;
        RECT 1553.510 1700.000 1553.790 1704.000 ;
        RECT 1553.580 1684.350 1553.720 1700.000 ;
        RECT 1521.320 1684.030 1521.580 1684.350 ;
        RECT 1553.520 1684.030 1553.780 1684.350 ;
        RECT 1521.380 14.610 1521.520 1684.030 ;
        RECT 1489.580 14.290 1489.840 14.610 ;
        RECT 1521.320 14.290 1521.580 14.610 ;
        RECT 1489.640 2.400 1489.780 14.290 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 0.300 ;
=======
      LAYER met1 ;
        RECT 1530.490 1683.920 1530.810 1683.980 ;
        RECT 1558.550 1683.920 1558.870 1683.980 ;
        RECT 1530.490 1683.780 1558.870 1683.920 ;
        RECT 1530.490 1683.720 1530.810 1683.780 ;
        RECT 1558.550 1683.720 1558.870 1683.780 ;
        RECT 1507.030 18.600 1507.350 18.660 ;
        RECT 1528.650 18.600 1528.970 18.660 ;
        RECT 1507.030 18.460 1528.970 18.600 ;
        RECT 1507.030 18.400 1507.350 18.460 ;
        RECT 1528.650 18.400 1528.970 18.460 ;
      LAYER via ;
        RECT 1530.520 1683.720 1530.780 1683.980 ;
        RECT 1558.580 1683.720 1558.840 1683.980 ;
        RECT 1507.060 18.400 1507.320 18.660 ;
        RECT 1528.680 18.400 1528.940 18.660 ;
      LAYER met2 ;
        RECT 1558.570 1700.000 1558.850 1704.000 ;
        RECT 1558.640 1684.010 1558.780 1700.000 ;
        RECT 1530.520 1683.690 1530.780 1684.010 ;
        RECT 1558.580 1683.690 1558.840 1684.010 ;
        RECT 1530.580 1671.170 1530.720 1683.690 ;
        RECT 1528.740 1671.030 1530.720 1671.170 ;
        RECT 1528.740 18.690 1528.880 1671.030 ;
        RECT 1507.060 18.370 1507.320 18.690 ;
        RECT 1528.680 18.370 1528.940 18.690 ;
        RECT 1507.120 2.400 1507.260 18.370 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 0.300 ;
=======
      LAYER met1 ;
        RECT 710.310 1639.040 710.630 1639.100 ;
        RECT 1340.050 1639.040 1340.370 1639.100 ;
        RECT 710.310 1638.900 1340.370 1639.040 ;
        RECT 710.310 1638.840 710.630 1638.900 ;
        RECT 1340.050 1638.840 1340.370 1638.900 ;
        RECT 704.330 20.980 704.650 21.040 ;
        RECT 710.310 20.980 710.630 21.040 ;
        RECT 704.330 20.840 710.630 20.980 ;
        RECT 704.330 20.780 704.650 20.840 ;
        RECT 710.310 20.780 710.630 20.840 ;
      LAYER via ;
        RECT 710.340 1638.840 710.600 1639.100 ;
        RECT 1340.080 1638.840 1340.340 1639.100 ;
        RECT 704.360 20.780 704.620 21.040 ;
        RECT 710.340 20.780 710.600 21.040 ;
      LAYER met2 ;
        RECT 1340.530 1700.410 1340.810 1704.000 ;
        RECT 1340.140 1700.270 1340.810 1700.410 ;
        RECT 1340.140 1639.130 1340.280 1700.270 ;
        RECT 1340.530 1700.000 1340.810 1700.270 ;
        RECT 710.340 1638.810 710.600 1639.130 ;
        RECT 1340.080 1638.810 1340.340 1639.130 ;
        RECT 710.400 21.070 710.540 1638.810 ;
        RECT 704.360 20.750 704.620 21.070 ;
        RECT 710.340 20.750 710.600 21.070 ;
        RECT 704.420 2.400 704.560 20.750 ;
        RECT 704.210 -4.800 704.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1541.990 1690.040 1542.310 1690.100 ;
        RECT 1563.150 1690.040 1563.470 1690.100 ;
        RECT 1541.990 1689.900 1563.470 1690.040 ;
        RECT 1541.990 1689.840 1542.310 1689.900 ;
        RECT 1563.150 1689.840 1563.470 1689.900 ;
        RECT 1524.970 15.200 1525.290 15.260 ;
        RECT 1541.990 15.200 1542.310 15.260 ;
        RECT 1524.970 15.060 1542.310 15.200 ;
        RECT 1524.970 15.000 1525.290 15.060 ;
        RECT 1541.990 15.000 1542.310 15.060 ;
      LAYER via ;
        RECT 1542.020 1689.840 1542.280 1690.100 ;
        RECT 1563.180 1689.840 1563.440 1690.100 ;
        RECT 1525.000 15.000 1525.260 15.260 ;
        RECT 1542.020 15.000 1542.280 15.260 ;
      LAYER met2 ;
        RECT 1563.170 1700.000 1563.450 1704.000 ;
        RECT 1563.240 1690.130 1563.380 1700.000 ;
        RECT 1542.020 1689.810 1542.280 1690.130 ;
        RECT 1563.180 1689.810 1563.440 1690.130 ;
        RECT 1542.080 15.290 1542.220 1689.810 ;
        RECT 1525.000 14.970 1525.260 15.290 ;
        RECT 1542.020 14.970 1542.280 15.290 ;
        RECT 1525.060 2.400 1525.200 14.970 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1545.210 1690.380 1545.530 1690.440 ;
        RECT 1568.210 1690.380 1568.530 1690.440 ;
        RECT 1545.210 1690.240 1568.530 1690.380 ;
        RECT 1545.210 1690.180 1545.530 1690.240 ;
        RECT 1568.210 1690.180 1568.530 1690.240 ;
        RECT 1542.910 20.640 1543.230 20.700 ;
        RECT 1545.210 20.640 1545.530 20.700 ;
        RECT 1542.910 20.500 1545.530 20.640 ;
        RECT 1542.910 20.440 1543.230 20.500 ;
        RECT 1545.210 20.440 1545.530 20.500 ;
      LAYER via ;
        RECT 1545.240 1690.180 1545.500 1690.440 ;
        RECT 1568.240 1690.180 1568.500 1690.440 ;
        RECT 1542.940 20.440 1543.200 20.700 ;
        RECT 1545.240 20.440 1545.500 20.700 ;
      LAYER met2 ;
        RECT 1568.230 1700.000 1568.510 1704.000 ;
        RECT 1568.300 1690.470 1568.440 1700.000 ;
        RECT 1545.240 1690.150 1545.500 1690.470 ;
        RECT 1568.240 1690.150 1568.500 1690.470 ;
        RECT 1545.300 20.730 1545.440 1690.150 ;
        RECT 1542.940 20.410 1543.200 20.730 ;
        RECT 1545.240 20.410 1545.500 20.730 ;
        RECT 1543.000 2.400 1543.140 20.410 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1565.910 1683.920 1566.230 1683.980 ;
        RECT 1572.810 1683.920 1573.130 1683.980 ;
        RECT 1565.910 1683.780 1573.130 1683.920 ;
        RECT 1565.910 1683.720 1566.230 1683.780 ;
        RECT 1572.810 1683.720 1573.130 1683.780 ;
        RECT 1560.850 20.640 1561.170 20.700 ;
        RECT 1565.910 20.640 1566.230 20.700 ;
        RECT 1560.850 20.500 1566.230 20.640 ;
        RECT 1560.850 20.440 1561.170 20.500 ;
        RECT 1565.910 20.440 1566.230 20.500 ;
      LAYER via ;
        RECT 1565.940 1683.720 1566.200 1683.980 ;
        RECT 1572.840 1683.720 1573.100 1683.980 ;
        RECT 1560.880 20.440 1561.140 20.700 ;
        RECT 1565.940 20.440 1566.200 20.700 ;
      LAYER met2 ;
        RECT 1572.830 1700.000 1573.110 1704.000 ;
        RECT 1572.900 1684.010 1573.040 1700.000 ;
        RECT 1565.940 1683.690 1566.200 1684.010 ;
        RECT 1572.840 1683.690 1573.100 1684.010 ;
        RECT 1566.000 20.730 1566.140 1683.690 ;
        RECT 1560.880 20.410 1561.140 20.730 ;
        RECT 1565.940 20.410 1566.200 20.730 ;
        RECT 1560.940 2.400 1561.080 20.410 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 0.300 ;
=======
      LAYER met1 ;
        RECT 1573.730 1678.140 1574.050 1678.200 ;
        RECT 1576.490 1678.140 1576.810 1678.200 ;
        RECT 1573.730 1678.000 1576.810 1678.140 ;
        RECT 1573.730 1677.940 1574.050 1678.000 ;
        RECT 1576.490 1677.940 1576.810 1678.000 ;
        RECT 1573.730 20.640 1574.050 20.700 ;
        RECT 1578.790 20.640 1579.110 20.700 ;
        RECT 1573.730 20.500 1579.110 20.640 ;
        RECT 1573.730 20.440 1574.050 20.500 ;
        RECT 1578.790 20.440 1579.110 20.500 ;
      LAYER via ;
        RECT 1573.760 1677.940 1574.020 1678.200 ;
        RECT 1576.520 1677.940 1576.780 1678.200 ;
        RECT 1573.760 20.440 1574.020 20.700 ;
        RECT 1578.820 20.440 1579.080 20.700 ;
      LAYER met2 ;
        RECT 1577.890 1700.410 1578.170 1704.000 ;
        RECT 1576.580 1700.270 1578.170 1700.410 ;
        RECT 1576.580 1678.230 1576.720 1700.270 ;
        RECT 1577.890 1700.000 1578.170 1700.270 ;
        RECT 1573.760 1677.910 1574.020 1678.230 ;
        RECT 1576.520 1677.910 1576.780 1678.230 ;
        RECT 1573.820 20.730 1573.960 1677.910 ;
        RECT 1573.760 20.410 1574.020 20.730 ;
        RECT 1578.820 20.410 1579.080 20.730 ;
        RECT 1578.880 2.400 1579.020 20.410 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 0.300 ;
=======
      LAYER met1 ;
        RECT 1582.470 1685.280 1582.790 1685.340 ;
        RECT 1594.430 1685.280 1594.750 1685.340 ;
        RECT 1582.470 1685.140 1594.750 1685.280 ;
        RECT 1582.470 1685.080 1582.790 1685.140 ;
        RECT 1594.430 1685.080 1594.750 1685.140 ;
        RECT 1593.970 2.960 1594.290 3.020 ;
        RECT 1596.270 2.960 1596.590 3.020 ;
        RECT 1593.970 2.820 1596.590 2.960 ;
        RECT 1593.970 2.760 1594.290 2.820 ;
        RECT 1596.270 2.760 1596.590 2.820 ;
      LAYER via ;
        RECT 1582.500 1685.080 1582.760 1685.340 ;
        RECT 1594.460 1685.080 1594.720 1685.340 ;
        RECT 1594.000 2.760 1594.260 3.020 ;
        RECT 1596.300 2.760 1596.560 3.020 ;
      LAYER met2 ;
        RECT 1582.490 1700.000 1582.770 1704.000 ;
        RECT 1582.560 1685.370 1582.700 1700.000 ;
        RECT 1582.500 1685.050 1582.760 1685.370 ;
        RECT 1594.460 1685.050 1594.720 1685.370 ;
        RECT 1594.520 1677.970 1594.660 1685.050 ;
        RECT 1594.060 1677.830 1594.660 1677.970 ;
        RECT 1594.060 3.050 1594.200 1677.830 ;
        RECT 1594.000 2.730 1594.260 3.050 ;
        RECT 1596.300 2.730 1596.560 3.050 ;
        RECT 1596.360 2.400 1596.500 2.730 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1587.530 1684.260 1587.850 1684.320 ;
        RECT 1597.650 1684.260 1597.970 1684.320 ;
        RECT 1587.530 1684.120 1597.970 1684.260 ;
        RECT 1587.530 1684.060 1587.850 1684.120 ;
        RECT 1597.650 1684.060 1597.970 1684.120 ;
        RECT 1597.650 17.580 1597.970 17.640 ;
        RECT 1614.210 17.580 1614.530 17.640 ;
        RECT 1597.650 17.440 1614.530 17.580 ;
        RECT 1597.650 17.380 1597.970 17.440 ;
        RECT 1614.210 17.380 1614.530 17.440 ;
      LAYER via ;
        RECT 1587.560 1684.060 1587.820 1684.320 ;
        RECT 1597.680 1684.060 1597.940 1684.320 ;
        RECT 1597.680 17.380 1597.940 17.640 ;
        RECT 1614.240 17.380 1614.500 17.640 ;
      LAYER met2 ;
        RECT 1587.550 1700.000 1587.830 1704.000 ;
        RECT 1587.620 1684.350 1587.760 1700.000 ;
        RECT 1587.560 1684.030 1587.820 1684.350 ;
        RECT 1597.680 1684.030 1597.940 1684.350 ;
        RECT 1597.740 17.670 1597.880 1684.030 ;
        RECT 1597.680 17.350 1597.940 17.670 ;
        RECT 1614.240 17.350 1614.500 17.670 ;
        RECT 1614.300 2.400 1614.440 17.350 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1592.130 1685.960 1592.450 1686.020 ;
        RECT 1604.550 1685.960 1604.870 1686.020 ;
        RECT 1592.130 1685.820 1604.870 1685.960 ;
        RECT 1592.130 1685.760 1592.450 1685.820 ;
        RECT 1604.550 1685.760 1604.870 1685.820 ;
        RECT 1604.550 20.300 1604.870 20.360 ;
        RECT 1632.150 20.300 1632.470 20.360 ;
        RECT 1604.550 20.160 1632.470 20.300 ;
        RECT 1604.550 20.100 1604.870 20.160 ;
        RECT 1632.150 20.100 1632.470 20.160 ;
      LAYER via ;
        RECT 1592.160 1685.760 1592.420 1686.020 ;
        RECT 1604.580 1685.760 1604.840 1686.020 ;
        RECT 1604.580 20.100 1604.840 20.360 ;
        RECT 1632.180 20.100 1632.440 20.360 ;
      LAYER met2 ;
        RECT 1592.150 1700.000 1592.430 1704.000 ;
        RECT 1592.220 1686.050 1592.360 1700.000 ;
        RECT 1592.160 1685.730 1592.420 1686.050 ;
        RECT 1604.580 1685.730 1604.840 1686.050 ;
        RECT 1604.640 20.390 1604.780 1685.730 ;
        RECT 1604.580 20.070 1604.840 20.390 ;
        RECT 1632.180 20.070 1632.440 20.390 ;
        RECT 1632.240 2.400 1632.380 20.070 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1597.190 1686.300 1597.510 1686.360 ;
        RECT 1610.990 1686.300 1611.310 1686.360 ;
        RECT 1597.190 1686.160 1611.310 1686.300 ;
        RECT 1597.190 1686.100 1597.510 1686.160 ;
        RECT 1610.990 1686.100 1611.310 1686.160 ;
        RECT 1610.990 16.900 1611.310 16.960 ;
        RECT 1650.090 16.900 1650.410 16.960 ;
        RECT 1610.990 16.760 1650.410 16.900 ;
        RECT 1610.990 16.700 1611.310 16.760 ;
        RECT 1650.090 16.700 1650.410 16.760 ;
      LAYER via ;
        RECT 1597.220 1686.100 1597.480 1686.360 ;
        RECT 1611.020 1686.100 1611.280 1686.360 ;
        RECT 1611.020 16.700 1611.280 16.960 ;
        RECT 1650.120 16.700 1650.380 16.960 ;
      LAYER met2 ;
        RECT 1597.210 1700.000 1597.490 1704.000 ;
        RECT 1597.280 1686.390 1597.420 1700.000 ;
        RECT 1597.220 1686.070 1597.480 1686.390 ;
        RECT 1611.020 1686.070 1611.280 1686.390 ;
        RECT 1611.080 16.990 1611.220 1686.070 ;
        RECT 1611.020 16.670 1611.280 16.990 ;
        RECT 1650.120 16.670 1650.380 16.990 ;
        RECT 1650.180 2.400 1650.320 16.670 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 0.300 ;
=======
      LAYER met1 ;
        RECT 1601.790 1684.260 1602.110 1684.320 ;
        RECT 1607.310 1684.260 1607.630 1684.320 ;
        RECT 1601.790 1684.120 1607.630 1684.260 ;
        RECT 1601.790 1684.060 1602.110 1684.120 ;
        RECT 1607.310 1684.060 1607.630 1684.120 ;
        RECT 1607.310 18.260 1607.630 18.320 ;
        RECT 1607.310 18.120 1631.920 18.260 ;
        RECT 1607.310 18.060 1607.630 18.120 ;
        RECT 1631.780 17.580 1631.920 18.120 ;
        RECT 1668.030 17.580 1668.350 17.640 ;
        RECT 1631.780 17.440 1668.350 17.580 ;
        RECT 1668.030 17.380 1668.350 17.440 ;
      LAYER via ;
        RECT 1601.820 1684.060 1602.080 1684.320 ;
        RECT 1607.340 1684.060 1607.600 1684.320 ;
        RECT 1607.340 18.060 1607.600 18.320 ;
        RECT 1668.060 17.380 1668.320 17.640 ;
      LAYER met2 ;
        RECT 1601.810 1700.000 1602.090 1704.000 ;
        RECT 1601.880 1684.350 1602.020 1700.000 ;
        RECT 1601.820 1684.030 1602.080 1684.350 ;
        RECT 1607.340 1684.030 1607.600 1684.350 ;
        RECT 1607.400 18.350 1607.540 1684.030 ;
        RECT 1607.340 18.030 1607.600 18.350 ;
        RECT 1668.060 17.350 1668.320 17.670 ;
        RECT 1668.120 2.400 1668.260 17.350 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 0.300 ;
=======
      LAYER li1 ;
        RECT 1674.085 17.425 1674.255 20.315 ;
      LAYER mcon ;
        RECT 1674.085 20.145 1674.255 20.315 ;
=======
>>>>>>> re-updated local openlane
      LAYER met1 ;
        RECT 1607.310 1687.660 1607.630 1687.720 ;
        RECT 1685.510 1687.660 1685.830 1687.720 ;
        RECT 1607.310 1687.520 1685.830 1687.660 ;
        RECT 1607.310 1687.460 1607.630 1687.520 ;
        RECT 1685.510 1687.460 1685.830 1687.520 ;
      LAYER via ;
        RECT 1607.340 1687.460 1607.600 1687.720 ;
        RECT 1685.540 1687.460 1685.800 1687.720 ;
      LAYER met2 ;
        RECT 1606.870 1700.410 1607.150 1704.000 ;
        RECT 1606.870 1700.270 1607.540 1700.410 ;
        RECT 1606.870 1700.000 1607.150 1700.270 ;
        RECT 1607.400 1687.750 1607.540 1700.270 ;
        RECT 1607.340 1687.430 1607.600 1687.750 ;
        RECT 1685.540 1687.430 1685.800 1687.750 ;
        RECT 1685.600 2.400 1685.740 1687.430 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 0.300 ;
=======
      LAYER li1 ;
        RECT 1340.585 1580.065 1340.755 1594.515 ;
        RECT 1340.585 1435.225 1340.755 1442.195 ;
        RECT 1340.585 565.845 1340.755 613.275 ;
        RECT 1341.045 421.345 1341.215 475.915 ;
        RECT 1341.045 324.785 1341.215 372.555 ;
        RECT 1341.045 276.165 1341.215 324.275 ;
      LAYER mcon ;
        RECT 1340.585 1594.345 1340.755 1594.515 ;
        RECT 1340.585 1442.025 1340.755 1442.195 ;
        RECT 1340.585 613.105 1340.755 613.275 ;
        RECT 1341.045 475.745 1341.215 475.915 ;
        RECT 1341.045 372.385 1341.215 372.555 ;
        RECT 1341.045 324.105 1341.215 324.275 ;
      LAYER met1 ;
        RECT 1341.430 1666.580 1341.750 1666.640 ;
        RECT 1344.190 1666.580 1344.510 1666.640 ;
        RECT 1341.430 1666.440 1344.510 1666.580 ;
        RECT 1341.430 1666.380 1341.750 1666.440 ;
        RECT 1344.190 1666.380 1344.510 1666.440 ;
        RECT 1340.525 1594.500 1340.815 1594.545 ;
        RECT 1341.430 1594.500 1341.750 1594.560 ;
        RECT 1340.525 1594.360 1341.750 1594.500 ;
        RECT 1340.525 1594.315 1340.815 1594.360 ;
        RECT 1341.430 1594.300 1341.750 1594.360 ;
        RECT 1340.510 1580.220 1340.830 1580.280 ;
        RECT 1340.315 1580.080 1340.830 1580.220 ;
        RECT 1340.510 1580.020 1340.830 1580.080 ;
        RECT 1340.525 1442.180 1340.815 1442.225 ;
        RECT 1340.970 1442.180 1341.290 1442.240 ;
        RECT 1340.525 1442.040 1341.290 1442.180 ;
        RECT 1340.525 1441.995 1340.815 1442.040 ;
        RECT 1340.970 1441.980 1341.290 1442.040 ;
        RECT 1340.510 1435.380 1340.830 1435.440 ;
        RECT 1340.315 1435.240 1340.830 1435.380 ;
        RECT 1340.510 1435.180 1340.830 1435.240 ;
        RECT 1340.510 1076.480 1340.830 1076.740 ;
        RECT 1340.600 1076.340 1340.740 1076.480 ;
        RECT 1340.970 1076.340 1341.290 1076.400 ;
        RECT 1340.600 1076.200 1341.290 1076.340 ;
        RECT 1340.970 1076.140 1341.290 1076.200 ;
        RECT 1340.510 917.900 1340.830 917.960 ;
        RECT 1341.430 917.900 1341.750 917.960 ;
        RECT 1340.510 917.760 1341.750 917.900 ;
        RECT 1340.510 917.700 1340.830 917.760 ;
        RECT 1341.430 917.700 1341.750 917.760 ;
        RECT 1340.510 613.740 1340.830 614.000 ;
        RECT 1340.600 613.305 1340.740 613.740 ;
        RECT 1340.525 613.075 1340.815 613.305 ;
        RECT 1340.510 566.000 1340.830 566.060 ;
        RECT 1340.315 565.860 1340.830 566.000 ;
        RECT 1340.510 565.800 1340.830 565.860 ;
        RECT 1340.970 475.900 1341.290 475.960 ;
        RECT 1340.775 475.760 1341.290 475.900 ;
        RECT 1340.970 475.700 1341.290 475.760 ;
        RECT 1340.510 421.500 1340.830 421.560 ;
        RECT 1340.985 421.500 1341.275 421.545 ;
        RECT 1340.510 421.360 1341.275 421.500 ;
        RECT 1340.510 421.300 1340.830 421.360 ;
        RECT 1340.985 421.315 1341.275 421.360 ;
        RECT 1340.510 420.820 1340.830 420.880 ;
        RECT 1341.430 420.820 1341.750 420.880 ;
        RECT 1340.510 420.680 1341.750 420.820 ;
        RECT 1340.510 420.620 1340.830 420.680 ;
        RECT 1341.430 420.620 1341.750 420.680 ;
        RECT 1340.970 372.540 1341.290 372.600 ;
        RECT 1340.775 372.400 1341.290 372.540 ;
        RECT 1340.970 372.340 1341.290 372.400 ;
        RECT 1340.970 324.940 1341.290 325.000 ;
        RECT 1340.775 324.800 1341.290 324.940 ;
        RECT 1340.970 324.740 1341.290 324.800 ;
        RECT 1340.970 324.260 1341.290 324.320 ;
        RECT 1340.775 324.120 1341.290 324.260 ;
        RECT 1340.970 324.060 1341.290 324.120 ;
        RECT 1340.985 276.320 1341.275 276.365 ;
        RECT 1341.430 276.320 1341.750 276.380 ;
        RECT 1340.985 276.180 1341.750 276.320 ;
        RECT 1340.985 276.135 1341.275 276.180 ;
        RECT 1341.430 276.120 1341.750 276.180 ;
        RECT 1340.970 234.840 1341.290 234.900 ;
        RECT 1340.600 234.700 1341.290 234.840 ;
        RECT 1340.600 234.220 1340.740 234.700 ;
        RECT 1340.970 234.640 1341.290 234.700 ;
        RECT 1340.510 233.960 1340.830 234.220 ;
        RECT 724.110 51.240 724.430 51.300 ;
        RECT 1340.510 51.240 1340.830 51.300 ;
        RECT 724.110 51.100 1340.830 51.240 ;
        RECT 724.110 51.040 724.430 51.100 ;
        RECT 1340.510 51.040 1340.830 51.100 ;
      LAYER via ;
        RECT 1341.460 1666.380 1341.720 1666.640 ;
        RECT 1344.220 1666.380 1344.480 1666.640 ;
        RECT 1341.460 1594.300 1341.720 1594.560 ;
        RECT 1340.540 1580.020 1340.800 1580.280 ;
        RECT 1341.000 1441.980 1341.260 1442.240 ;
        RECT 1340.540 1435.180 1340.800 1435.440 ;
        RECT 1340.540 1076.480 1340.800 1076.740 ;
        RECT 1341.000 1076.140 1341.260 1076.400 ;
        RECT 1340.540 917.700 1340.800 917.960 ;
        RECT 1341.460 917.700 1341.720 917.960 ;
        RECT 1340.540 613.740 1340.800 614.000 ;
        RECT 1340.540 565.800 1340.800 566.060 ;
        RECT 1341.000 475.700 1341.260 475.960 ;
        RECT 1340.540 421.300 1340.800 421.560 ;
        RECT 1340.540 420.620 1340.800 420.880 ;
        RECT 1341.460 420.620 1341.720 420.880 ;
        RECT 1341.000 372.340 1341.260 372.600 ;
        RECT 1341.000 324.740 1341.260 325.000 ;
        RECT 1341.000 324.060 1341.260 324.320 ;
        RECT 1341.460 276.120 1341.720 276.380 ;
        RECT 1341.000 234.640 1341.260 234.900 ;
        RECT 1340.540 233.960 1340.800 234.220 ;
        RECT 724.140 51.040 724.400 51.300 ;
        RECT 1340.540 51.040 1340.800 51.300 ;
      LAYER met2 ;
        RECT 1344.670 1700.410 1344.950 1704.000 ;
        RECT 1344.280 1700.270 1344.950 1700.410 ;
        RECT 1344.280 1666.670 1344.420 1700.270 ;
        RECT 1344.670 1700.000 1344.950 1700.270 ;
        RECT 1341.460 1666.350 1341.720 1666.670 ;
        RECT 1344.220 1666.350 1344.480 1666.670 ;
        RECT 1341.520 1594.590 1341.660 1666.350 ;
        RECT 1341.460 1594.270 1341.720 1594.590 ;
        RECT 1340.540 1580.165 1340.800 1580.310 ;
        RECT 1340.530 1579.795 1340.810 1580.165 ;
        RECT 1340.990 1537.635 1341.270 1538.005 ;
        RECT 1341.060 1442.270 1341.200 1537.635 ;
        RECT 1341.000 1441.950 1341.260 1442.270 ;
        RECT 1340.540 1435.150 1340.800 1435.470 ;
        RECT 1340.600 1076.770 1340.740 1435.150 ;
        RECT 1340.540 1076.450 1340.800 1076.770 ;
        RECT 1341.000 1076.110 1341.260 1076.430 ;
        RECT 1341.060 983.010 1341.200 1076.110 ;
        RECT 1341.060 982.870 1341.660 983.010 ;
        RECT 1341.520 917.990 1341.660 982.870 ;
        RECT 1340.540 917.670 1340.800 917.990 ;
        RECT 1341.460 917.670 1341.720 917.990 ;
        RECT 1340.600 821.965 1340.740 917.670 ;
        RECT 1340.530 821.595 1340.810 821.965 ;
        RECT 1340.530 820.915 1340.810 821.285 ;
        RECT 1340.600 719.285 1340.740 820.915 ;
        RECT 1340.530 718.915 1340.810 719.285 ;
        RECT 1340.530 717.555 1340.810 717.925 ;
        RECT 1340.600 614.030 1340.740 717.555 ;
        RECT 1340.540 613.710 1340.800 614.030 ;
        RECT 1340.540 565.770 1340.800 566.090 ;
        RECT 1340.600 549.170 1340.740 565.770 ;
        RECT 1340.600 549.030 1341.200 549.170 ;
        RECT 1341.060 475.990 1341.200 549.030 ;
        RECT 1341.000 475.670 1341.260 475.990 ;
        RECT 1340.540 421.270 1340.800 421.590 ;
        RECT 1340.600 420.910 1340.740 421.270 ;
        RECT 1340.540 420.590 1340.800 420.910 ;
        RECT 1341.460 420.590 1341.720 420.910 ;
        RECT 1341.520 373.050 1341.660 420.590 ;
        RECT 1341.060 372.910 1341.660 373.050 ;
        RECT 1341.060 372.630 1341.200 372.910 ;
        RECT 1341.000 372.310 1341.260 372.630 ;
        RECT 1341.000 324.710 1341.260 325.030 ;
        RECT 1341.060 324.350 1341.200 324.710 ;
        RECT 1341.000 324.030 1341.260 324.350 ;
        RECT 1341.460 276.090 1341.720 276.410 ;
        RECT 1341.520 275.810 1341.660 276.090 ;
        RECT 1341.060 275.670 1341.660 275.810 ;
        RECT 1341.060 234.930 1341.200 275.670 ;
        RECT 1341.000 234.610 1341.260 234.930 ;
        RECT 1340.540 233.930 1340.800 234.250 ;
        RECT 1340.600 51.330 1340.740 233.930 ;
        RECT 724.140 51.010 724.400 51.330 ;
        RECT 1340.540 51.010 1340.800 51.330 ;
        RECT 724.200 3.130 724.340 51.010 ;
        RECT 722.360 2.990 724.340 3.130 ;
        RECT 722.360 2.400 722.500 2.990 ;
        RECT 722.150 -4.800 722.710 2.400 ;
      LAYER via2 ;
        RECT 1340.530 1579.840 1340.810 1580.120 ;
        RECT 1340.990 1537.680 1341.270 1537.960 ;
        RECT 1340.530 821.640 1340.810 821.920 ;
        RECT 1340.530 820.960 1340.810 821.240 ;
        RECT 1340.530 718.960 1340.810 719.240 ;
        RECT 1340.530 717.600 1340.810 717.880 ;
      LAYER met3 ;
        RECT 1340.505 1580.140 1340.835 1580.145 ;
        RECT 1340.505 1580.130 1341.090 1580.140 ;
        RECT 1340.505 1579.830 1341.290 1580.130 ;
        RECT 1340.505 1579.820 1341.090 1579.830 ;
        RECT 1340.505 1579.815 1340.835 1579.820 ;
        RECT 1340.965 1537.980 1341.295 1537.985 ;
        RECT 1340.710 1537.970 1341.295 1537.980 ;
        RECT 1340.510 1537.670 1341.295 1537.970 ;
        RECT 1340.710 1537.660 1341.295 1537.670 ;
        RECT 1340.965 1537.655 1341.295 1537.660 ;
        RECT 1340.505 821.930 1340.835 821.945 ;
        RECT 1340.505 821.615 1341.050 821.930 ;
        RECT 1340.750 821.265 1341.050 821.615 ;
        RECT 1340.505 820.950 1341.050 821.265 ;
        RECT 1340.505 820.935 1340.835 820.950 ;
        RECT 1340.505 719.250 1340.835 719.265 ;
        RECT 1340.505 718.935 1341.050 719.250 ;
        RECT 1340.750 717.905 1341.050 718.935 ;
        RECT 1340.505 717.590 1341.050 717.905 ;
        RECT 1340.505 717.575 1340.835 717.590 ;
      LAYER via3 ;
        RECT 1340.740 1579.820 1341.060 1580.140 ;
        RECT 1340.740 1537.660 1341.060 1537.980 ;
      LAYER met4 ;
        RECT 1340.735 1579.815 1341.065 1580.145 ;
        RECT 1340.750 1537.985 1341.050 1579.815 ;
        RECT 1340.735 1537.655 1341.065 1537.985 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1345.570 1694.120 1345.890 1694.180 ;
        RECT 1347.410 1694.120 1347.730 1694.180 ;
        RECT 1345.570 1693.980 1347.730 1694.120 ;
        RECT 1345.570 1693.920 1345.890 1693.980 ;
        RECT 1347.410 1693.920 1347.730 1693.980 ;
        RECT 724.110 1618.300 724.430 1618.360 ;
        RECT 1347.410 1618.300 1347.730 1618.360 ;
        RECT 724.110 1618.160 1347.730 1618.300 ;
        RECT 724.110 1618.100 724.430 1618.160 ;
        RECT 1347.410 1618.100 1347.730 1618.160 ;
      LAYER via ;
        RECT 1345.600 1693.920 1345.860 1694.180 ;
        RECT 1347.440 1693.920 1347.700 1694.180 ;
        RECT 724.140 1618.100 724.400 1618.360 ;
        RECT 1347.440 1618.100 1347.700 1618.360 ;
      LAYER met2 ;
        RECT 1345.590 1700.000 1345.870 1704.000 ;
        RECT 1345.660 1694.210 1345.800 1700.000 ;
        RECT 1345.600 1693.890 1345.860 1694.210 ;
        RECT 1347.440 1693.890 1347.700 1694.210 ;
        RECT 1347.500 1618.390 1347.640 1693.890 ;
        RECT 724.140 1618.070 724.400 1618.390 ;
        RECT 1347.440 1618.070 1347.700 1618.390 ;
        RECT 724.200 3.130 724.340 1618.070 ;
        RECT 722.360 2.990 724.340 3.130 ;
        RECT 722.360 2.400 722.500 2.990 ;
        RECT 722.150 -4.800 722.710 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 0.300 ;
=======
      LAYER met1 ;
        RECT 1609.610 1686.300 1609.930 1686.360 ;
        RECT 1613.750 1686.300 1614.070 1686.360 ;
        RECT 1609.610 1686.160 1614.070 1686.300 ;
        RECT 1609.610 1686.100 1609.930 1686.160 ;
        RECT 1613.750 1686.100 1614.070 1686.160 ;
        RECT 1613.750 18.940 1614.070 19.000 ;
        RECT 1703.450 18.940 1703.770 19.000 ;
        RECT 1613.750 18.800 1703.770 18.940 ;
        RECT 1613.750 18.740 1614.070 18.800 ;
        RECT 1703.450 18.740 1703.770 18.800 ;
      LAYER via ;
        RECT 1609.640 1686.100 1609.900 1686.360 ;
        RECT 1613.780 1686.100 1614.040 1686.360 ;
        RECT 1613.780 18.740 1614.040 19.000 ;
        RECT 1703.480 18.740 1703.740 19.000 ;
      LAYER met2 ;
        RECT 1609.630 1700.000 1609.910 1704.000 ;
        RECT 1609.700 1686.390 1609.840 1700.000 ;
        RECT 1609.640 1686.070 1609.900 1686.390 ;
        RECT 1613.780 1686.070 1614.040 1686.390 ;
        RECT 1613.840 19.030 1613.980 1686.070 ;
        RECT 1613.780 18.710 1614.040 19.030 ;
        RECT 1703.480 18.710 1703.740 19.030 ;
        RECT 1703.540 2.400 1703.680 18.710 ;
=======
      LAYER li1 ;
        RECT 1652.465 14.025 1652.635 15.215 ;
      LAYER mcon ;
        RECT 1652.465 15.045 1652.635 15.215 ;
      LAYER met1 ;
        RECT 1611.450 1689.700 1611.770 1689.760 ;
        RECT 1613.750 1689.700 1614.070 1689.760 ;
        RECT 1611.450 1689.560 1614.070 1689.700 ;
        RECT 1611.450 1689.500 1611.770 1689.560 ;
        RECT 1613.750 1689.500 1614.070 1689.560 ;
        RECT 1652.405 15.200 1652.695 15.245 ;
        RECT 1703.450 15.200 1703.770 15.260 ;
        RECT 1652.405 15.060 1703.770 15.200 ;
        RECT 1652.405 15.015 1652.695 15.060 ;
        RECT 1703.450 15.000 1703.770 15.060 ;
        RECT 1612.830 14.180 1613.150 14.240 ;
        RECT 1652.405 14.180 1652.695 14.225 ;
        RECT 1612.830 14.040 1652.695 14.180 ;
        RECT 1612.830 13.980 1613.150 14.040 ;
        RECT 1652.405 13.995 1652.695 14.040 ;
      LAYER via ;
        RECT 1611.480 1689.500 1611.740 1689.760 ;
        RECT 1613.780 1689.500 1614.040 1689.760 ;
        RECT 1703.480 15.000 1703.740 15.260 ;
        RECT 1612.860 13.980 1613.120 14.240 ;
      LAYER met2 ;
        RECT 1611.470 1700.000 1611.750 1704.000 ;
        RECT 1611.540 1689.790 1611.680 1700.000 ;
        RECT 1611.480 1689.470 1611.740 1689.790 ;
        RECT 1613.780 1689.470 1614.040 1689.790 ;
        RECT 1613.840 39.170 1613.980 1689.470 ;
        RECT 1612.920 39.030 1613.980 39.170 ;
        RECT 1612.920 14.270 1613.060 39.030 ;
        RECT 1703.480 14.970 1703.740 15.290 ;
        RECT 1612.860 13.950 1613.120 14.270 ;
        RECT 1703.540 2.400 1703.680 14.970 ;
>>>>>>> re-updated local openlane
        RECT 1703.330 -4.800 1703.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 0.300 ;
=======
      LAYER met1 ;
        RECT 1616.510 1684.940 1616.830 1685.000 ;
        RECT 1651.010 1684.940 1651.330 1685.000 ;
        RECT 1616.510 1684.800 1651.330 1684.940 ;
        RECT 1616.510 1684.740 1616.830 1684.800 ;
        RECT 1651.010 1684.740 1651.330 1684.800 ;
        RECT 1652.390 51.580 1652.710 51.640 ;
        RECT 1718.170 51.580 1718.490 51.640 ;
        RECT 1652.390 51.440 1718.490 51.580 ;
        RECT 1652.390 51.380 1652.710 51.440 ;
        RECT 1718.170 51.380 1718.490 51.440 ;
        RECT 1718.170 2.960 1718.490 3.020 ;
        RECT 1721.390 2.960 1721.710 3.020 ;
        RECT 1718.170 2.820 1721.710 2.960 ;
        RECT 1718.170 2.760 1718.490 2.820 ;
        RECT 1721.390 2.760 1721.710 2.820 ;
      LAYER via ;
        RECT 1616.540 1684.740 1616.800 1685.000 ;
        RECT 1651.040 1684.740 1651.300 1685.000 ;
        RECT 1652.420 51.380 1652.680 51.640 ;
        RECT 1718.200 51.380 1718.460 51.640 ;
        RECT 1718.200 2.760 1718.460 3.020 ;
        RECT 1721.420 2.760 1721.680 3.020 ;
      LAYER met2 ;
        RECT 1616.530 1700.000 1616.810 1704.000 ;
        RECT 1616.600 1685.030 1616.740 1700.000 ;
        RECT 1616.540 1684.710 1616.800 1685.030 ;
        RECT 1651.040 1684.710 1651.300 1685.030 ;
        RECT 1651.100 1676.610 1651.240 1684.710 ;
        RECT 1651.100 1676.470 1652.620 1676.610 ;
        RECT 1652.480 51.670 1652.620 1676.470 ;
        RECT 1652.420 51.350 1652.680 51.670 ;
        RECT 1718.200 51.350 1718.460 51.670 ;
        RECT 1718.260 3.050 1718.400 51.350 ;
        RECT 1718.200 2.730 1718.460 3.050 ;
        RECT 1721.420 2.730 1721.680 3.050 ;
        RECT 1721.480 2.400 1721.620 2.730 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1619.730 1683.920 1620.050 1683.980 ;
        RECT 1621.110 1683.920 1621.430 1683.980 ;
        RECT 1619.730 1683.780 1621.430 1683.920 ;
        RECT 1619.730 1683.720 1620.050 1683.780 ;
        RECT 1621.110 1683.720 1621.430 1683.780 ;
        RECT 1619.730 20.980 1620.050 21.040 ;
        RECT 1739.330 20.980 1739.650 21.040 ;
        RECT 1619.730 20.840 1739.650 20.980 ;
        RECT 1619.730 20.780 1620.050 20.840 ;
        RECT 1739.330 20.780 1739.650 20.840 ;
      LAYER via ;
        RECT 1619.760 1683.720 1620.020 1683.980 ;
        RECT 1621.140 1683.720 1621.400 1683.980 ;
        RECT 1619.760 20.780 1620.020 21.040 ;
        RECT 1739.360 20.780 1739.620 21.040 ;
      LAYER met2 ;
        RECT 1621.130 1700.000 1621.410 1704.000 ;
        RECT 1621.200 1684.010 1621.340 1700.000 ;
        RECT 1619.760 1683.690 1620.020 1684.010 ;
        RECT 1621.140 1683.690 1621.400 1684.010 ;
        RECT 1619.820 21.070 1619.960 1683.690 ;
        RECT 1619.760 20.750 1620.020 21.070 ;
        RECT 1739.360 20.750 1739.620 21.070 ;
        RECT 1739.420 2.400 1739.560 20.750 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1626.630 21.320 1626.950 21.380 ;
        RECT 1756.810 21.320 1757.130 21.380 ;
        RECT 1626.630 21.180 1757.130 21.320 ;
        RECT 1626.630 21.120 1626.950 21.180 ;
        RECT 1756.810 21.120 1757.130 21.180 ;
      LAYER via ;
        RECT 1626.660 21.120 1626.920 21.380 ;
        RECT 1756.840 21.120 1757.100 21.380 ;
      LAYER met2 ;
        RECT 1626.190 1700.410 1626.470 1704.000 ;
        RECT 1626.190 1700.270 1626.860 1700.410 ;
        RECT 1626.190 1700.000 1626.470 1700.270 ;
        RECT 1626.720 21.410 1626.860 1700.270 ;
        RECT 1626.660 21.090 1626.920 21.410 ;
        RECT 1756.840 21.090 1757.100 21.410 ;
        RECT 1756.900 2.400 1757.040 21.090 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1630.770 1685.620 1631.090 1685.680 ;
        RECT 1633.530 1685.620 1633.850 1685.680 ;
        RECT 1630.770 1685.480 1633.850 1685.620 ;
        RECT 1630.770 1685.420 1631.090 1685.480 ;
        RECT 1633.530 1685.420 1633.850 1685.480 ;
        RECT 1633.530 21.660 1633.850 21.720 ;
        RECT 1774.750 21.660 1775.070 21.720 ;
        RECT 1633.530 21.520 1775.070 21.660 ;
        RECT 1633.530 21.460 1633.850 21.520 ;
        RECT 1774.750 21.460 1775.070 21.520 ;
      LAYER via ;
        RECT 1630.800 1685.420 1631.060 1685.680 ;
        RECT 1633.560 1685.420 1633.820 1685.680 ;
        RECT 1633.560 21.460 1633.820 21.720 ;
        RECT 1774.780 21.460 1775.040 21.720 ;
      LAYER met2 ;
        RECT 1630.790 1700.000 1631.070 1704.000 ;
        RECT 1630.860 1685.710 1631.000 1700.000 ;
        RECT 1630.800 1685.390 1631.060 1685.710 ;
        RECT 1633.560 1685.390 1633.820 1685.710 ;
        RECT 1633.620 21.750 1633.760 1685.390 ;
        RECT 1633.560 21.430 1633.820 21.750 ;
        RECT 1774.780 21.430 1775.040 21.750 ;
        RECT 1774.840 2.400 1774.980 21.430 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 0.300 ;
=======
      LAYER met1 ;
        RECT 1635.830 1684.600 1636.150 1684.660 ;
        RECT 1641.350 1684.600 1641.670 1684.660 ;
        RECT 1635.830 1684.460 1641.670 1684.600 ;
        RECT 1635.830 1684.400 1636.150 1684.460 ;
        RECT 1641.350 1684.400 1641.670 1684.460 ;
        RECT 1641.350 22.000 1641.670 22.060 ;
        RECT 1792.690 22.000 1793.010 22.060 ;
        RECT 1641.350 21.860 1793.010 22.000 ;
        RECT 1641.350 21.800 1641.670 21.860 ;
        RECT 1792.690 21.800 1793.010 21.860 ;
      LAYER via ;
        RECT 1635.860 1684.400 1636.120 1684.660 ;
        RECT 1641.380 1684.400 1641.640 1684.660 ;
        RECT 1641.380 21.800 1641.640 22.060 ;
        RECT 1792.720 21.800 1792.980 22.060 ;
      LAYER met2 ;
        RECT 1635.850 1700.000 1636.130 1704.000 ;
        RECT 1635.920 1684.690 1636.060 1700.000 ;
        RECT 1635.860 1684.370 1636.120 1684.690 ;
        RECT 1641.380 1684.370 1641.640 1684.690 ;
        RECT 1641.440 22.090 1641.580 1684.370 ;
        RECT 1641.380 21.770 1641.640 22.090 ;
        RECT 1792.720 21.770 1792.980 22.090 ;
        RECT 1792.780 2.400 1792.920 21.770 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 0.300 ;
=======
      LAYER met1 ;
        RECT 1640.430 23.020 1640.750 23.080 ;
        RECT 1810.630 23.020 1810.950 23.080 ;
        RECT 1640.430 22.880 1810.950 23.020 ;
        RECT 1640.430 22.820 1640.750 22.880 ;
        RECT 1810.630 22.820 1810.950 22.880 ;
      LAYER via ;
        RECT 1640.460 22.820 1640.720 23.080 ;
        RECT 1810.660 22.820 1810.920 23.080 ;
      LAYER met2 ;
        RECT 1640.450 1700.000 1640.730 1704.000 ;
        RECT 1640.520 23.110 1640.660 1700.000 ;
        RECT 1640.460 22.790 1640.720 23.110 ;
        RECT 1810.660 22.790 1810.920 23.110 ;
        RECT 1810.720 2.400 1810.860 22.790 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1645.490 1683.920 1645.810 1683.980 ;
        RECT 1647.790 1683.920 1648.110 1683.980 ;
        RECT 1645.490 1683.780 1648.110 1683.920 ;
        RECT 1645.490 1683.720 1645.810 1683.780 ;
        RECT 1647.790 1683.720 1648.110 1683.780 ;
        RECT 1647.790 23.360 1648.110 23.420 ;
        RECT 1828.570 23.360 1828.890 23.420 ;
        RECT 1647.790 23.220 1828.890 23.360 ;
        RECT 1647.790 23.160 1648.110 23.220 ;
        RECT 1828.570 23.160 1828.890 23.220 ;
      LAYER via ;
        RECT 1645.520 1683.720 1645.780 1683.980 ;
        RECT 1647.820 1683.720 1648.080 1683.980 ;
        RECT 1647.820 23.160 1648.080 23.420 ;
        RECT 1828.600 23.160 1828.860 23.420 ;
      LAYER met2 ;
        RECT 1645.510 1700.000 1645.790 1704.000 ;
        RECT 1645.580 1684.010 1645.720 1700.000 ;
        RECT 1645.520 1683.690 1645.780 1684.010 ;
        RECT 1647.820 1683.690 1648.080 1684.010 ;
        RECT 1647.880 23.450 1648.020 1683.690 ;
        RECT 1647.820 23.130 1648.080 23.450 ;
        RECT 1828.600 23.130 1828.860 23.450 ;
        RECT 1828.660 2.400 1828.800 23.130 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1654.230 27.440 1654.550 27.500 ;
        RECT 1846.050 27.440 1846.370 27.500 ;
        RECT 1654.230 27.300 1846.370 27.440 ;
        RECT 1654.230 27.240 1654.550 27.300 ;
        RECT 1846.050 27.240 1846.370 27.300 ;
      LAYER via ;
        RECT 1654.260 27.240 1654.520 27.500 ;
        RECT 1846.080 27.240 1846.340 27.500 ;
      LAYER met2 ;
        RECT 1650.110 1700.410 1650.390 1704.000 ;
        RECT 1650.110 1700.270 1651.700 1700.410 ;
        RECT 1650.110 1700.000 1650.390 1700.270 ;
        RECT 1651.560 1677.290 1651.700 1700.270 ;
        RECT 1651.560 1677.150 1654.460 1677.290 ;
        RECT 1654.320 27.530 1654.460 1677.150 ;
        RECT 1654.260 27.210 1654.520 27.530 ;
        RECT 1846.080 27.210 1846.340 27.530 ;
        RECT 1846.140 2.400 1846.280 27.210 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 0.300 ;
=======
      LAYER li1 ;
        RECT 1802.425 22.865 1802.595 26.775 ;
      LAYER mcon ;
        RECT 1802.425 26.605 1802.595 26.775 ;
      LAYER met1 ;
        RECT 1654.690 26.760 1655.010 26.820 ;
        RECT 1802.365 26.760 1802.655 26.805 ;
        RECT 1654.690 26.620 1802.655 26.760 ;
        RECT 1654.690 26.560 1655.010 26.620 ;
        RECT 1802.365 26.575 1802.655 26.620 ;
        RECT 1802.365 23.020 1802.655 23.065 ;
        RECT 1863.990 23.020 1864.310 23.080 ;
        RECT 1802.365 22.880 1864.310 23.020 ;
        RECT 1802.365 22.835 1802.655 22.880 ;
        RECT 1863.990 22.820 1864.310 22.880 ;
      LAYER via ;
        RECT 1654.720 26.560 1654.980 26.820 ;
        RECT 1864.020 22.820 1864.280 23.080 ;
      LAYER met2 ;
        RECT 1652.870 1700.410 1653.150 1704.000 ;
        RECT 1652.870 1700.270 1654.460 1700.410 ;
        RECT 1652.870 1700.000 1653.150 1700.270 ;
        RECT 1654.320 1688.850 1654.460 1700.270 ;
        RECT 1654.320 1688.710 1654.920 1688.850 ;
        RECT 1654.780 26.850 1654.920 1688.710 ;
        RECT 1654.720 26.530 1654.980 26.850 ;
        RECT 1864.020 22.790 1864.280 23.110 ;
        RECT 1864.080 2.400 1864.220 22.790 ;
=======
      LAYER met1 ;
        RECT 1655.150 26.760 1655.470 26.820 ;
        RECT 1863.990 26.760 1864.310 26.820 ;
        RECT 1655.150 26.620 1864.310 26.760 ;
        RECT 1655.150 26.560 1655.470 26.620 ;
        RECT 1863.990 26.560 1864.310 26.620 ;
      LAYER via ;
        RECT 1655.180 26.560 1655.440 26.820 ;
        RECT 1864.020 26.560 1864.280 26.820 ;
      LAYER met2 ;
        RECT 1655.170 1700.000 1655.450 1704.000 ;
        RECT 1655.240 26.850 1655.380 1700.000 ;
        RECT 1655.180 26.530 1655.440 26.850 ;
        RECT 1864.020 26.530 1864.280 26.850 ;
        RECT 1864.080 2.400 1864.220 26.530 ;
>>>>>>> re-updated local openlane
        RECT 1863.870 -4.800 1864.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1346.030 1664.540 1346.350 1664.600 ;
        RECT 1349.250 1664.540 1349.570 1664.600 ;
        RECT 1346.030 1664.400 1349.570 1664.540 ;
        RECT 1346.030 1664.340 1346.350 1664.400 ;
        RECT 1349.250 1664.340 1349.570 1664.400 ;
        RECT 744.810 65.520 745.130 65.580 ;
        RECT 1346.030 65.520 1346.350 65.580 ;
        RECT 744.810 65.380 1346.350 65.520 ;
        RECT 744.810 65.320 745.130 65.380 ;
        RECT 1346.030 65.320 1346.350 65.380 ;
        RECT 740.210 2.960 740.530 3.020 ;
        RECT 744.810 2.960 745.130 3.020 ;
        RECT 740.210 2.820 745.130 2.960 ;
        RECT 740.210 2.760 740.530 2.820 ;
        RECT 744.810 2.760 745.130 2.820 ;
      LAYER via ;
        RECT 1346.060 1664.340 1346.320 1664.600 ;
        RECT 1349.280 1664.340 1349.540 1664.600 ;
        RECT 744.840 65.320 745.100 65.580 ;
        RECT 1346.060 65.320 1346.320 65.580 ;
        RECT 740.240 2.760 740.500 3.020 ;
        RECT 744.840 2.760 745.100 3.020 ;
      LAYER met2 ;
        RECT 1350.190 1700.410 1350.470 1704.000 ;
        RECT 1349.340 1700.270 1350.470 1700.410 ;
        RECT 1349.340 1664.630 1349.480 1700.270 ;
        RECT 1350.190 1700.000 1350.470 1700.270 ;
        RECT 1346.060 1664.310 1346.320 1664.630 ;
        RECT 1349.280 1664.310 1349.540 1664.630 ;
        RECT 1346.120 65.610 1346.260 1664.310 ;
        RECT 744.840 65.290 745.100 65.610 ;
        RECT 1346.060 65.290 1346.320 65.610 ;
        RECT 744.900 3.050 745.040 65.290 ;
        RECT 740.240 2.730 740.500 3.050 ;
        RECT 744.840 2.730 745.100 3.050 ;
        RECT 740.300 2.400 740.440 2.730 ;
        RECT 740.090 -4.800 740.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 0.300 ;
=======
      LAYER met1 ;
        RECT 1659.750 1683.920 1660.070 1683.980 ;
        RECT 1662.050 1683.920 1662.370 1683.980 ;
        RECT 1659.750 1683.780 1662.370 1683.920 ;
        RECT 1659.750 1683.720 1660.070 1683.780 ;
        RECT 1662.050 1683.720 1662.370 1683.780 ;
        RECT 1662.050 26.080 1662.370 26.140 ;
        RECT 1881.930 26.080 1882.250 26.140 ;
        RECT 1662.050 25.940 1882.250 26.080 ;
        RECT 1662.050 25.880 1662.370 25.940 ;
        RECT 1881.930 25.880 1882.250 25.940 ;
      LAYER via ;
        RECT 1659.780 1683.720 1660.040 1683.980 ;
        RECT 1662.080 1683.720 1662.340 1683.980 ;
        RECT 1662.080 25.880 1662.340 26.140 ;
        RECT 1881.960 25.880 1882.220 26.140 ;
      LAYER met2 ;
        RECT 1659.770 1700.000 1660.050 1704.000 ;
        RECT 1659.840 1684.010 1659.980 1700.000 ;
        RECT 1659.780 1683.690 1660.040 1684.010 ;
        RECT 1662.080 1683.690 1662.340 1684.010 ;
        RECT 1662.140 26.170 1662.280 1683.690 ;
        RECT 1662.080 25.850 1662.340 26.170 ;
        RECT 1881.960 25.850 1882.220 26.170 ;
        RECT 1882.020 2.400 1882.160 25.850 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1664.810 1684.260 1665.130 1684.320 ;
        RECT 1668.490 1684.260 1668.810 1684.320 ;
        RECT 1664.810 1684.120 1668.810 1684.260 ;
        RECT 1664.810 1684.060 1665.130 1684.120 ;
        RECT 1668.490 1684.060 1668.810 1684.120 ;
        RECT 1668.490 25.400 1668.810 25.460 ;
        RECT 1899.870 25.400 1900.190 25.460 ;
        RECT 1668.490 25.260 1900.190 25.400 ;
        RECT 1668.490 25.200 1668.810 25.260 ;
        RECT 1899.870 25.200 1900.190 25.260 ;
      LAYER via ;
        RECT 1664.840 1684.060 1665.100 1684.320 ;
        RECT 1668.520 1684.060 1668.780 1684.320 ;
        RECT 1668.520 25.200 1668.780 25.460 ;
        RECT 1899.900 25.200 1900.160 25.460 ;
      LAYER met2 ;
        RECT 1664.830 1700.000 1665.110 1704.000 ;
        RECT 1664.900 1684.350 1665.040 1700.000 ;
        RECT 1664.840 1684.030 1665.100 1684.350 ;
        RECT 1668.520 1684.030 1668.780 1684.350 ;
        RECT 1668.580 25.490 1668.720 1684.030 ;
        RECT 1668.520 25.170 1668.780 25.490 ;
        RECT 1899.900 25.170 1900.160 25.490 ;
        RECT 1899.960 2.400 1900.100 25.170 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1668.030 1683.920 1668.350 1683.980 ;
        RECT 1669.410 1683.920 1669.730 1683.980 ;
        RECT 1668.030 1683.780 1669.730 1683.920 ;
        RECT 1668.030 1683.720 1668.350 1683.780 ;
        RECT 1669.410 1683.720 1669.730 1683.780 ;
        RECT 1668.030 24.380 1668.350 24.440 ;
        RECT 1917.810 24.380 1918.130 24.440 ;
        RECT 1668.030 24.240 1918.130 24.380 ;
        RECT 1668.030 24.180 1668.350 24.240 ;
        RECT 1917.810 24.180 1918.130 24.240 ;
      LAYER via ;
        RECT 1668.060 1683.720 1668.320 1683.980 ;
        RECT 1669.440 1683.720 1669.700 1683.980 ;
        RECT 1668.060 24.180 1668.320 24.440 ;
        RECT 1917.840 24.180 1918.100 24.440 ;
      LAYER met2 ;
        RECT 1669.430 1700.000 1669.710 1704.000 ;
        RECT 1669.500 1684.010 1669.640 1700.000 ;
        RECT 1668.060 1683.690 1668.320 1684.010 ;
        RECT 1669.440 1683.690 1669.700 1684.010 ;
        RECT 1668.120 24.470 1668.260 1683.690 ;
        RECT 1668.060 24.150 1668.320 24.470 ;
        RECT 1917.840 24.150 1918.100 24.470 ;
        RECT 1917.900 2.400 1918.040 24.150 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 0.300 ;
=======
      LAYER li1 ;
        RECT 1919.265 24.055 1919.435 24.735 ;
        RECT 1918.345 23.885 1919.435 24.055 ;
      LAYER mcon ;
        RECT 1919.265 24.565 1919.435 24.735 ;
      LAYER met1 ;
        RECT 1672.170 1688.680 1672.490 1688.740 ;
        RECT 1675.390 1688.680 1675.710 1688.740 ;
        RECT 1672.170 1688.540 1675.710 1688.680 ;
        RECT 1672.170 1688.480 1672.490 1688.540 ;
        RECT 1675.390 1688.480 1675.710 1688.540 ;
        RECT 1919.205 24.720 1919.495 24.765 ;
        RECT 1935.290 24.720 1935.610 24.780 ;
        RECT 1919.205 24.580 1935.610 24.720 ;
        RECT 1919.205 24.535 1919.495 24.580 ;
        RECT 1935.290 24.520 1935.610 24.580 ;
        RECT 1675.390 24.040 1675.710 24.100 ;
        RECT 1918.285 24.040 1918.575 24.085 ;
        RECT 1675.390 23.900 1918.575 24.040 ;
        RECT 1675.390 23.840 1675.710 23.900 ;
        RECT 1918.285 23.855 1918.575 23.900 ;
      LAYER via ;
        RECT 1672.200 1688.480 1672.460 1688.740 ;
        RECT 1675.420 1688.480 1675.680 1688.740 ;
        RECT 1935.320 24.520 1935.580 24.780 ;
        RECT 1675.420 23.840 1675.680 24.100 ;
      LAYER met2 ;
        RECT 1672.190 1700.000 1672.470 1704.000 ;
        RECT 1672.260 1688.770 1672.400 1700.000 ;
        RECT 1672.200 1688.450 1672.460 1688.770 ;
        RECT 1675.420 1688.450 1675.680 1688.770 ;
        RECT 1675.480 24.130 1675.620 1688.450 ;
        RECT 1935.320 24.490 1935.580 24.810 ;
        RECT 1675.420 23.810 1675.680 24.130 ;
        RECT 1935.380 2.400 1935.520 24.490 ;
=======
      LAYER met1 ;
        RECT 1674.470 1683.920 1674.790 1683.980 ;
        RECT 1675.850 1683.920 1676.170 1683.980 ;
        RECT 1674.470 1683.780 1676.170 1683.920 ;
        RECT 1674.470 1683.720 1674.790 1683.780 ;
        RECT 1675.850 1683.720 1676.170 1683.780 ;
        RECT 1675.850 24.040 1676.170 24.100 ;
        RECT 1935.290 24.040 1935.610 24.100 ;
        RECT 1675.850 23.900 1935.610 24.040 ;
        RECT 1675.850 23.840 1676.170 23.900 ;
        RECT 1935.290 23.840 1935.610 23.900 ;
      LAYER via ;
        RECT 1674.500 1683.720 1674.760 1683.980 ;
        RECT 1675.880 1683.720 1676.140 1683.980 ;
        RECT 1675.880 23.840 1676.140 24.100 ;
        RECT 1935.320 23.840 1935.580 24.100 ;
      LAYER met2 ;
        RECT 1674.490 1700.000 1674.770 1704.000 ;
        RECT 1674.560 1684.010 1674.700 1700.000 ;
        RECT 1674.500 1683.690 1674.760 1684.010 ;
        RECT 1675.880 1683.690 1676.140 1684.010 ;
        RECT 1675.940 24.130 1676.080 1683.690 ;
        RECT 1675.880 23.810 1676.140 24.130 ;
        RECT 1935.320 23.810 1935.580 24.130 ;
        RECT 1935.380 2.400 1935.520 23.810 ;
>>>>>>> re-updated local openlane
        RECT 1935.170 -4.800 1935.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1679.070 1683.920 1679.390 1683.980 ;
        RECT 1682.750 1683.920 1683.070 1683.980 ;
        RECT 1679.070 1683.780 1683.070 1683.920 ;
        RECT 1679.070 1683.720 1679.390 1683.780 ;
        RECT 1682.750 1683.720 1683.070 1683.780 ;
      LAYER via ;
        RECT 1679.100 1683.720 1679.360 1683.980 ;
        RECT 1682.780 1683.720 1683.040 1683.980 ;
      LAYER met2 ;
        RECT 1679.090 1700.000 1679.370 1704.000 ;
        RECT 1679.160 1684.010 1679.300 1700.000 ;
        RECT 1679.100 1683.690 1679.360 1684.010 ;
        RECT 1682.780 1683.690 1683.040 1684.010 ;
        RECT 1682.840 24.325 1682.980 1683.690 ;
        RECT 1682.770 23.955 1683.050 24.325 ;
        RECT 1953.250 23.955 1953.530 24.325 ;
        RECT 1953.320 2.400 1953.460 23.955 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
      LAYER via2 ;
        RECT 1682.770 24.000 1683.050 24.280 ;
        RECT 1953.250 24.000 1953.530 24.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1682.745 27.690 1683.075 27.705 ;
        RECT 1953.225 27.690 1953.555 27.705 ;
        RECT 1682.745 27.390 1953.555 27.690 ;
        RECT 1682.745 27.375 1683.075 27.390 ;
        RECT 1953.225 27.375 1953.555 27.390 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1682.745 24.290 1683.075 24.305 ;
        RECT 1953.225 24.290 1953.555 24.305 ;
        RECT 1682.745 23.990 1953.555 24.290 ;
        RECT 1682.745 23.975 1683.075 23.990 ;
        RECT 1953.225 23.975 1953.555 23.990 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1684.130 1673.380 1684.450 1673.440 ;
        RECT 1966.570 1673.380 1966.890 1673.440 ;
        RECT 1684.130 1673.240 1966.890 1673.380 ;
        RECT 1684.130 1673.180 1684.450 1673.240 ;
        RECT 1966.570 1673.180 1966.890 1673.240 ;
        RECT 1966.570 62.120 1966.890 62.180 ;
        RECT 1971.170 62.120 1971.490 62.180 ;
        RECT 1966.570 61.980 1971.490 62.120 ;
        RECT 1966.570 61.920 1966.890 61.980 ;
        RECT 1971.170 61.920 1971.490 61.980 ;
      LAYER via ;
        RECT 1684.160 1673.180 1684.420 1673.440 ;
        RECT 1966.600 1673.180 1966.860 1673.440 ;
        RECT 1966.600 61.920 1966.860 62.180 ;
        RECT 1971.200 61.920 1971.460 62.180 ;
      LAYER met2 ;
        RECT 1684.150 1700.000 1684.430 1704.000 ;
        RECT 1684.220 1673.470 1684.360 1700.000 ;
        RECT 1684.160 1673.150 1684.420 1673.470 ;
        RECT 1966.600 1673.150 1966.860 1673.470 ;
        RECT 1966.660 62.210 1966.800 1673.150 ;
        RECT 1966.600 61.890 1966.860 62.210 ;
        RECT 1971.200 61.890 1971.460 62.210 ;
        RECT 1971.260 2.400 1971.400 61.890 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1688.270 42.060 1688.590 42.120 ;
        RECT 1989.110 42.060 1989.430 42.120 ;
        RECT 1688.270 41.920 1989.430 42.060 ;
        RECT 1688.270 41.860 1688.590 41.920 ;
        RECT 1989.110 41.860 1989.430 41.920 ;
      LAYER via ;
        RECT 1688.300 41.860 1688.560 42.120 ;
        RECT 1989.140 41.860 1989.400 42.120 ;
      LAYER met2 ;
        RECT 1686.910 1700.410 1687.190 1704.000 ;
        RECT 1686.910 1700.270 1687.580 1700.410 ;
        RECT 1686.910 1700.000 1687.190 1700.270 ;
        RECT 1687.440 1688.680 1687.580 1700.270 ;
        RECT 1687.440 1688.540 1688.500 1688.680 ;
        RECT 1688.360 42.150 1688.500 1688.540 ;
        RECT 1688.300 41.830 1688.560 42.150 ;
        RECT 1989.140 41.830 1989.400 42.150 ;
        RECT 1989.200 2.400 1989.340 41.830 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1987.345 1587.205 1987.515 1618.315 ;
        RECT 1987.345 959.225 1987.515 1006.995 ;
        RECT 1987.345 766.105 1987.515 814.215 ;
        RECT 1987.345 669.545 1987.515 717.655 ;
        RECT 1987.345 572.645 1987.515 620.755 ;
        RECT 1987.345 476.085 1987.515 524.195 ;
        RECT 1987.345 379.525 1987.515 427.635 ;
        RECT 1987.345 282.965 1987.515 331.075 ;
        RECT 1986.425 186.405 1986.595 234.515 ;
        RECT 1987.345 61.285 1987.515 137.955 ;
      LAYER mcon ;
        RECT 1987.345 1618.145 1987.515 1618.315 ;
        RECT 1987.345 1006.825 1987.515 1006.995 ;
        RECT 1987.345 814.045 1987.515 814.215 ;
        RECT 1987.345 717.485 1987.515 717.655 ;
        RECT 1987.345 620.585 1987.515 620.755 ;
        RECT 1987.345 524.025 1987.515 524.195 ;
        RECT 1987.345 427.465 1987.515 427.635 ;
        RECT 1987.345 330.905 1987.515 331.075 ;
        RECT 1986.425 234.345 1986.595 234.515 ;
        RECT 1987.345 137.785 1987.515 137.955 ;
      LAYER met1 ;
        RECT 1689.650 1618.300 1689.970 1618.360 ;
        RECT 1987.285 1618.300 1987.575 1618.345 ;
        RECT 1689.650 1618.160 1987.575 1618.300 ;
        RECT 1689.650 1618.100 1689.970 1618.160 ;
        RECT 1987.285 1618.115 1987.575 1618.160 ;
        RECT 1987.270 1587.360 1987.590 1587.420 ;
        RECT 1987.075 1587.220 1987.590 1587.360 ;
        RECT 1987.270 1587.160 1987.590 1587.220 ;
        RECT 1986.810 1539.080 1987.130 1539.140 ;
        RECT 1987.270 1539.080 1987.590 1539.140 ;
        RECT 1986.810 1538.940 1987.590 1539.080 ;
        RECT 1986.810 1538.880 1987.130 1538.940 ;
        RECT 1987.270 1538.880 1987.590 1538.940 ;
        RECT 1987.270 1442.180 1987.590 1442.240 ;
        RECT 1987.730 1442.180 1988.050 1442.240 ;
        RECT 1987.270 1442.040 1988.050 1442.180 ;
        RECT 1987.270 1441.980 1987.590 1442.040 ;
        RECT 1987.730 1441.980 1988.050 1442.040 ;
        RECT 1987.270 1006.980 1987.590 1007.040 ;
        RECT 1987.075 1006.840 1987.590 1006.980 ;
        RECT 1987.270 1006.780 1987.590 1006.840 ;
        RECT 1987.270 959.380 1987.590 959.440 ;
        RECT 1987.075 959.240 1987.590 959.380 ;
        RECT 1987.270 959.180 1987.590 959.240 ;
        RECT 1986.810 821.340 1987.130 821.400 ;
        RECT 1987.270 821.340 1987.590 821.400 ;
        RECT 1986.810 821.200 1987.590 821.340 ;
        RECT 1986.810 821.140 1987.130 821.200 ;
        RECT 1987.270 821.140 1987.590 821.200 ;
        RECT 1987.270 814.200 1987.590 814.260 ;
        RECT 1987.075 814.060 1987.590 814.200 ;
        RECT 1987.270 814.000 1987.590 814.060 ;
        RECT 1987.270 766.260 1987.590 766.320 ;
        RECT 1987.075 766.120 1987.590 766.260 ;
        RECT 1987.270 766.060 1987.590 766.120 ;
        RECT 1987.270 717.640 1987.590 717.700 ;
        RECT 1987.075 717.500 1987.590 717.640 ;
        RECT 1987.270 717.440 1987.590 717.500 ;
        RECT 1987.270 669.700 1987.590 669.760 ;
        RECT 1987.075 669.560 1987.590 669.700 ;
        RECT 1987.270 669.500 1987.590 669.560 ;
        RECT 1987.270 620.740 1987.590 620.800 ;
        RECT 1987.075 620.600 1987.590 620.740 ;
        RECT 1987.270 620.540 1987.590 620.600 ;
        RECT 1987.270 572.800 1987.590 572.860 ;
        RECT 1987.075 572.660 1987.590 572.800 ;
        RECT 1987.270 572.600 1987.590 572.660 ;
        RECT 1987.270 524.180 1987.590 524.240 ;
        RECT 1987.075 524.040 1987.590 524.180 ;
        RECT 1987.270 523.980 1987.590 524.040 ;
        RECT 1987.270 476.240 1987.590 476.300 ;
        RECT 1987.075 476.100 1987.590 476.240 ;
        RECT 1987.270 476.040 1987.590 476.100 ;
        RECT 1987.270 427.620 1987.590 427.680 ;
        RECT 1987.075 427.480 1987.590 427.620 ;
        RECT 1987.270 427.420 1987.590 427.480 ;
        RECT 1987.270 379.680 1987.590 379.740 ;
        RECT 1987.075 379.540 1987.590 379.680 ;
        RECT 1987.270 379.480 1987.590 379.540 ;
        RECT 1987.270 331.060 1987.590 331.120 ;
        RECT 1987.075 330.920 1987.590 331.060 ;
        RECT 1987.270 330.860 1987.590 330.920 ;
        RECT 1987.270 283.120 1987.590 283.180 ;
        RECT 1987.075 282.980 1987.590 283.120 ;
        RECT 1987.270 282.920 1987.590 282.980 ;
        RECT 1986.365 234.500 1986.655 234.545 ;
        RECT 1987.270 234.500 1987.590 234.560 ;
        RECT 1986.365 234.360 1987.590 234.500 ;
        RECT 1986.365 234.315 1986.655 234.360 ;
        RECT 1987.270 234.300 1987.590 234.360 ;
        RECT 1986.350 186.560 1986.670 186.620 ;
        RECT 1986.155 186.420 1986.670 186.560 ;
        RECT 1986.350 186.360 1986.670 186.420 ;
        RECT 1987.270 137.940 1987.590 138.000 ;
        RECT 1987.075 137.800 1987.590 137.940 ;
        RECT 1987.270 137.740 1987.590 137.800 ;
        RECT 1987.285 61.440 1987.575 61.485 ;
        RECT 1989.110 61.440 1989.430 61.500 ;
        RECT 1987.285 61.300 1989.430 61.440 ;
        RECT 1987.285 61.255 1987.575 61.300 ;
        RECT 1989.110 61.240 1989.430 61.300 ;
      LAYER via ;
        RECT 1689.680 1618.100 1689.940 1618.360 ;
        RECT 1987.300 1587.160 1987.560 1587.420 ;
        RECT 1986.840 1538.880 1987.100 1539.140 ;
        RECT 1987.300 1538.880 1987.560 1539.140 ;
        RECT 1987.300 1441.980 1987.560 1442.240 ;
        RECT 1987.760 1441.980 1988.020 1442.240 ;
        RECT 1987.300 1006.780 1987.560 1007.040 ;
        RECT 1987.300 959.180 1987.560 959.440 ;
        RECT 1986.840 821.140 1987.100 821.400 ;
        RECT 1987.300 821.140 1987.560 821.400 ;
        RECT 1987.300 814.000 1987.560 814.260 ;
        RECT 1987.300 766.060 1987.560 766.320 ;
        RECT 1987.300 717.440 1987.560 717.700 ;
        RECT 1987.300 669.500 1987.560 669.760 ;
        RECT 1987.300 620.540 1987.560 620.800 ;
        RECT 1987.300 572.600 1987.560 572.860 ;
        RECT 1987.300 523.980 1987.560 524.240 ;
        RECT 1987.300 476.040 1987.560 476.300 ;
        RECT 1987.300 427.420 1987.560 427.680 ;
        RECT 1987.300 379.480 1987.560 379.740 ;
        RECT 1987.300 330.860 1987.560 331.120 ;
        RECT 1987.300 282.920 1987.560 283.180 ;
        RECT 1987.300 234.300 1987.560 234.560 ;
        RECT 1986.380 186.360 1986.640 186.620 ;
        RECT 1987.300 137.740 1987.560 138.000 ;
        RECT 1989.140 61.240 1989.400 61.500 ;
      LAYER met2 ;
        RECT 1689.210 1700.410 1689.490 1704.000 ;
        RECT 1689.210 1700.270 1689.880 1700.410 ;
        RECT 1689.210 1700.000 1689.490 1700.270 ;
        RECT 1689.740 1618.390 1689.880 1700.270 ;
        RECT 1689.680 1618.070 1689.940 1618.390 ;
        RECT 1987.300 1587.130 1987.560 1587.450 ;
        RECT 1987.360 1586.850 1987.500 1587.130 ;
        RECT 1986.900 1586.710 1987.500 1586.850 ;
        RECT 1986.900 1539.170 1987.040 1586.710 ;
        RECT 1986.840 1538.850 1987.100 1539.170 ;
        RECT 1987.300 1538.850 1987.560 1539.170 ;
        RECT 1987.360 1490.290 1987.500 1538.850 ;
        RECT 1987.360 1490.150 1987.960 1490.290 ;
        RECT 1987.820 1442.270 1987.960 1490.150 ;
        RECT 1987.300 1441.950 1987.560 1442.270 ;
        RECT 1987.760 1441.950 1988.020 1442.270 ;
        RECT 1987.360 1007.070 1987.500 1441.950 ;
        RECT 1987.300 1006.750 1987.560 1007.070 ;
        RECT 1987.300 959.150 1987.560 959.470 ;
        RECT 1987.360 869.450 1987.500 959.150 ;
        RECT 1986.900 869.310 1987.500 869.450 ;
        RECT 1986.900 821.430 1987.040 869.310 ;
        RECT 1986.840 821.110 1987.100 821.430 ;
        RECT 1987.300 821.110 1987.560 821.430 ;
        RECT 1987.360 814.290 1987.500 821.110 ;
        RECT 1987.300 813.970 1987.560 814.290 ;
        RECT 1987.300 766.030 1987.560 766.350 ;
        RECT 1987.360 717.730 1987.500 766.030 ;
        RECT 1987.300 717.410 1987.560 717.730 ;
        RECT 1987.300 669.470 1987.560 669.790 ;
        RECT 1987.360 620.830 1987.500 669.470 ;
        RECT 1987.300 620.510 1987.560 620.830 ;
        RECT 1987.300 572.570 1987.560 572.890 ;
        RECT 1987.360 524.270 1987.500 572.570 ;
        RECT 1987.300 523.950 1987.560 524.270 ;
        RECT 1987.300 476.010 1987.560 476.330 ;
        RECT 1987.360 427.710 1987.500 476.010 ;
        RECT 1987.300 427.390 1987.560 427.710 ;
        RECT 1987.300 379.450 1987.560 379.770 ;
        RECT 1987.360 331.150 1987.500 379.450 ;
        RECT 1987.300 330.830 1987.560 331.150 ;
        RECT 1987.300 282.890 1987.560 283.210 ;
        RECT 1987.360 234.590 1987.500 282.890 ;
        RECT 1987.300 234.270 1987.560 234.590 ;
        RECT 1986.380 186.330 1986.640 186.650 ;
        RECT 1986.440 145.365 1986.580 186.330 ;
        RECT 1986.370 144.995 1986.650 145.365 ;
        RECT 1987.290 144.995 1987.570 145.365 ;
        RECT 1987.360 138.030 1987.500 144.995 ;
        RECT 1987.300 137.710 1987.560 138.030 ;
        RECT 1989.140 61.210 1989.400 61.530 ;
        RECT 1989.200 2.400 1989.340 61.210 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
      LAYER via2 ;
        RECT 1986.370 145.040 1986.650 145.320 ;
        RECT 1987.290 145.040 1987.570 145.320 ;
      LAYER met3 ;
        RECT 1986.345 145.330 1986.675 145.345 ;
        RECT 1987.265 145.330 1987.595 145.345 ;
        RECT 1986.345 145.030 1987.595 145.330 ;
        RECT 1986.345 145.015 1986.675 145.030 ;
        RECT 1987.265 145.015 1987.595 145.030 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1695.630 58.720 1695.950 58.780 ;
        RECT 2006.590 58.720 2006.910 58.780 ;
        RECT 1695.630 58.580 2006.910 58.720 ;
        RECT 1695.630 58.520 1695.950 58.580 ;
        RECT 2006.590 58.520 2006.910 58.580 ;
      LAYER via ;
        RECT 1695.660 58.520 1695.920 58.780 ;
        RECT 2006.620 58.520 2006.880 58.780 ;
      LAYER met2 ;
        RECT 1693.810 1700.410 1694.090 1704.000 ;
        RECT 1693.810 1700.270 1694.940 1700.410 ;
        RECT 1693.810 1700.000 1694.090 1700.270 ;
        RECT 1694.800 1656.210 1694.940 1700.270 ;
        RECT 1694.800 1656.070 1695.860 1656.210 ;
        RECT 1695.720 58.810 1695.860 1656.070 ;
        RECT 1695.660 58.490 1695.920 58.810 ;
        RECT 2006.620 58.490 2006.880 58.810 ;
        RECT 2006.680 2.400 2006.820 58.490 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 0.300 ;
=======
      LAYER met1 ;
        RECT 1698.850 1683.920 1699.170 1683.980 ;
        RECT 1702.990 1683.920 1703.310 1683.980 ;
        RECT 1698.850 1683.780 1703.310 1683.920 ;
        RECT 1698.850 1683.720 1699.170 1683.780 ;
        RECT 1702.990 1683.720 1703.310 1683.780 ;
        RECT 1702.990 1625.100 1703.310 1625.160 ;
        RECT 2021.770 1625.100 2022.090 1625.160 ;
        RECT 1702.990 1624.960 2022.090 1625.100 ;
        RECT 1702.990 1624.900 1703.310 1624.960 ;
        RECT 2021.770 1624.900 2022.090 1624.960 ;
        RECT 2021.770 62.120 2022.090 62.180 ;
        RECT 2024.530 62.120 2024.850 62.180 ;
        RECT 2021.770 61.980 2024.850 62.120 ;
        RECT 2021.770 61.920 2022.090 61.980 ;
        RECT 2024.530 61.920 2024.850 61.980 ;
      LAYER via ;
        RECT 1698.880 1683.720 1699.140 1683.980 ;
        RECT 1703.020 1683.720 1703.280 1683.980 ;
        RECT 1703.020 1624.900 1703.280 1625.160 ;
        RECT 2021.800 1624.900 2022.060 1625.160 ;
        RECT 2021.800 61.920 2022.060 62.180 ;
        RECT 2024.560 61.920 2024.820 62.180 ;
      LAYER met2 ;
        RECT 1698.870 1700.000 1699.150 1704.000 ;
        RECT 1698.940 1684.010 1699.080 1700.000 ;
        RECT 1698.880 1683.690 1699.140 1684.010 ;
        RECT 1703.020 1683.690 1703.280 1684.010 ;
        RECT 1703.080 1625.190 1703.220 1683.690 ;
        RECT 1703.020 1624.870 1703.280 1625.190 ;
        RECT 2021.800 1624.870 2022.060 1625.190 ;
        RECT 2021.860 62.210 2022.000 1624.870 ;
        RECT 2021.800 61.890 2022.060 62.210 ;
        RECT 2024.560 61.890 2024.820 62.210 ;
        RECT 2024.620 2.400 2024.760 61.890 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1703.910 1666.920 1704.230 1666.980 ;
        RECT 2042.470 1666.920 2042.790 1666.980 ;
        RECT 1703.910 1666.780 2042.790 1666.920 ;
        RECT 1703.910 1666.720 1704.230 1666.780 ;
        RECT 2042.470 1666.720 2042.790 1666.780 ;
      LAYER via ;
        RECT 1703.940 1666.720 1704.200 1666.980 ;
        RECT 2042.500 1666.720 2042.760 1666.980 ;
      LAYER met2 ;
        RECT 1703.470 1700.410 1703.750 1704.000 ;
        RECT 1703.470 1700.270 1704.140 1700.410 ;
        RECT 1703.470 1700.000 1703.750 1700.270 ;
        RECT 1704.000 1667.010 1704.140 1700.270 ;
        RECT 1703.940 1666.690 1704.200 1667.010 ;
        RECT 2042.500 1666.690 2042.760 1667.010 ;
        RECT 2042.560 2.400 2042.700 1666.690 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 0.300 ;
=======
      LAYER met1 ;
        RECT 758.610 1673.040 758.930 1673.100 ;
        RECT 1355.230 1673.040 1355.550 1673.100 ;
        RECT 758.610 1672.900 1355.550 1673.040 ;
        RECT 758.610 1672.840 758.930 1672.900 ;
        RECT 1355.230 1672.840 1355.550 1672.900 ;
        RECT 757.690 2.960 758.010 3.020 ;
        RECT 758.610 2.960 758.930 3.020 ;
        RECT 757.690 2.820 758.930 2.960 ;
        RECT 757.690 2.760 758.010 2.820 ;
        RECT 758.610 2.760 758.930 2.820 ;
      LAYER via ;
        RECT 758.640 1672.840 758.900 1673.100 ;
        RECT 1355.260 1672.840 1355.520 1673.100 ;
        RECT 757.720 2.760 757.980 3.020 ;
        RECT 758.640 2.760 758.900 3.020 ;
      LAYER met2 ;
        RECT 1355.250 1700.000 1355.530 1704.000 ;
        RECT 1355.320 1673.130 1355.460 1700.000 ;
        RECT 758.640 1672.810 758.900 1673.130 ;
        RECT 1355.260 1672.810 1355.520 1673.130 ;
        RECT 758.700 3.050 758.840 1672.810 ;
        RECT 757.720 2.730 757.980 3.050 ;
        RECT 758.640 2.730 758.900 3.050 ;
        RECT 757.780 2.400 757.920 2.730 ;
        RECT 757.570 -4.800 758.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1708.510 1684.260 1708.830 1684.320 ;
        RECT 1709.890 1684.260 1710.210 1684.320 ;
        RECT 1708.510 1684.120 1710.210 1684.260 ;
        RECT 1708.510 1684.060 1708.830 1684.120 ;
        RECT 1709.890 1684.060 1710.210 1684.120 ;
        RECT 1709.890 1604.700 1710.210 1604.760 ;
        RECT 2056.270 1604.700 2056.590 1604.760 ;
        RECT 1709.890 1604.560 2056.590 1604.700 ;
        RECT 1709.890 1604.500 1710.210 1604.560 ;
        RECT 2056.270 1604.500 2056.590 1604.560 ;
        RECT 2056.270 62.120 2056.590 62.180 ;
        RECT 2060.410 62.120 2060.730 62.180 ;
        RECT 2056.270 61.980 2060.730 62.120 ;
        RECT 2056.270 61.920 2056.590 61.980 ;
        RECT 2060.410 61.920 2060.730 61.980 ;
      LAYER via ;
        RECT 1708.540 1684.060 1708.800 1684.320 ;
        RECT 1709.920 1684.060 1710.180 1684.320 ;
        RECT 1709.920 1604.500 1710.180 1604.760 ;
        RECT 2056.300 1604.500 2056.560 1604.760 ;
        RECT 2056.300 61.920 2056.560 62.180 ;
        RECT 2060.440 61.920 2060.700 62.180 ;
      LAYER met2 ;
        RECT 1708.530 1700.000 1708.810 1704.000 ;
        RECT 1708.600 1684.350 1708.740 1700.000 ;
        RECT 1708.540 1684.030 1708.800 1684.350 ;
        RECT 1709.920 1684.030 1710.180 1684.350 ;
        RECT 1709.980 1604.790 1710.120 1684.030 ;
        RECT 1709.920 1604.470 1710.180 1604.790 ;
        RECT 2056.300 1604.470 2056.560 1604.790 ;
        RECT 2056.360 62.210 2056.500 1604.470 ;
        RECT 2056.300 61.890 2056.560 62.210 ;
        RECT 2060.440 61.890 2060.700 62.210 ;
        RECT 2060.500 2.400 2060.640 61.890 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 0.300 ;
=======
      LAYER met1 ;
        RECT 1709.430 28.460 1709.750 28.520 ;
        RECT 2078.350 28.460 2078.670 28.520 ;
        RECT 1709.430 28.320 2078.670 28.460 ;
        RECT 1709.430 28.260 1709.750 28.320 ;
        RECT 2078.350 28.260 2078.670 28.320 ;
      LAYER via ;
        RECT 1709.460 28.260 1709.720 28.520 ;
        RECT 2078.380 28.260 2078.640 28.520 ;
      LAYER met2 ;
        RECT 1710.830 1700.410 1711.110 1704.000 ;
        RECT 1709.980 1700.270 1711.110 1700.410 ;
        RECT 1709.980 1688.680 1710.120 1700.270 ;
        RECT 1710.830 1700.000 1711.110 1700.270 ;
        RECT 1709.520 1688.540 1710.120 1688.680 ;
        RECT 1709.520 28.550 1709.660 1688.540 ;
        RECT 1709.460 28.230 1709.720 28.550 ;
        RECT 2078.380 28.230 2078.640 28.550 ;
        RECT 2078.440 2.400 2078.580 28.230 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 2077.045 1594.005 2077.215 1642.115 ;
        RECT 2077.045 1497.445 2077.215 1545.555 ;
        RECT 2077.045 1400.885 2077.215 1448.995 ;
        RECT 2077.045 1304.325 2077.215 1352.435 ;
        RECT 2077.045 1207.425 2077.215 1255.875 ;
        RECT 2077.045 628.065 2077.215 675.835 ;
        RECT 2077.045 531.505 2077.215 579.615 ;
        RECT 2077.045 434.945 2077.215 483.055 ;
        RECT 2077.045 338.045 2077.215 386.155 ;
        RECT 2077.045 48.365 2077.215 96.475 ;
      LAYER mcon ;
        RECT 2077.045 1641.945 2077.215 1642.115 ;
        RECT 2077.045 1545.385 2077.215 1545.555 ;
        RECT 2077.045 1448.825 2077.215 1448.995 ;
        RECT 2077.045 1352.265 2077.215 1352.435 ;
        RECT 2077.045 1255.705 2077.215 1255.875 ;
        RECT 2077.045 675.665 2077.215 675.835 ;
        RECT 2077.045 579.445 2077.215 579.615 ;
        RECT 2077.045 482.885 2077.215 483.055 ;
        RECT 2077.045 385.985 2077.215 386.155 ;
        RECT 2077.045 96.305 2077.215 96.475 ;
      LAYER met1 ;
        RECT 1713.110 1680.860 1713.430 1680.920 ;
        RECT 2076.970 1680.860 2077.290 1680.920 ;
        RECT 1713.110 1680.720 2077.290 1680.860 ;
        RECT 1713.110 1680.660 1713.430 1680.720 ;
        RECT 2076.970 1680.660 2077.290 1680.720 ;
        RECT 2076.970 1642.100 2077.290 1642.160 ;
        RECT 2076.970 1641.960 2077.485 1642.100 ;
        RECT 2076.970 1641.900 2077.290 1641.960 ;
        RECT 2076.970 1594.160 2077.290 1594.220 ;
        RECT 2076.970 1594.020 2077.485 1594.160 ;
        RECT 2076.970 1593.960 2077.290 1594.020 ;
        RECT 2076.970 1545.540 2077.290 1545.600 ;
        RECT 2076.970 1545.400 2077.485 1545.540 ;
        RECT 2076.970 1545.340 2077.290 1545.400 ;
        RECT 2076.970 1497.600 2077.290 1497.660 ;
        RECT 2076.970 1497.460 2077.485 1497.600 ;
        RECT 2076.970 1497.400 2077.290 1497.460 ;
        RECT 2076.970 1448.980 2077.290 1449.040 ;
        RECT 2076.970 1448.840 2077.485 1448.980 ;
        RECT 2076.970 1448.780 2077.290 1448.840 ;
        RECT 2076.970 1401.040 2077.290 1401.100 ;
        RECT 2076.970 1400.900 2077.485 1401.040 ;
        RECT 2076.970 1400.840 2077.290 1400.900 ;
        RECT 2076.970 1352.420 2077.290 1352.480 ;
        RECT 2076.970 1352.280 2077.485 1352.420 ;
        RECT 2076.970 1352.220 2077.290 1352.280 ;
        RECT 2076.970 1304.480 2077.290 1304.540 ;
        RECT 2076.970 1304.340 2077.485 1304.480 ;
        RECT 2076.970 1304.280 2077.290 1304.340 ;
        RECT 2076.970 1255.860 2077.290 1255.920 ;
        RECT 2076.970 1255.720 2077.485 1255.860 ;
        RECT 2076.970 1255.660 2077.290 1255.720 ;
        RECT 2076.970 1207.580 2077.290 1207.640 ;
        RECT 2076.970 1207.440 2077.485 1207.580 ;
        RECT 2076.970 1207.380 2077.290 1207.440 ;
        RECT 2076.970 1111.020 2077.290 1111.080 ;
        RECT 2077.890 1111.020 2078.210 1111.080 ;
        RECT 2076.970 1110.880 2078.210 1111.020 ;
        RECT 2076.970 1110.820 2077.290 1110.880 ;
        RECT 2077.890 1110.820 2078.210 1110.880 ;
        RECT 2076.970 1014.460 2077.290 1014.520 ;
        RECT 2077.890 1014.460 2078.210 1014.520 ;
        RECT 2076.970 1014.320 2078.210 1014.460 ;
        RECT 2076.970 1014.260 2077.290 1014.320 ;
        RECT 2077.890 1014.260 2078.210 1014.320 ;
        RECT 2076.970 917.900 2077.290 917.960 ;
        RECT 2077.890 917.900 2078.210 917.960 ;
        RECT 2076.970 917.760 2078.210 917.900 ;
        RECT 2076.970 917.700 2077.290 917.760 ;
        RECT 2077.890 917.700 2078.210 917.760 ;
        RECT 2076.970 772.720 2077.290 772.780 ;
        RECT 2077.890 772.720 2078.210 772.780 ;
        RECT 2076.970 772.580 2078.210 772.720 ;
        RECT 2076.970 772.520 2077.290 772.580 ;
        RECT 2077.890 772.520 2078.210 772.580 ;
        RECT 2076.970 675.820 2077.290 675.880 ;
        RECT 2076.970 675.680 2077.485 675.820 ;
        RECT 2076.970 675.620 2077.290 675.680 ;
        RECT 2076.970 628.220 2077.290 628.280 ;
        RECT 2076.970 628.080 2077.485 628.220 ;
        RECT 2076.970 628.020 2077.290 628.080 ;
        RECT 2076.970 579.600 2077.290 579.660 ;
        RECT 2076.970 579.460 2077.485 579.600 ;
        RECT 2076.970 579.400 2077.290 579.460 ;
        RECT 2076.970 531.660 2077.290 531.720 ;
        RECT 2076.970 531.520 2077.485 531.660 ;
        RECT 2076.970 531.460 2077.290 531.520 ;
        RECT 2076.970 483.040 2077.290 483.100 ;
        RECT 2076.970 482.900 2077.485 483.040 ;
        RECT 2076.970 482.840 2077.290 482.900 ;
        RECT 2076.970 435.100 2077.290 435.160 ;
        RECT 2076.970 434.960 2077.485 435.100 ;
        RECT 2076.970 434.900 2077.290 434.960 ;
        RECT 2076.970 386.140 2077.290 386.200 ;
        RECT 2076.970 386.000 2077.485 386.140 ;
        RECT 2076.970 385.940 2077.290 386.000 ;
        RECT 2076.970 338.200 2077.290 338.260 ;
        RECT 2076.970 338.060 2077.485 338.200 ;
        RECT 2076.970 338.000 2077.290 338.060 ;
        RECT 2076.970 96.460 2077.290 96.520 ;
        RECT 2076.970 96.320 2077.485 96.460 ;
        RECT 2076.970 96.260 2077.290 96.320 ;
        RECT 2076.985 48.520 2077.275 48.565 ;
        RECT 2078.350 48.520 2078.670 48.580 ;
        RECT 2076.985 48.380 2078.670 48.520 ;
        RECT 2076.985 48.335 2077.275 48.380 ;
        RECT 2078.350 48.320 2078.670 48.380 ;
      LAYER via ;
        RECT 1713.140 1680.660 1713.400 1680.920 ;
        RECT 2077.000 1680.660 2077.260 1680.920 ;
        RECT 2077.000 1641.900 2077.260 1642.160 ;
        RECT 2077.000 1593.960 2077.260 1594.220 ;
        RECT 2077.000 1545.340 2077.260 1545.600 ;
        RECT 2077.000 1497.400 2077.260 1497.660 ;
        RECT 2077.000 1448.780 2077.260 1449.040 ;
        RECT 2077.000 1400.840 2077.260 1401.100 ;
        RECT 2077.000 1352.220 2077.260 1352.480 ;
        RECT 2077.000 1304.280 2077.260 1304.540 ;
        RECT 2077.000 1255.660 2077.260 1255.920 ;
        RECT 2077.000 1207.380 2077.260 1207.640 ;
        RECT 2077.000 1110.820 2077.260 1111.080 ;
        RECT 2077.920 1110.820 2078.180 1111.080 ;
        RECT 2077.000 1014.260 2077.260 1014.520 ;
        RECT 2077.920 1014.260 2078.180 1014.520 ;
        RECT 2077.000 917.700 2077.260 917.960 ;
        RECT 2077.920 917.700 2078.180 917.960 ;
        RECT 2077.000 772.520 2077.260 772.780 ;
        RECT 2077.920 772.520 2078.180 772.780 ;
        RECT 2077.000 675.620 2077.260 675.880 ;
        RECT 2077.000 628.020 2077.260 628.280 ;
        RECT 2077.000 579.400 2077.260 579.660 ;
        RECT 2077.000 531.460 2077.260 531.720 ;
        RECT 2077.000 482.840 2077.260 483.100 ;
        RECT 2077.000 434.900 2077.260 435.160 ;
        RECT 2077.000 385.940 2077.260 386.200 ;
        RECT 2077.000 338.000 2077.260 338.260 ;
        RECT 2077.000 96.260 2077.260 96.520 ;
        RECT 2078.380 48.320 2078.640 48.580 ;
      LAYER met2 ;
        RECT 1713.130 1700.000 1713.410 1704.000 ;
        RECT 1713.200 1680.950 1713.340 1700.000 ;
        RECT 1713.140 1680.630 1713.400 1680.950 ;
        RECT 2077.000 1680.630 2077.260 1680.950 ;
        RECT 2077.060 1642.190 2077.200 1680.630 ;
        RECT 2077.000 1641.870 2077.260 1642.190 ;
        RECT 2077.000 1593.930 2077.260 1594.250 ;
        RECT 2077.060 1545.630 2077.200 1593.930 ;
        RECT 2077.000 1545.310 2077.260 1545.630 ;
        RECT 2077.000 1497.370 2077.260 1497.690 ;
        RECT 2077.060 1449.070 2077.200 1497.370 ;
        RECT 2077.000 1448.750 2077.260 1449.070 ;
        RECT 2077.000 1400.810 2077.260 1401.130 ;
        RECT 2077.060 1353.725 2077.200 1400.810 ;
        RECT 2076.990 1353.355 2077.270 1353.725 ;
        RECT 2076.990 1352.675 2077.270 1353.045 ;
        RECT 2077.060 1352.510 2077.200 1352.675 ;
        RECT 2077.000 1352.190 2077.260 1352.510 ;
        RECT 2077.000 1304.250 2077.260 1304.570 ;
        RECT 2077.060 1257.165 2077.200 1304.250 ;
        RECT 2076.990 1256.795 2077.270 1257.165 ;
        RECT 2076.990 1256.115 2077.270 1256.485 ;
        RECT 2077.060 1255.950 2077.200 1256.115 ;
        RECT 2077.000 1255.630 2077.260 1255.950 ;
        RECT 2077.000 1207.350 2077.260 1207.670 ;
        RECT 2077.060 1159.245 2077.200 1207.350 ;
        RECT 2076.990 1158.875 2077.270 1159.245 ;
        RECT 2077.910 1158.875 2078.190 1159.245 ;
        RECT 2077.980 1111.110 2078.120 1158.875 ;
        RECT 2077.000 1110.790 2077.260 1111.110 ;
        RECT 2077.920 1110.790 2078.180 1111.110 ;
        RECT 2077.060 1062.685 2077.200 1110.790 ;
        RECT 2076.990 1062.315 2077.270 1062.685 ;
        RECT 2077.910 1062.315 2078.190 1062.685 ;
        RECT 2077.980 1014.550 2078.120 1062.315 ;
        RECT 2077.000 1014.230 2077.260 1014.550 ;
        RECT 2077.920 1014.230 2078.180 1014.550 ;
        RECT 2077.060 966.125 2077.200 1014.230 ;
        RECT 2076.990 965.755 2077.270 966.125 ;
        RECT 2077.910 965.755 2078.190 966.125 ;
        RECT 2077.980 917.990 2078.120 965.755 ;
        RECT 2077.000 917.670 2077.260 917.990 ;
        RECT 2077.920 917.670 2078.180 917.990 ;
        RECT 2077.060 869.565 2077.200 917.670 ;
        RECT 2076.990 869.195 2077.270 869.565 ;
        RECT 2077.910 869.195 2078.190 869.565 ;
        RECT 2077.980 821.285 2078.120 869.195 ;
        RECT 2076.990 820.915 2077.270 821.285 ;
        RECT 2077.910 820.915 2078.190 821.285 ;
        RECT 2077.060 772.810 2077.200 820.915 ;
        RECT 2077.000 772.490 2077.260 772.810 ;
        RECT 2077.920 772.490 2078.180 772.810 ;
        RECT 2077.980 724.725 2078.120 772.490 ;
        RECT 2076.990 724.355 2077.270 724.725 ;
        RECT 2077.910 724.355 2078.190 724.725 ;
        RECT 2077.060 675.910 2077.200 724.355 ;
        RECT 2077.000 675.590 2077.260 675.910 ;
        RECT 2077.000 627.990 2077.260 628.310 ;
        RECT 2077.060 579.690 2077.200 627.990 ;
        RECT 2077.000 579.370 2077.260 579.690 ;
        RECT 2077.000 531.430 2077.260 531.750 ;
        RECT 2077.060 483.130 2077.200 531.430 ;
        RECT 2077.000 482.810 2077.260 483.130 ;
        RECT 2077.000 434.870 2077.260 435.190 ;
        RECT 2077.060 386.230 2077.200 434.870 ;
        RECT 2077.000 385.910 2077.260 386.230 ;
        RECT 2077.000 337.970 2077.260 338.290 ;
        RECT 2077.060 290.885 2077.200 337.970 ;
        RECT 2076.990 290.515 2077.270 290.885 ;
        RECT 2076.990 289.835 2077.270 290.205 ;
        RECT 2077.060 96.550 2077.200 289.835 ;
        RECT 2077.000 96.230 2077.260 96.550 ;
        RECT 2078.380 48.290 2078.640 48.610 ;
        RECT 2078.440 2.400 2078.580 48.290 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
      LAYER via2 ;
        RECT 2076.990 1353.400 2077.270 1353.680 ;
        RECT 2076.990 1352.720 2077.270 1353.000 ;
        RECT 2076.990 1256.840 2077.270 1257.120 ;
        RECT 2076.990 1256.160 2077.270 1256.440 ;
        RECT 2076.990 1158.920 2077.270 1159.200 ;
        RECT 2077.910 1158.920 2078.190 1159.200 ;
        RECT 2076.990 1062.360 2077.270 1062.640 ;
        RECT 2077.910 1062.360 2078.190 1062.640 ;
        RECT 2076.990 965.800 2077.270 966.080 ;
        RECT 2077.910 965.800 2078.190 966.080 ;
        RECT 2076.990 869.240 2077.270 869.520 ;
        RECT 2077.910 869.240 2078.190 869.520 ;
        RECT 2076.990 820.960 2077.270 821.240 ;
        RECT 2077.910 820.960 2078.190 821.240 ;
        RECT 2076.990 724.400 2077.270 724.680 ;
        RECT 2077.910 724.400 2078.190 724.680 ;
        RECT 2076.990 290.560 2077.270 290.840 ;
        RECT 2076.990 289.880 2077.270 290.160 ;
      LAYER met3 ;
        RECT 2076.965 1353.690 2077.295 1353.705 ;
        RECT 2076.750 1353.375 2077.295 1353.690 ;
        RECT 2076.750 1353.025 2077.050 1353.375 ;
        RECT 2076.750 1352.710 2077.295 1353.025 ;
        RECT 2076.965 1352.695 2077.295 1352.710 ;
        RECT 2076.965 1257.130 2077.295 1257.145 ;
        RECT 2076.750 1256.815 2077.295 1257.130 ;
        RECT 2076.750 1256.465 2077.050 1256.815 ;
        RECT 2076.750 1256.150 2077.295 1256.465 ;
        RECT 2076.965 1256.135 2077.295 1256.150 ;
        RECT 2076.965 1159.210 2077.295 1159.225 ;
        RECT 2077.885 1159.210 2078.215 1159.225 ;
        RECT 2076.965 1158.910 2078.215 1159.210 ;
        RECT 2076.965 1158.895 2077.295 1158.910 ;
        RECT 2077.885 1158.895 2078.215 1158.910 ;
        RECT 2076.965 1062.650 2077.295 1062.665 ;
        RECT 2077.885 1062.650 2078.215 1062.665 ;
        RECT 2076.965 1062.350 2078.215 1062.650 ;
        RECT 2076.965 1062.335 2077.295 1062.350 ;
        RECT 2077.885 1062.335 2078.215 1062.350 ;
        RECT 2076.965 966.090 2077.295 966.105 ;
        RECT 2077.885 966.090 2078.215 966.105 ;
        RECT 2076.965 965.790 2078.215 966.090 ;
        RECT 2076.965 965.775 2077.295 965.790 ;
        RECT 2077.885 965.775 2078.215 965.790 ;
        RECT 2076.965 869.530 2077.295 869.545 ;
        RECT 2077.885 869.530 2078.215 869.545 ;
        RECT 2076.965 869.230 2078.215 869.530 ;
        RECT 2076.965 869.215 2077.295 869.230 ;
        RECT 2077.885 869.215 2078.215 869.230 ;
        RECT 2076.965 821.250 2077.295 821.265 ;
        RECT 2077.885 821.250 2078.215 821.265 ;
        RECT 2076.965 820.950 2078.215 821.250 ;
        RECT 2076.965 820.935 2077.295 820.950 ;
        RECT 2077.885 820.935 2078.215 820.950 ;
        RECT 2076.965 724.690 2077.295 724.705 ;
        RECT 2077.885 724.690 2078.215 724.705 ;
        RECT 2076.965 724.390 2078.215 724.690 ;
        RECT 2076.965 724.375 2077.295 724.390 ;
        RECT 2077.885 724.375 2078.215 724.390 ;
        RECT 2076.965 290.850 2077.295 290.865 ;
        RECT 2076.750 290.535 2077.295 290.850 ;
        RECT 2076.750 290.185 2077.050 290.535 ;
        RECT 2076.750 289.870 2077.295 290.185 ;
        RECT 2076.965 289.855 2077.295 289.870 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1718.170 1685.280 1718.490 1685.340 ;
        RECT 1728.290 1685.280 1728.610 1685.340 ;
        RECT 1718.170 1685.140 1728.610 1685.280 ;
        RECT 1718.170 1685.080 1718.490 1685.140 ;
        RECT 1728.290 1685.080 1728.610 1685.140 ;
        RECT 1728.290 65.520 1728.610 65.580 ;
        RECT 2090.770 65.520 2091.090 65.580 ;
        RECT 1728.290 65.380 2091.090 65.520 ;
        RECT 1728.290 65.320 1728.610 65.380 ;
        RECT 2090.770 65.320 2091.090 65.380 ;
        RECT 2090.770 62.120 2091.090 62.180 ;
        RECT 2095.830 62.120 2096.150 62.180 ;
        RECT 2090.770 61.980 2096.150 62.120 ;
        RECT 2090.770 61.920 2091.090 61.980 ;
        RECT 2095.830 61.920 2096.150 61.980 ;
      LAYER via ;
        RECT 1718.200 1685.080 1718.460 1685.340 ;
        RECT 1728.320 1685.080 1728.580 1685.340 ;
        RECT 1728.320 65.320 1728.580 65.580 ;
        RECT 2090.800 65.320 2091.060 65.580 ;
        RECT 2090.800 61.920 2091.060 62.180 ;
        RECT 2095.860 61.920 2096.120 62.180 ;
      LAYER met2 ;
        RECT 1718.190 1700.000 1718.470 1704.000 ;
        RECT 1718.260 1685.370 1718.400 1700.000 ;
        RECT 1718.200 1685.050 1718.460 1685.370 ;
        RECT 1728.320 1685.050 1728.580 1685.370 ;
        RECT 1728.380 65.610 1728.520 1685.050 ;
        RECT 1728.320 65.290 1728.580 65.610 ;
        RECT 2090.800 65.290 2091.060 65.610 ;
        RECT 2090.860 62.210 2091.000 65.290 ;
        RECT 2090.800 61.890 2091.060 62.210 ;
        RECT 2095.860 61.890 2096.120 62.210 ;
        RECT 2095.920 2.400 2096.060 61.890 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 0.300 ;
=======
      LAYER met1 ;
        RECT 1722.770 1683.920 1723.090 1683.980 ;
        RECT 1724.150 1683.920 1724.470 1683.980 ;
        RECT 1722.770 1683.780 1724.470 1683.920 ;
        RECT 1722.770 1683.720 1723.090 1683.780 ;
        RECT 1724.150 1683.720 1724.470 1683.780 ;
        RECT 1724.150 27.780 1724.470 27.840 ;
        RECT 2113.770 27.780 2114.090 27.840 ;
        RECT 1724.150 27.640 2114.090 27.780 ;
        RECT 1724.150 27.580 1724.470 27.640 ;
        RECT 2113.770 27.580 2114.090 27.640 ;
      LAYER via ;
        RECT 1722.800 1683.720 1723.060 1683.980 ;
        RECT 1724.180 1683.720 1724.440 1683.980 ;
        RECT 1724.180 27.580 1724.440 27.840 ;
        RECT 2113.800 27.580 2114.060 27.840 ;
      LAYER met2 ;
        RECT 1722.790 1700.000 1723.070 1704.000 ;
        RECT 1722.860 1684.010 1723.000 1700.000 ;
        RECT 1722.800 1683.690 1723.060 1684.010 ;
        RECT 1724.180 1683.690 1724.440 1684.010 ;
        RECT 1724.240 27.870 1724.380 1683.690 ;
        RECT 1724.180 27.550 1724.440 27.870 ;
        RECT 2113.800 27.550 2114.060 27.870 ;
        RECT 2113.860 2.400 2114.000 27.550 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 0.300 ;
=======
      LAYER met1 ;
        RECT 1727.830 1683.920 1728.150 1683.980 ;
        RECT 1731.050 1683.920 1731.370 1683.980 ;
        RECT 1727.830 1683.780 1731.370 1683.920 ;
        RECT 1727.830 1683.720 1728.150 1683.780 ;
        RECT 1731.050 1683.720 1731.370 1683.780 ;
        RECT 1731.050 28.120 1731.370 28.180 ;
        RECT 2131.710 28.120 2132.030 28.180 ;
        RECT 1731.050 27.980 2132.030 28.120 ;
        RECT 1731.050 27.920 1731.370 27.980 ;
        RECT 2131.710 27.920 2132.030 27.980 ;
      LAYER via ;
        RECT 1727.860 1683.720 1728.120 1683.980 ;
        RECT 1731.080 1683.720 1731.340 1683.980 ;
        RECT 1731.080 27.920 1731.340 28.180 ;
        RECT 2131.740 27.920 2132.000 28.180 ;
      LAYER met2 ;
        RECT 1727.850 1700.000 1728.130 1704.000 ;
        RECT 1727.920 1684.010 1728.060 1700.000 ;
        RECT 1727.860 1683.690 1728.120 1684.010 ;
        RECT 1731.080 1683.690 1731.340 1684.010 ;
        RECT 1731.140 28.210 1731.280 1683.690 ;
        RECT 1731.080 27.890 1731.340 28.210 ;
        RECT 2131.740 27.890 2132.000 28.210 ;
        RECT 2131.800 2.400 2131.940 27.890 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1732.430 1684.260 1732.750 1684.320 ;
        RECT 1738.410 1684.260 1738.730 1684.320 ;
        RECT 1732.430 1684.120 1738.730 1684.260 ;
        RECT 1732.430 1684.060 1732.750 1684.120 ;
        RECT 1738.410 1684.060 1738.730 1684.120 ;
        RECT 1738.410 28.460 1738.730 28.520 ;
        RECT 2149.650 28.460 2149.970 28.520 ;
        RECT 1738.410 28.320 2149.970 28.460 ;
        RECT 1738.410 28.260 1738.730 28.320 ;
        RECT 2149.650 28.260 2149.970 28.320 ;
      LAYER via ;
        RECT 1732.460 1684.060 1732.720 1684.320 ;
        RECT 1738.440 1684.060 1738.700 1684.320 ;
        RECT 1738.440 28.260 1738.700 28.520 ;
        RECT 2149.680 28.260 2149.940 28.520 ;
      LAYER met2 ;
        RECT 1732.450 1700.000 1732.730 1704.000 ;
        RECT 1732.520 1684.350 1732.660 1700.000 ;
        RECT 1732.460 1684.030 1732.720 1684.350 ;
        RECT 1738.440 1684.030 1738.700 1684.350 ;
        RECT 1738.500 28.550 1738.640 1684.030 ;
        RECT 1738.440 28.230 1738.700 28.550 ;
        RECT 2149.680 28.230 2149.940 28.550 ;
        RECT 2149.740 2.400 2149.880 28.230 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1737.950 28.800 1738.270 28.860 ;
        RECT 2167.590 28.800 2167.910 28.860 ;
        RECT 1737.950 28.660 2167.910 28.800 ;
        RECT 1737.950 28.600 1738.270 28.660 ;
        RECT 2167.590 28.600 2167.910 28.660 ;
      LAYER via ;
        RECT 1737.980 28.600 1738.240 28.860 ;
        RECT 2167.620 28.600 2167.880 28.860 ;
      LAYER met2 ;
        RECT 1737.510 1700.410 1737.790 1704.000 ;
        RECT 1737.510 1700.270 1738.180 1700.410 ;
        RECT 1737.510 1700.000 1737.790 1700.270 ;
        RECT 1738.040 28.890 1738.180 1700.270 ;
        RECT 1737.980 28.570 1738.240 28.890 ;
        RECT 2167.620 28.570 2167.880 28.890 ;
        RECT 2167.680 2.400 2167.820 28.570 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 0.300 ;
=======
      LAYER met1 ;
        RECT 1742.090 1683.920 1742.410 1683.980 ;
        RECT 1744.850 1683.920 1745.170 1683.980 ;
        RECT 1742.090 1683.780 1745.170 1683.920 ;
        RECT 1742.090 1683.720 1742.410 1683.780 ;
        RECT 1744.850 1683.720 1745.170 1683.780 ;
        RECT 1744.850 29.140 1745.170 29.200 ;
        RECT 2185.070 29.140 2185.390 29.200 ;
        RECT 1744.850 29.000 2185.390 29.140 ;
        RECT 1744.850 28.940 1745.170 29.000 ;
        RECT 2185.070 28.940 2185.390 29.000 ;
      LAYER via ;
        RECT 1742.120 1683.720 1742.380 1683.980 ;
        RECT 1744.880 1683.720 1745.140 1683.980 ;
        RECT 1744.880 28.940 1745.140 29.200 ;
        RECT 2185.100 28.940 2185.360 29.200 ;
      LAYER met2 ;
        RECT 1742.110 1700.000 1742.390 1704.000 ;
        RECT 1742.180 1684.010 1742.320 1700.000 ;
        RECT 1742.120 1683.690 1742.380 1684.010 ;
        RECT 1744.880 1683.690 1745.140 1684.010 ;
        RECT 1744.940 29.230 1745.080 1683.690 ;
        RECT 1744.880 28.910 1745.140 29.230 ;
        RECT 2185.100 28.910 2185.360 29.230 ;
        RECT 2185.160 2.400 2185.300 28.910 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1747.150 1684.260 1747.470 1684.320 ;
        RECT 1751.750 1684.260 1752.070 1684.320 ;
        RECT 1747.150 1684.120 1752.070 1684.260 ;
        RECT 1747.150 1684.060 1747.470 1684.120 ;
        RECT 1751.750 1684.060 1752.070 1684.120 ;
        RECT 1751.750 29.480 1752.070 29.540 ;
        RECT 2203.010 29.480 2203.330 29.540 ;
        RECT 1751.750 29.340 2203.330 29.480 ;
        RECT 1751.750 29.280 1752.070 29.340 ;
        RECT 2203.010 29.280 2203.330 29.340 ;
      LAYER via ;
        RECT 1747.180 1684.060 1747.440 1684.320 ;
        RECT 1751.780 1684.060 1752.040 1684.320 ;
        RECT 1751.780 29.280 1752.040 29.540 ;
        RECT 2203.040 29.280 2203.300 29.540 ;
      LAYER met2 ;
        RECT 1747.170 1700.000 1747.450 1704.000 ;
        RECT 1747.240 1684.350 1747.380 1700.000 ;
        RECT 1747.180 1684.030 1747.440 1684.350 ;
        RECT 1751.780 1684.030 1752.040 1684.350 ;
        RECT 1751.840 29.570 1751.980 1684.030 ;
        RECT 1751.780 29.250 1752.040 29.570 ;
        RECT 2203.040 29.250 2203.300 29.570 ;
        RECT 2203.100 2.400 2203.240 29.250 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1751.290 29.820 1751.610 29.880 ;
        RECT 2220.950 29.820 2221.270 29.880 ;
        RECT 1751.290 29.680 2221.270 29.820 ;
        RECT 1751.290 29.620 1751.610 29.680 ;
        RECT 2220.950 29.620 2221.270 29.680 ;
      LAYER via ;
        RECT 1751.320 29.620 1751.580 29.880 ;
        RECT 2220.980 29.620 2221.240 29.880 ;
      LAYER met2 ;
        RECT 1751.770 1700.410 1752.050 1704.000 ;
        RECT 1751.380 1700.270 1752.050 1700.410 ;
        RECT 1751.380 29.910 1751.520 1700.270 ;
        RECT 1751.770 1700.000 1752.050 1700.270 ;
        RECT 1751.320 29.590 1751.580 29.910 ;
        RECT 2220.980 29.590 2221.240 29.910 ;
        RECT 2221.040 2.400 2221.180 29.590 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 0.300 ;
=======
      LAYER li1 ;
        RECT 1354.385 1607.605 1354.555 1642.115 ;
        RECT 1354.385 1545.725 1354.555 1593.835 ;
        RECT 1354.385 1400.885 1354.555 1414.995 ;
        RECT 1354.385 1207.425 1354.555 1255.875 ;
        RECT 1354.385 1062.585 1354.555 1110.695 ;
        RECT 1354.385 821.185 1354.555 910.775 ;
        RECT 1354.385 766.105 1354.555 814.215 ;
        RECT 1354.385 524.365 1354.555 572.475 ;
        RECT 1354.845 469.285 1355.015 517.395 ;
      LAYER mcon ;
        RECT 1354.385 1641.945 1354.555 1642.115 ;
        RECT 1354.385 1593.665 1354.555 1593.835 ;
        RECT 1354.385 1414.825 1354.555 1414.995 ;
        RECT 1354.385 1255.705 1354.555 1255.875 ;
        RECT 1354.385 1110.525 1354.555 1110.695 ;
        RECT 1354.385 910.605 1354.555 910.775 ;
        RECT 1354.385 814.045 1354.555 814.215 ;
        RECT 1354.385 572.305 1354.555 572.475 ;
        RECT 1354.845 517.225 1355.015 517.395 ;
      LAYER met1 ;
        RECT 1354.310 1642.100 1354.630 1642.160 ;
        RECT 1354.115 1641.960 1354.630 1642.100 ;
        RECT 1354.310 1641.900 1354.630 1641.960 ;
        RECT 1354.310 1607.760 1354.630 1607.820 ;
        RECT 1354.115 1607.620 1354.630 1607.760 ;
        RECT 1354.310 1607.560 1354.630 1607.620 ;
        RECT 1354.310 1593.820 1354.630 1593.880 ;
        RECT 1354.115 1593.680 1354.630 1593.820 ;
        RECT 1354.310 1593.620 1354.630 1593.680 ;
        RECT 1354.325 1545.880 1354.615 1545.925 ;
        RECT 1354.770 1545.880 1355.090 1545.940 ;
        RECT 1354.325 1545.740 1355.090 1545.880 ;
        RECT 1354.325 1545.695 1354.615 1545.740 ;
        RECT 1354.770 1545.680 1355.090 1545.740 ;
        RECT 1354.325 1414.980 1354.615 1415.025 ;
        RECT 1354.770 1414.980 1355.090 1415.040 ;
        RECT 1354.325 1414.840 1355.090 1414.980 ;
        RECT 1354.325 1414.795 1354.615 1414.840 ;
        RECT 1354.770 1414.780 1355.090 1414.840 ;
        RECT 1354.310 1401.040 1354.630 1401.100 ;
        RECT 1354.115 1400.900 1354.630 1401.040 ;
        RECT 1354.310 1400.840 1354.630 1400.900 ;
        RECT 1354.770 1304.820 1355.090 1304.880 ;
        RECT 1354.400 1304.680 1355.090 1304.820 ;
        RECT 1354.400 1304.540 1354.540 1304.680 ;
        RECT 1354.770 1304.620 1355.090 1304.680 ;
        RECT 1354.310 1304.280 1354.630 1304.540 ;
        RECT 1354.310 1255.860 1354.630 1255.920 ;
        RECT 1354.115 1255.720 1354.630 1255.860 ;
        RECT 1354.310 1255.660 1354.630 1255.720 ;
        RECT 1354.310 1207.580 1354.630 1207.640 ;
        RECT 1354.115 1207.440 1354.630 1207.580 ;
        RECT 1354.310 1207.380 1354.630 1207.440 ;
        RECT 1354.310 1110.680 1354.630 1110.740 ;
        RECT 1354.115 1110.540 1354.630 1110.680 ;
        RECT 1354.310 1110.480 1354.630 1110.540 ;
        RECT 1354.325 1062.740 1354.615 1062.785 ;
        RECT 1354.770 1062.740 1355.090 1062.800 ;
        RECT 1354.325 1062.600 1355.090 1062.740 ;
        RECT 1354.325 1062.555 1354.615 1062.600 ;
        RECT 1354.770 1062.540 1355.090 1062.600 ;
        RECT 1354.310 918.240 1354.630 918.300 ;
        RECT 1354.770 918.240 1355.090 918.300 ;
        RECT 1354.310 918.100 1355.090 918.240 ;
        RECT 1354.310 918.040 1354.630 918.100 ;
        RECT 1354.770 918.040 1355.090 918.100 ;
        RECT 1354.310 910.760 1354.630 910.820 ;
        RECT 1354.115 910.620 1354.630 910.760 ;
        RECT 1354.310 910.560 1354.630 910.620 ;
        RECT 1354.310 821.340 1354.630 821.400 ;
        RECT 1354.115 821.200 1354.630 821.340 ;
        RECT 1354.310 821.140 1354.630 821.200 ;
        RECT 1354.310 814.200 1354.630 814.260 ;
        RECT 1354.115 814.060 1354.630 814.200 ;
        RECT 1354.310 814.000 1354.630 814.060 ;
        RECT 1354.310 766.260 1354.630 766.320 ;
        RECT 1354.115 766.120 1354.630 766.260 ;
        RECT 1354.310 766.060 1354.630 766.120 ;
        RECT 1354.310 765.580 1354.630 765.640 ;
        RECT 1355.230 765.580 1355.550 765.640 ;
        RECT 1354.310 765.440 1355.550 765.580 ;
        RECT 1354.310 765.380 1354.630 765.440 ;
        RECT 1355.230 765.380 1355.550 765.440 ;
        RECT 1354.310 717.640 1354.630 717.700 ;
        RECT 1354.770 717.640 1355.090 717.700 ;
        RECT 1354.310 717.500 1355.090 717.640 ;
        RECT 1354.310 717.440 1354.630 717.500 ;
        RECT 1354.770 717.440 1355.090 717.500 ;
        RECT 1354.310 572.460 1354.630 572.520 ;
        RECT 1354.115 572.320 1354.630 572.460 ;
        RECT 1354.310 572.260 1354.630 572.320 ;
        RECT 1354.325 524.520 1354.615 524.565 ;
        RECT 1354.770 524.520 1355.090 524.580 ;
        RECT 1354.325 524.380 1355.090 524.520 ;
        RECT 1354.325 524.335 1354.615 524.380 ;
        RECT 1354.770 524.320 1355.090 524.380 ;
        RECT 1354.770 517.380 1355.090 517.440 ;
        RECT 1354.575 517.240 1355.090 517.380 ;
        RECT 1354.770 517.180 1355.090 517.240 ;
        RECT 1354.770 469.440 1355.090 469.500 ;
        RECT 1354.575 469.300 1355.090 469.440 ;
        RECT 1354.770 469.240 1355.090 469.300 ;
        RECT 1354.310 427.960 1354.630 428.020 ;
        RECT 1354.770 427.960 1355.090 428.020 ;
        RECT 1354.310 427.820 1355.090 427.960 ;
        RECT 1354.310 427.760 1354.630 427.820 ;
        RECT 1354.770 427.760 1355.090 427.820 ;
        RECT 1354.310 283.120 1354.630 283.180 ;
        RECT 1354.770 283.120 1355.090 283.180 ;
        RECT 1354.310 282.980 1355.090 283.120 ;
        RECT 1354.310 282.920 1354.630 282.980 ;
        RECT 1354.770 282.920 1355.090 282.980 ;
        RECT 775.630 31.520 775.950 31.580 ;
        RECT 1354.770 31.520 1355.090 31.580 ;
        RECT 775.630 31.380 1355.090 31.520 ;
        RECT 775.630 31.320 775.950 31.380 ;
        RECT 1354.770 31.320 1355.090 31.380 ;
      LAYER via ;
        RECT 1354.340 1641.900 1354.600 1642.160 ;
        RECT 1354.340 1607.560 1354.600 1607.820 ;
        RECT 1354.340 1593.620 1354.600 1593.880 ;
        RECT 1354.800 1545.680 1355.060 1545.940 ;
        RECT 1354.800 1414.780 1355.060 1415.040 ;
        RECT 1354.340 1400.840 1354.600 1401.100 ;
        RECT 1354.800 1304.620 1355.060 1304.880 ;
        RECT 1354.340 1304.280 1354.600 1304.540 ;
        RECT 1354.340 1255.660 1354.600 1255.920 ;
        RECT 1354.340 1207.380 1354.600 1207.640 ;
        RECT 1354.340 1110.480 1354.600 1110.740 ;
        RECT 1354.800 1062.540 1355.060 1062.800 ;
        RECT 1354.340 918.040 1354.600 918.300 ;
        RECT 1354.800 918.040 1355.060 918.300 ;
        RECT 1354.340 910.560 1354.600 910.820 ;
        RECT 1354.340 821.140 1354.600 821.400 ;
        RECT 1354.340 814.000 1354.600 814.260 ;
        RECT 1354.340 766.060 1354.600 766.320 ;
        RECT 1354.340 765.380 1354.600 765.640 ;
        RECT 1355.260 765.380 1355.520 765.640 ;
        RECT 1354.340 717.440 1354.600 717.700 ;
        RECT 1354.800 717.440 1355.060 717.700 ;
        RECT 1354.340 572.260 1354.600 572.520 ;
        RECT 1354.800 524.320 1355.060 524.580 ;
        RECT 1354.800 517.180 1355.060 517.440 ;
        RECT 1354.800 469.240 1355.060 469.500 ;
        RECT 1354.340 427.760 1354.600 428.020 ;
        RECT 1354.800 427.760 1355.060 428.020 ;
        RECT 1354.340 282.920 1354.600 283.180 ;
        RECT 1354.800 282.920 1355.060 283.180 ;
        RECT 775.660 31.320 775.920 31.580 ;
        RECT 1354.800 31.320 1355.060 31.580 ;
      LAYER met2 ;
        RECT 1358.930 1700.410 1359.210 1704.000 ;
        RECT 1358.540 1700.270 1359.210 1700.410 ;
        RECT 1358.540 1676.610 1358.680 1700.270 ;
        RECT 1358.930 1700.000 1359.210 1700.270 ;
        RECT 1354.400 1676.470 1358.680 1676.610 ;
        RECT 1354.400 1642.190 1354.540 1676.470 ;
        RECT 1354.340 1641.870 1354.600 1642.190 ;
        RECT 1354.340 1607.530 1354.600 1607.850 ;
        RECT 1354.400 1593.910 1354.540 1607.530 ;
        RECT 1354.340 1593.590 1354.600 1593.910 ;
        RECT 1354.800 1545.650 1355.060 1545.970 ;
        RECT 1354.860 1415.070 1355.000 1545.650 ;
        RECT 1354.800 1414.750 1355.060 1415.070 ;
        RECT 1354.340 1400.810 1354.600 1401.130 ;
        RECT 1354.400 1352.250 1354.540 1400.810 ;
        RECT 1354.400 1352.110 1355.000 1352.250 ;
        RECT 1354.860 1304.910 1355.000 1352.110 ;
        RECT 1354.800 1304.590 1355.060 1304.910 ;
        RECT 1354.340 1304.250 1354.600 1304.570 ;
        RECT 1354.400 1255.950 1354.540 1304.250 ;
        RECT 1354.340 1255.630 1354.600 1255.950 ;
        RECT 1354.340 1207.350 1354.600 1207.670 ;
        RECT 1354.400 1110.770 1354.540 1207.350 ;
        RECT 1354.340 1110.450 1354.600 1110.770 ;
        RECT 1354.800 1062.510 1355.060 1062.830 ;
        RECT 1354.860 918.330 1355.000 1062.510 ;
        RECT 1354.340 918.010 1354.600 918.330 ;
        RECT 1354.800 918.010 1355.060 918.330 ;
        RECT 1354.400 910.850 1354.540 918.010 ;
        RECT 1354.340 910.530 1354.600 910.850 ;
        RECT 1354.340 821.110 1354.600 821.430 ;
        RECT 1354.400 814.290 1354.540 821.110 ;
        RECT 1354.340 813.970 1354.600 814.290 ;
        RECT 1354.340 766.030 1354.600 766.350 ;
        RECT 1354.400 765.670 1354.540 766.030 ;
        RECT 1354.340 765.350 1354.600 765.670 ;
        RECT 1355.260 765.350 1355.520 765.670 ;
        RECT 1355.320 717.925 1355.460 765.350 ;
        RECT 1354.330 717.555 1354.610 717.925 ;
        RECT 1354.340 717.410 1354.600 717.555 ;
        RECT 1354.800 717.410 1355.060 717.730 ;
        RECT 1355.250 717.555 1355.530 717.925 ;
        RECT 1354.860 671.005 1355.000 717.410 ;
        RECT 1354.790 670.635 1355.070 671.005 ;
        RECT 1354.330 669.275 1354.610 669.645 ;
        RECT 1354.400 572.550 1354.540 669.275 ;
        RECT 1354.340 572.230 1354.600 572.550 ;
        RECT 1354.800 524.290 1355.060 524.610 ;
        RECT 1354.860 517.470 1355.000 524.290 ;
        RECT 1354.800 517.150 1355.060 517.470 ;
        RECT 1354.800 469.210 1355.060 469.530 ;
        RECT 1354.860 428.050 1355.000 469.210 ;
        RECT 1354.340 427.730 1354.600 428.050 ;
        RECT 1354.800 427.730 1355.060 428.050 ;
        RECT 1354.400 283.210 1354.540 427.730 ;
        RECT 1354.340 282.890 1354.600 283.210 ;
        RECT 1354.800 282.890 1355.060 283.210 ;
        RECT 1354.860 207.130 1355.000 282.890 ;
        RECT 1354.400 206.990 1355.000 207.130 ;
        RECT 1354.400 144.685 1354.540 206.990 ;
        RECT 1354.330 144.315 1354.610 144.685 ;
        RECT 1354.790 143.635 1355.070 144.005 ;
        RECT 1354.860 31.610 1355.000 143.635 ;
        RECT 775.660 31.290 775.920 31.610 ;
        RECT 1354.800 31.290 1355.060 31.610 ;
        RECT 775.720 2.400 775.860 31.290 ;
        RECT 775.510 -4.800 776.070 2.400 ;
      LAYER via2 ;
        RECT 1354.330 717.600 1354.610 717.880 ;
        RECT 1355.250 717.600 1355.530 717.880 ;
        RECT 1354.790 670.680 1355.070 670.960 ;
        RECT 1354.330 669.320 1354.610 669.600 ;
        RECT 1354.330 144.360 1354.610 144.640 ;
        RECT 1354.790 143.680 1355.070 143.960 ;
      LAYER met3 ;
        RECT 1354.305 717.890 1354.635 717.905 ;
        RECT 1355.225 717.890 1355.555 717.905 ;
        RECT 1354.305 717.590 1355.555 717.890 ;
        RECT 1354.305 717.575 1354.635 717.590 ;
        RECT 1355.225 717.575 1355.555 717.590 ;
        RECT 1354.765 670.970 1355.095 670.985 ;
        RECT 1353.630 670.670 1355.095 670.970 ;
        RECT 1353.630 669.610 1353.930 670.670 ;
        RECT 1354.765 670.655 1355.095 670.670 ;
        RECT 1354.305 669.610 1354.635 669.625 ;
        RECT 1353.630 669.310 1354.635 669.610 ;
        RECT 1354.305 669.295 1354.635 669.310 ;
        RECT 1354.305 144.650 1354.635 144.665 ;
        RECT 1353.630 144.350 1354.635 144.650 ;
        RECT 1353.630 143.970 1353.930 144.350 ;
        RECT 1354.305 144.335 1354.635 144.350 ;
        RECT 1354.765 143.970 1355.095 143.985 ;
        RECT 1353.630 143.670 1355.095 143.970 ;
        RECT 1354.765 143.655 1355.095 143.670 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 779.310 1597.560 779.630 1597.620 ;
        RECT 1360.290 1597.560 1360.610 1597.620 ;
        RECT 779.310 1597.420 1360.610 1597.560 ;
        RECT 779.310 1597.360 779.630 1597.420 ;
        RECT 1360.290 1597.360 1360.610 1597.420 ;
        RECT 775.630 2.960 775.950 3.020 ;
        RECT 779.310 2.960 779.630 3.020 ;
        RECT 775.630 2.820 779.630 2.960 ;
        RECT 775.630 2.760 775.950 2.820 ;
        RECT 779.310 2.760 779.630 2.820 ;
      LAYER via ;
        RECT 779.340 1597.360 779.600 1597.620 ;
        RECT 1360.320 1597.360 1360.580 1597.620 ;
        RECT 775.660 2.760 775.920 3.020 ;
        RECT 779.340 2.760 779.600 3.020 ;
      LAYER met2 ;
        RECT 1359.850 1700.410 1360.130 1704.000 ;
        RECT 1359.850 1700.270 1360.520 1700.410 ;
        RECT 1359.850 1700.000 1360.130 1700.270 ;
        RECT 1360.380 1597.650 1360.520 1700.270 ;
        RECT 779.340 1597.330 779.600 1597.650 ;
        RECT 1360.320 1597.330 1360.580 1597.650 ;
        RECT 779.400 3.050 779.540 1597.330 ;
        RECT 775.660 2.730 775.920 3.050 ;
        RECT 779.340 2.730 779.600 3.050 ;
        RECT 775.720 2.400 775.860 2.730 ;
        RECT 775.510 -4.800 776.070 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1756.810 1683.920 1757.130 1683.980 ;
        RECT 1759.110 1683.920 1759.430 1683.980 ;
        RECT 1756.810 1683.780 1759.430 1683.920 ;
        RECT 1756.810 1683.720 1757.130 1683.780 ;
        RECT 1759.110 1683.720 1759.430 1683.780 ;
        RECT 1759.110 30.160 1759.430 30.220 ;
        RECT 2238.890 30.160 2239.210 30.220 ;
        RECT 1759.110 30.020 2239.210 30.160 ;
        RECT 1759.110 29.960 1759.430 30.020 ;
        RECT 2238.890 29.960 2239.210 30.020 ;
      LAYER via ;
        RECT 1756.840 1683.720 1757.100 1683.980 ;
        RECT 1759.140 1683.720 1759.400 1683.980 ;
        RECT 1759.140 29.960 1759.400 30.220 ;
        RECT 2238.920 29.960 2239.180 30.220 ;
      LAYER met2 ;
        RECT 1756.830 1700.000 1757.110 1704.000 ;
        RECT 1756.900 1684.010 1757.040 1700.000 ;
        RECT 1756.840 1683.690 1757.100 1684.010 ;
        RECT 1759.140 1683.690 1759.400 1684.010 ;
        RECT 1759.200 30.250 1759.340 1683.690 ;
        RECT 1759.140 29.930 1759.400 30.250 ;
        RECT 2238.920 29.930 2239.180 30.250 ;
        RECT 2238.980 2.400 2239.120 29.930 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1761.410 1683.920 1761.730 1683.980 ;
        RECT 1765.550 1683.920 1765.870 1683.980 ;
        RECT 1761.410 1683.780 1765.870 1683.920 ;
        RECT 1761.410 1683.720 1761.730 1683.780 ;
        RECT 1765.550 1683.720 1765.870 1683.780 ;
        RECT 1765.550 30.500 1765.870 30.560 ;
        RECT 2256.830 30.500 2257.150 30.560 ;
        RECT 1765.550 30.360 2257.150 30.500 ;
        RECT 1765.550 30.300 1765.870 30.360 ;
        RECT 2256.830 30.300 2257.150 30.360 ;
      LAYER via ;
        RECT 1761.440 1683.720 1761.700 1683.980 ;
        RECT 1765.580 1683.720 1765.840 1683.980 ;
        RECT 1765.580 30.300 1765.840 30.560 ;
        RECT 2256.860 30.300 2257.120 30.560 ;
      LAYER met2 ;
        RECT 1761.430 1700.000 1761.710 1704.000 ;
        RECT 1761.500 1684.010 1761.640 1700.000 ;
        RECT 1761.440 1683.690 1761.700 1684.010 ;
        RECT 1765.580 1683.690 1765.840 1684.010 ;
        RECT 1765.640 30.590 1765.780 1683.690 ;
        RECT 1765.580 30.270 1765.840 30.590 ;
        RECT 2256.860 30.270 2257.120 30.590 ;
        RECT 2256.920 5.170 2257.060 30.270 ;
        RECT 2256.460 5.030 2257.060 5.170 ;
        RECT 2256.460 2.400 2256.600 5.030 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1766.470 1683.920 1766.790 1683.980 ;
        RECT 1771.990 1683.920 1772.310 1683.980 ;
        RECT 1766.470 1683.780 1772.310 1683.920 ;
        RECT 1766.470 1683.720 1766.790 1683.780 ;
        RECT 1771.990 1683.720 1772.310 1683.780 ;
        RECT 1771.990 34.240 1772.310 34.300 ;
        RECT 2274.310 34.240 2274.630 34.300 ;
        RECT 1771.990 34.100 2274.630 34.240 ;
        RECT 1771.990 34.040 1772.310 34.100 ;
        RECT 2274.310 34.040 2274.630 34.100 ;
      LAYER via ;
        RECT 1766.500 1683.720 1766.760 1683.980 ;
        RECT 1772.020 1683.720 1772.280 1683.980 ;
        RECT 1772.020 34.040 1772.280 34.300 ;
        RECT 2274.340 34.040 2274.600 34.300 ;
      LAYER met2 ;
        RECT 1766.490 1700.000 1766.770 1704.000 ;
        RECT 1766.560 1684.010 1766.700 1700.000 ;
        RECT 1766.500 1683.690 1766.760 1684.010 ;
        RECT 1772.020 1683.690 1772.280 1684.010 ;
        RECT 1772.080 34.330 1772.220 1683.690 ;
        RECT 1772.020 34.010 1772.280 34.330 ;
        RECT 2274.340 34.010 2274.600 34.330 ;
        RECT 2274.400 2.400 2274.540 34.010 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1772.450 33.900 1772.770 33.960 ;
        RECT 2292.250 33.900 2292.570 33.960 ;
        RECT 1772.450 33.760 2292.570 33.900 ;
        RECT 1772.450 33.700 1772.770 33.760 ;
        RECT 2292.250 33.700 2292.570 33.760 ;
      LAYER via ;
        RECT 1772.480 33.700 1772.740 33.960 ;
        RECT 2292.280 33.700 2292.540 33.960 ;
      LAYER met2 ;
        RECT 1771.090 1700.410 1771.370 1704.000 ;
        RECT 1771.090 1700.270 1772.680 1700.410 ;
        RECT 1771.090 1700.000 1771.370 1700.270 ;
        RECT 1772.540 33.990 1772.680 1700.270 ;
        RECT 1772.480 33.670 1772.740 33.990 ;
        RECT 2292.280 33.670 2292.540 33.990 ;
        RECT 2292.340 2.400 2292.480 33.670 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 0.300 ;
=======
      LAYER met1 ;
        RECT 1776.130 1683.920 1776.450 1683.980 ;
        RECT 1779.350 1683.920 1779.670 1683.980 ;
        RECT 1776.130 1683.780 1779.670 1683.920 ;
        RECT 1776.130 1683.720 1776.450 1683.780 ;
        RECT 1779.350 1683.720 1779.670 1683.780 ;
        RECT 1779.350 33.560 1779.670 33.620 ;
        RECT 2310.190 33.560 2310.510 33.620 ;
        RECT 1779.350 33.420 2310.510 33.560 ;
        RECT 1779.350 33.360 1779.670 33.420 ;
        RECT 2310.190 33.360 2310.510 33.420 ;
      LAYER via ;
        RECT 1776.160 1683.720 1776.420 1683.980 ;
        RECT 1779.380 1683.720 1779.640 1683.980 ;
        RECT 1779.380 33.360 1779.640 33.620 ;
        RECT 2310.220 33.360 2310.480 33.620 ;
      LAYER met2 ;
        RECT 1776.150 1700.000 1776.430 1704.000 ;
        RECT 1776.220 1684.010 1776.360 1700.000 ;
        RECT 1776.160 1683.690 1776.420 1684.010 ;
        RECT 1779.380 1683.690 1779.640 1684.010 ;
        RECT 1779.440 33.650 1779.580 1683.690 ;
        RECT 1779.380 33.330 1779.640 33.650 ;
        RECT 2310.220 33.330 2310.480 33.650 ;
        RECT 2310.280 2.400 2310.420 33.330 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1780.730 1684.600 1781.050 1684.660 ;
        RECT 1786.250 1684.600 1786.570 1684.660 ;
        RECT 1780.730 1684.460 1786.570 1684.600 ;
        RECT 1780.730 1684.400 1781.050 1684.460 ;
        RECT 1786.250 1684.400 1786.570 1684.460 ;
        RECT 1786.250 33.220 1786.570 33.280 ;
        RECT 2328.130 33.220 2328.450 33.280 ;
        RECT 1786.250 33.080 2328.450 33.220 ;
        RECT 1786.250 33.020 1786.570 33.080 ;
        RECT 2328.130 33.020 2328.450 33.080 ;
      LAYER via ;
        RECT 1780.760 1684.400 1781.020 1684.660 ;
        RECT 1786.280 1684.400 1786.540 1684.660 ;
        RECT 1786.280 33.020 1786.540 33.280 ;
        RECT 2328.160 33.020 2328.420 33.280 ;
      LAYER met2 ;
        RECT 1780.750 1700.000 1781.030 1704.000 ;
        RECT 1780.820 1684.690 1780.960 1700.000 ;
        RECT 1780.760 1684.370 1781.020 1684.690 ;
        RECT 1786.280 1684.370 1786.540 1684.690 ;
        RECT 1786.340 33.310 1786.480 1684.370 ;
        RECT 1786.280 32.990 1786.540 33.310 ;
        RECT 2328.160 32.990 2328.420 33.310 ;
        RECT 2328.220 2.400 2328.360 32.990 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1786.710 32.880 1787.030 32.940 ;
        RECT 2345.610 32.880 2345.930 32.940 ;
        RECT 1786.710 32.740 2345.930 32.880 ;
        RECT 1786.710 32.680 1787.030 32.740 ;
        RECT 2345.610 32.680 2345.930 32.740 ;
      LAYER via ;
        RECT 1786.740 32.680 1787.000 32.940 ;
        RECT 2345.640 32.680 2345.900 32.940 ;
      LAYER met2 ;
        RECT 1785.810 1700.410 1786.090 1704.000 ;
        RECT 1785.810 1700.270 1786.940 1700.410 ;
        RECT 1785.810 1700.000 1786.090 1700.270 ;
        RECT 1786.800 32.970 1786.940 1700.270 ;
        RECT 1786.740 32.650 1787.000 32.970 ;
        RECT 2345.640 32.650 2345.900 32.970 ;
        RECT 2345.700 2.400 2345.840 32.650 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1790.390 1683.920 1790.710 1683.980 ;
        RECT 1793.150 1683.920 1793.470 1683.980 ;
        RECT 1790.390 1683.780 1793.470 1683.920 ;
        RECT 1790.390 1683.720 1790.710 1683.780 ;
        RECT 1793.150 1683.720 1793.470 1683.780 ;
        RECT 1793.150 32.540 1793.470 32.600 ;
        RECT 2363.550 32.540 2363.870 32.600 ;
        RECT 1793.150 32.400 2363.870 32.540 ;
        RECT 1793.150 32.340 1793.470 32.400 ;
        RECT 2363.550 32.340 2363.870 32.400 ;
      LAYER via ;
        RECT 1790.420 1683.720 1790.680 1683.980 ;
        RECT 1793.180 1683.720 1793.440 1683.980 ;
        RECT 1793.180 32.340 1793.440 32.600 ;
        RECT 2363.580 32.340 2363.840 32.600 ;
      LAYER met2 ;
        RECT 1790.410 1700.000 1790.690 1704.000 ;
        RECT 1790.480 1684.010 1790.620 1700.000 ;
        RECT 1790.420 1683.690 1790.680 1684.010 ;
        RECT 1793.180 1683.690 1793.440 1684.010 ;
        RECT 1793.240 32.630 1793.380 1683.690 ;
        RECT 1793.180 32.310 1793.440 32.630 ;
        RECT 2363.580 32.310 2363.840 32.630 ;
        RECT 2363.640 2.400 2363.780 32.310 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1795.450 1684.600 1795.770 1684.660 ;
        RECT 1800.050 1684.600 1800.370 1684.660 ;
        RECT 1795.450 1684.460 1800.370 1684.600 ;
        RECT 1795.450 1684.400 1795.770 1684.460 ;
        RECT 1800.050 1684.400 1800.370 1684.460 ;
        RECT 1800.050 32.200 1800.370 32.260 ;
        RECT 2381.490 32.200 2381.810 32.260 ;
        RECT 1800.050 32.060 2381.810 32.200 ;
        RECT 1800.050 32.000 1800.370 32.060 ;
        RECT 2381.490 32.000 2381.810 32.060 ;
      LAYER via ;
        RECT 1795.480 1684.400 1795.740 1684.660 ;
        RECT 1800.080 1684.400 1800.340 1684.660 ;
        RECT 1800.080 32.000 1800.340 32.260 ;
        RECT 2381.520 32.000 2381.780 32.260 ;
      LAYER met2 ;
        RECT 1795.470 1700.000 1795.750 1704.000 ;
        RECT 1795.540 1684.690 1795.680 1700.000 ;
        RECT 1795.480 1684.370 1795.740 1684.690 ;
        RECT 1800.080 1684.370 1800.340 1684.690 ;
        RECT 1800.140 32.290 1800.280 1684.370 ;
        RECT 1800.080 31.970 1800.340 32.290 ;
        RECT 2381.520 31.970 2381.780 32.290 ;
        RECT 2381.580 2.400 2381.720 31.970 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 0.300 ;
=======
      LAYER met1 ;
        RECT 1799.590 31.860 1799.910 31.920 ;
        RECT 2399.430 31.860 2399.750 31.920 ;
        RECT 1799.590 31.720 2399.750 31.860 ;
        RECT 1799.590 31.660 1799.910 31.720 ;
        RECT 2399.430 31.660 2399.750 31.720 ;
      LAYER via ;
        RECT 1799.620 31.660 1799.880 31.920 ;
        RECT 2399.460 31.660 2399.720 31.920 ;
      LAYER met2 ;
        RECT 1800.070 1700.410 1800.350 1704.000 ;
        RECT 1799.680 1700.270 1800.350 1700.410 ;
        RECT 1799.680 31.950 1799.820 1700.270 ;
        RECT 1800.070 1700.000 1800.350 1700.270 ;
        RECT 1799.620 31.630 1799.880 31.950 ;
        RECT 2399.460 31.630 2399.720 31.950 ;
        RECT 2399.520 2.400 2399.660 31.630 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1800.070 33.520 1800.350 33.800 ;
        RECT 2399.450 33.520 2399.730 33.800 ;
      LAYER met3 ;
        RECT 1800.045 33.810 1800.375 33.825 ;
        RECT 2399.425 33.810 2399.755 33.825 ;
        RECT 1800.045 33.510 2399.755 33.810 ;
        RECT 1800.045 33.495 1800.375 33.510 ;
        RECT 2399.425 33.495 2399.755 33.510 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 0.300 ;
=======
      LAYER li1 ;
        RECT 1360.825 1545.725 1360.995 1593.835 ;
        RECT 1360.825 1400.885 1360.995 1448.995 ;
        RECT 1360.825 1207.425 1360.995 1255.875 ;
        RECT 1360.825 1062.585 1360.995 1110.695 ;
        RECT 1360.825 821.185 1360.995 910.775 ;
        RECT 1361.285 517.565 1361.455 565.675 ;
      LAYER mcon ;
        RECT 1360.825 1593.665 1360.995 1593.835 ;
        RECT 1360.825 1448.825 1360.995 1448.995 ;
        RECT 1360.825 1255.705 1360.995 1255.875 ;
        RECT 1360.825 1110.525 1360.995 1110.695 ;
        RECT 1360.825 910.605 1360.995 910.775 ;
        RECT 1361.285 565.505 1361.455 565.675 ;
      LAYER met1 ;
        RECT 1360.750 1593.820 1361.070 1593.880 ;
        RECT 1360.555 1593.680 1361.070 1593.820 ;
        RECT 1360.750 1593.620 1361.070 1593.680 ;
        RECT 1360.765 1545.880 1361.055 1545.925 ;
        RECT 1361.210 1545.880 1361.530 1545.940 ;
        RECT 1360.765 1545.740 1361.530 1545.880 ;
        RECT 1360.765 1545.695 1361.055 1545.740 ;
        RECT 1361.210 1545.680 1361.530 1545.740 ;
        RECT 1360.765 1448.980 1361.055 1449.025 ;
        RECT 1361.210 1448.980 1361.530 1449.040 ;
        RECT 1360.765 1448.840 1361.530 1448.980 ;
        RECT 1360.765 1448.795 1361.055 1448.840 ;
        RECT 1361.210 1448.780 1361.530 1448.840 ;
        RECT 1360.750 1401.040 1361.070 1401.100 ;
        RECT 1360.555 1400.900 1361.070 1401.040 ;
        RECT 1360.750 1400.840 1361.070 1400.900 ;
        RECT 1361.210 1304.820 1361.530 1304.880 ;
        RECT 1360.840 1304.680 1361.530 1304.820 ;
        RECT 1360.840 1304.540 1360.980 1304.680 ;
        RECT 1361.210 1304.620 1361.530 1304.680 ;
        RECT 1360.750 1304.280 1361.070 1304.540 ;
        RECT 1360.750 1255.860 1361.070 1255.920 ;
        RECT 1360.555 1255.720 1361.070 1255.860 ;
        RECT 1360.750 1255.660 1361.070 1255.720 ;
        RECT 1360.750 1207.580 1361.070 1207.640 ;
        RECT 1360.555 1207.440 1361.070 1207.580 ;
        RECT 1360.750 1207.380 1361.070 1207.440 ;
        RECT 1360.750 1110.680 1361.070 1110.740 ;
        RECT 1360.555 1110.540 1361.070 1110.680 ;
        RECT 1360.750 1110.480 1361.070 1110.540 ;
        RECT 1360.765 1062.740 1361.055 1062.785 ;
        RECT 1361.210 1062.740 1361.530 1062.800 ;
        RECT 1360.765 1062.600 1361.530 1062.740 ;
        RECT 1360.765 1062.555 1361.055 1062.600 ;
        RECT 1361.210 1062.540 1361.530 1062.600 ;
        RECT 1360.750 918.240 1361.070 918.300 ;
        RECT 1361.210 918.240 1361.530 918.300 ;
        RECT 1360.750 918.100 1361.530 918.240 ;
        RECT 1360.750 918.040 1361.070 918.100 ;
        RECT 1361.210 918.040 1361.530 918.100 ;
        RECT 1360.750 910.760 1361.070 910.820 ;
        RECT 1360.555 910.620 1361.070 910.760 ;
        RECT 1360.750 910.560 1361.070 910.620 ;
        RECT 1360.750 821.340 1361.070 821.400 ;
        RECT 1360.555 821.200 1361.070 821.340 ;
        RECT 1360.750 821.140 1361.070 821.200 ;
        RECT 1358.910 814.200 1359.230 814.260 ;
        RECT 1360.750 814.200 1361.070 814.260 ;
        RECT 1358.910 814.060 1361.070 814.200 ;
        RECT 1358.910 814.000 1359.230 814.060 ;
        RECT 1360.750 814.000 1361.070 814.060 ;
        RECT 1360.750 765.920 1361.070 765.980 ;
        RECT 1361.670 765.920 1361.990 765.980 ;
        RECT 1360.750 765.780 1361.990 765.920 ;
        RECT 1360.750 765.720 1361.070 765.780 ;
        RECT 1361.670 765.720 1361.990 765.780 ;
        RECT 1358.910 717.640 1359.230 717.700 ;
        RECT 1360.750 717.640 1361.070 717.700 ;
        RECT 1358.910 717.500 1361.070 717.640 ;
        RECT 1358.910 717.440 1359.230 717.500 ;
        RECT 1360.750 717.440 1361.070 717.500 ;
        RECT 1361.225 565.660 1361.515 565.705 ;
        RECT 1361.670 565.660 1361.990 565.720 ;
        RECT 1361.225 565.520 1361.990 565.660 ;
        RECT 1361.225 565.475 1361.515 565.520 ;
        RECT 1361.670 565.460 1361.990 565.520 ;
        RECT 1361.210 517.720 1361.530 517.780 ;
        RECT 1361.015 517.580 1361.530 517.720 ;
        RECT 1361.210 517.520 1361.530 517.580 ;
        RECT 1360.750 427.960 1361.070 428.020 ;
        RECT 1361.210 427.960 1361.530 428.020 ;
        RECT 1360.750 427.820 1361.530 427.960 ;
        RECT 1360.750 427.760 1361.070 427.820 ;
        RECT 1361.210 427.760 1361.530 427.820 ;
        RECT 1360.750 283.120 1361.070 283.180 ;
        RECT 1361.210 283.120 1361.530 283.180 ;
        RECT 1360.750 282.980 1361.530 283.120 ;
        RECT 1360.750 282.920 1361.070 282.980 ;
        RECT 1361.210 282.920 1361.530 282.980 ;
        RECT 800.010 50.900 800.330 50.960 ;
        RECT 1361.210 50.900 1361.530 50.960 ;
        RECT 800.010 50.760 1361.530 50.900 ;
        RECT 800.010 50.700 800.330 50.760 ;
        RECT 1361.210 50.700 1361.530 50.760 ;
=======
      LAYER met1 ;
        RECT 1360.750 1678.140 1361.070 1678.200 ;
        RECT 1363.510 1678.140 1363.830 1678.200 ;
        RECT 1360.750 1678.000 1363.830 1678.140 ;
        RECT 1360.750 1677.940 1361.070 1678.000 ;
        RECT 1363.510 1677.940 1363.830 1678.000 ;
        RECT 800.010 1604.700 800.330 1604.760 ;
        RECT 1360.750 1604.700 1361.070 1604.760 ;
        RECT 800.010 1604.560 1361.070 1604.700 ;
        RECT 800.010 1604.500 800.330 1604.560 ;
        RECT 1360.750 1604.500 1361.070 1604.560 ;
>>>>>>> re-updated local openlane
        RECT 793.570 20.980 793.890 21.040 ;
        RECT 800.010 20.980 800.330 21.040 ;
        RECT 793.570 20.840 800.330 20.980 ;
        RECT 793.570 20.780 793.890 20.840 ;
        RECT 800.010 20.780 800.330 20.840 ;
      LAYER via ;
        RECT 1360.780 1677.940 1361.040 1678.200 ;
        RECT 1363.540 1677.940 1363.800 1678.200 ;
        RECT 800.040 1604.500 800.300 1604.760 ;
        RECT 1360.780 1604.500 1361.040 1604.760 ;
        RECT 793.600 20.780 793.860 21.040 ;
        RECT 800.040 20.780 800.300 21.040 ;
      LAYER met2 ;
        RECT 1364.910 1700.410 1365.190 1704.000 ;
        RECT 1363.600 1700.270 1365.190 1700.410 ;
        RECT 1363.600 1678.230 1363.740 1700.270 ;
        RECT 1364.910 1700.000 1365.190 1700.270 ;
        RECT 1360.780 1677.910 1361.040 1678.230 ;
        RECT 1363.540 1677.910 1363.800 1678.230 ;
        RECT 1360.840 1604.790 1360.980 1677.910 ;
        RECT 800.040 1604.470 800.300 1604.790 ;
        RECT 1360.780 1604.470 1361.040 1604.790 ;
        RECT 800.100 21.070 800.240 1604.470 ;
        RECT 793.600 20.750 793.860 21.070 ;
        RECT 800.040 20.750 800.300 21.070 ;
        RECT 793.660 2.400 793.800 20.750 ;
        RECT 793.450 -4.800 794.010 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1358.930 765.880 1359.210 766.160 ;
        RECT 1360.770 765.880 1361.050 766.160 ;
        RECT 1360.770 717.600 1361.050 717.880 ;
        RECT 1361.690 717.600 1361.970 717.880 ;
        RECT 1358.930 669.320 1359.210 669.600 ;
        RECT 1360.770 669.320 1361.050 669.600 ;
        RECT 1360.770 470.080 1361.050 470.360 ;
        RECT 1361.230 469.400 1361.510 469.680 ;
        RECT 1360.770 144.360 1361.050 144.640 ;
        RECT 1361.230 143.680 1361.510 143.960 ;
      LAYER met3 ;
        RECT 1358.905 766.170 1359.235 766.185 ;
        RECT 1360.745 766.170 1361.075 766.185 ;
        RECT 1358.905 765.870 1361.075 766.170 ;
        RECT 1358.905 765.855 1359.235 765.870 ;
        RECT 1360.745 765.855 1361.075 765.870 ;
        RECT 1360.745 717.890 1361.075 717.905 ;
        RECT 1361.665 717.890 1361.995 717.905 ;
        RECT 1360.745 717.590 1361.995 717.890 ;
        RECT 1360.745 717.575 1361.075 717.590 ;
        RECT 1361.665 717.575 1361.995 717.590 ;
        RECT 1358.905 669.610 1359.235 669.625 ;
        RECT 1360.745 669.610 1361.075 669.625 ;
        RECT 1358.905 669.310 1361.075 669.610 ;
        RECT 1358.905 669.295 1359.235 669.310 ;
        RECT 1360.745 669.295 1361.075 669.310 ;
        RECT 1360.745 470.370 1361.075 470.385 ;
        RECT 1360.745 470.070 1362.210 470.370 ;
        RECT 1360.745 470.055 1361.075 470.070 ;
        RECT 1361.205 469.690 1361.535 469.705 ;
        RECT 1361.910 469.690 1362.210 470.070 ;
        RECT 1361.205 469.390 1362.210 469.690 ;
        RECT 1361.205 469.375 1361.535 469.390 ;
        RECT 1360.745 144.650 1361.075 144.665 ;
        RECT 1360.070 144.350 1361.075 144.650 ;
        RECT 1360.070 143.970 1360.370 144.350 ;
        RECT 1360.745 144.335 1361.075 144.350 ;
        RECT 1361.205 143.970 1361.535 143.985 ;
        RECT 1360.070 143.670 1361.535 143.970 ;
        RECT 1361.205 143.655 1361.535 143.670 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1293.590 1688.340 1293.910 1688.400 ;
        RECT 1323.030 1688.340 1323.350 1688.400 ;
        RECT 1293.590 1688.200 1323.350 1688.340 ;
        RECT 1293.590 1688.140 1293.910 1688.200 ;
        RECT 1323.030 1688.140 1323.350 1688.200 ;
        RECT 641.310 1611.160 641.630 1611.220 ;
        RECT 1293.590 1611.160 1293.910 1611.220 ;
        RECT 641.310 1611.020 1293.910 1611.160 ;
        RECT 641.310 1610.960 641.630 1611.020 ;
        RECT 1293.590 1610.960 1293.910 1611.020 ;
      LAYER via ;
        RECT 1293.620 1688.140 1293.880 1688.400 ;
        RECT 1323.060 1688.140 1323.320 1688.400 ;
        RECT 641.340 1610.960 641.600 1611.220 ;
        RECT 1293.620 1610.960 1293.880 1611.220 ;
      LAYER met2 ;
        RECT 1323.050 1700.000 1323.330 1704.000 ;
        RECT 1323.120 1688.430 1323.260 1700.000 ;
        RECT 1293.620 1688.110 1293.880 1688.430 ;
        RECT 1323.060 1688.110 1323.320 1688.430 ;
        RECT 1293.680 1611.250 1293.820 1688.110 ;
        RECT 641.340 1610.930 641.600 1611.250 ;
        RECT 1293.620 1610.930 1293.880 1611.250 ;
        RECT 641.400 17.410 641.540 1610.930 ;
        RECT 639.100 17.270 641.540 17.410 ;
        RECT 639.100 2.400 639.240 17.270 ;
        RECT 638.890 -4.800 639.450 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 639.030 32.840 639.310 33.120 ;
        RECT 1318.450 32.840 1318.730 33.120 ;
      LAYER met3 ;
        RECT 639.005 33.130 639.335 33.145 ;
        RECT 1318.425 33.130 1318.755 33.145 ;
        RECT 639.005 32.830 1318.755 33.130 ;
        RECT 639.005 32.815 639.335 32.830 ;
        RECT 1318.425 32.815 1318.755 32.830 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1806.950 31.520 1807.270 31.580 ;
        RECT 2422.890 31.520 2423.210 31.580 ;
        RECT 1806.950 31.380 2423.210 31.520 ;
        RECT 1806.950 31.320 1807.270 31.380 ;
        RECT 2422.890 31.320 2423.210 31.380 ;
      LAYER via ;
        RECT 1806.980 31.320 1807.240 31.580 ;
        RECT 2422.920 31.320 2423.180 31.580 ;
      LAYER met2 ;
        RECT 1806.510 1700.410 1806.790 1704.000 ;
        RECT 1806.510 1700.270 1807.180 1700.410 ;
        RECT 1806.510 1700.000 1806.790 1700.270 ;
        RECT 1807.040 31.610 1807.180 1700.270 ;
        RECT 1806.980 31.290 1807.240 31.610 ;
        RECT 2422.920 31.290 2423.180 31.610 ;
        RECT 2422.980 2.400 2423.120 31.290 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1807.430 32.840 1807.710 33.120 ;
        RECT 2422.910 32.840 2423.190 33.120 ;
      LAYER met3 ;
        RECT 1807.405 33.130 1807.735 33.145 ;
        RECT 2422.885 33.130 2423.215 33.145 ;
        RECT 1807.405 32.830 2423.215 33.130 ;
        RECT 1807.405 32.815 1807.735 32.830 ;
        RECT 2422.885 32.815 2423.215 32.830 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1811.550 1683.920 1811.870 1683.980 ;
        RECT 1814.310 1683.920 1814.630 1683.980 ;
        RECT 1811.550 1683.780 1814.630 1683.920 ;
        RECT 1811.550 1683.720 1811.870 1683.780 ;
        RECT 1814.310 1683.720 1814.630 1683.780 ;
        RECT 1814.310 31.180 1814.630 31.240 ;
        RECT 2440.830 31.180 2441.150 31.240 ;
        RECT 1814.310 31.040 2441.150 31.180 ;
        RECT 1814.310 30.980 1814.630 31.040 ;
        RECT 2440.830 30.980 2441.150 31.040 ;
      LAYER via ;
        RECT 1811.580 1683.720 1811.840 1683.980 ;
        RECT 1814.340 1683.720 1814.600 1683.980 ;
        RECT 1814.340 30.980 1814.600 31.240 ;
        RECT 2440.860 30.980 2441.120 31.240 ;
      LAYER met2 ;
        RECT 1811.570 1700.000 1811.850 1704.000 ;
        RECT 1811.640 1684.010 1811.780 1700.000 ;
        RECT 1811.580 1683.690 1811.840 1684.010 ;
        RECT 1814.340 1683.690 1814.600 1684.010 ;
        RECT 1814.400 31.270 1814.540 1683.690 ;
        RECT 1814.340 30.950 1814.600 31.270 ;
        RECT 2440.860 30.950 2441.120 31.270 ;
        RECT 2440.920 2.400 2441.060 30.950 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1814.330 32.160 1814.610 32.440 ;
        RECT 2440.850 32.160 2441.130 32.440 ;
      LAYER met3 ;
        RECT 1814.305 32.450 1814.635 32.465 ;
        RECT 2440.825 32.450 2441.155 32.465 ;
        RECT 1814.305 32.150 2441.155 32.450 ;
        RECT 1814.305 32.135 1814.635 32.150 ;
        RECT 2440.825 32.135 2441.155 32.150 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2458.650 -4.800 2459.210 0.300 ;
=======
        RECT 1813.870 1700.000 1814.150 1704.000 ;
        RECT 1813.940 31.805 1814.080 1700.000 ;
        RECT 1813.870 31.435 1814.150 31.805 ;
        RECT 2458.790 31.435 2459.070 31.805 ;
        RECT 2458.860 2.400 2459.000 31.435 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
      LAYER via2 ;
        RECT 1813.870 31.480 1814.150 31.760 ;
        RECT 2458.790 31.480 2459.070 31.760 ;
      LAYER met3 ;
        RECT 1813.845 31.770 1814.175 31.785 ;
        RECT 2458.765 31.770 2459.095 31.785 ;
        RECT 1813.845 31.470 2459.095 31.770 ;
        RECT 1813.845 31.455 1814.175 31.470 ;
        RECT 2458.765 31.455 2459.095 31.470 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1816.150 1683.920 1816.470 1683.980 ;
        RECT 1818.910 1683.920 1819.230 1683.980 ;
        RECT 1816.150 1683.780 1819.230 1683.920 ;
        RECT 1816.150 1683.720 1816.470 1683.780 ;
        RECT 1818.910 1683.720 1819.230 1683.780 ;
        RECT 1819.370 30.840 1819.690 30.900 ;
        RECT 2458.770 30.840 2459.090 30.900 ;
        RECT 1819.370 30.700 2459.090 30.840 ;
        RECT 1819.370 30.640 1819.690 30.700 ;
        RECT 2458.770 30.640 2459.090 30.700 ;
      LAYER via ;
        RECT 1816.180 1683.720 1816.440 1683.980 ;
        RECT 1818.940 1683.720 1819.200 1683.980 ;
        RECT 1819.400 30.640 1819.660 30.900 ;
        RECT 2458.800 30.640 2459.060 30.900 ;
      LAYER met2 ;
        RECT 1816.170 1700.000 1816.450 1704.000 ;
        RECT 1816.240 1684.010 1816.380 1700.000 ;
        RECT 1816.180 1683.690 1816.440 1684.010 ;
        RECT 1818.940 1683.690 1819.200 1684.010 ;
        RECT 1819.000 1656.210 1819.140 1683.690 ;
        RECT 1819.000 1656.070 1819.600 1656.210 ;
        RECT 1819.460 30.930 1819.600 1656.070 ;
        RECT 1819.400 30.610 1819.660 30.930 ;
        RECT 2458.800 30.610 2459.060 30.930 ;
        RECT 2458.860 2.400 2459.000 30.610 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2476.590 -4.800 2477.150 0.300 ;
=======
        RECT 1818.470 1700.410 1818.750 1704.000 ;
        RECT 1818.470 1700.270 1820.060 1700.410 ;
        RECT 1818.470 1700.000 1818.750 1700.270 ;
        RECT 1819.920 1670.490 1820.060 1700.270 ;
        RECT 1819.920 1670.350 1820.520 1670.490 ;
        RECT 1820.380 31.125 1820.520 1670.350 ;
        RECT 1820.310 30.755 1820.590 31.125 ;
        RECT 2476.730 30.755 2477.010 31.125 ;
        RECT 2476.800 2.400 2476.940 30.755 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
      LAYER via2 ;
        RECT 1820.310 30.800 1820.590 31.080 ;
        RECT 2476.730 30.800 2477.010 31.080 ;
      LAYER met3 ;
        RECT 1820.285 31.090 1820.615 31.105 ;
        RECT 2476.705 31.090 2477.035 31.105 ;
        RECT 1820.285 30.790 2477.035 31.090 ;
        RECT 1820.285 30.775 1820.615 30.790 ;
        RECT 2476.705 30.775 2477.035 30.790 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1820.290 72.320 1820.610 72.380 ;
        RECT 2470.270 72.320 2470.590 72.380 ;
        RECT 1820.290 72.180 2470.590 72.320 ;
        RECT 1820.290 72.120 1820.610 72.180 ;
        RECT 2470.270 72.120 2470.590 72.180 ;
        RECT 2470.270 35.940 2470.590 36.000 ;
        RECT 2476.710 35.940 2477.030 36.000 ;
        RECT 2470.270 35.800 2477.030 35.940 ;
        RECT 2470.270 35.740 2470.590 35.800 ;
        RECT 2476.710 35.740 2477.030 35.800 ;
      LAYER via ;
        RECT 1820.320 72.120 1820.580 72.380 ;
        RECT 2470.300 72.120 2470.560 72.380 ;
        RECT 2470.300 35.740 2470.560 36.000 ;
        RECT 2476.740 35.740 2477.000 36.000 ;
      LAYER met2 ;
        RECT 1821.230 1700.410 1821.510 1704.000 ;
        RECT 1820.380 1700.270 1821.510 1700.410 ;
        RECT 1820.380 72.410 1820.520 1700.270 ;
        RECT 1821.230 1700.000 1821.510 1700.270 ;
        RECT 1820.320 72.090 1820.580 72.410 ;
        RECT 2470.300 72.090 2470.560 72.410 ;
        RECT 2470.360 36.030 2470.500 72.090 ;
        RECT 2470.300 35.710 2470.560 36.030 ;
        RECT 2476.740 35.710 2477.000 36.030 ;
        RECT 2476.800 2.400 2476.940 35.710 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1826.270 1673.040 1826.590 1673.100 ;
        RECT 2490.970 1673.040 2491.290 1673.100 ;
        RECT 1826.270 1672.900 2491.290 1673.040 ;
        RECT 1826.270 1672.840 1826.590 1672.900 ;
        RECT 2490.970 1672.840 2491.290 1672.900 ;
      LAYER via ;
        RECT 1826.300 1672.840 1826.560 1673.100 ;
        RECT 2491.000 1672.840 2491.260 1673.100 ;
      LAYER met2 ;
        RECT 1826.290 1700.000 1826.570 1704.000 ;
        RECT 1826.360 1673.130 1826.500 1700.000 ;
        RECT 1826.300 1672.810 1826.560 1673.130 ;
        RECT 2491.000 1672.810 2491.260 1673.130 ;
        RECT 2491.060 16.730 2491.200 1672.810 ;
        RECT 2491.060 16.590 2494.880 16.730 ;
        RECT 2494.740 2.400 2494.880 16.590 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1826.290 46.440 1826.570 46.720 ;
        RECT 2494.670 46.440 2494.950 46.720 ;
      LAYER met3 ;
        RECT 1826.265 46.730 1826.595 46.745 ;
        RECT 2494.645 46.730 2494.975 46.745 ;
        RECT 1826.265 46.430 2494.975 46.730 ;
        RECT 1826.265 46.415 1826.595 46.430 ;
        RECT 2494.645 46.415 2494.975 46.430 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1830.870 1684.940 1831.190 1685.000 ;
        RECT 1834.550 1684.940 1834.870 1685.000 ;
        RECT 1830.870 1684.800 1834.870 1684.940 ;
        RECT 1830.870 1684.740 1831.190 1684.800 ;
        RECT 1834.550 1684.740 1834.870 1684.800 ;
        RECT 1834.550 879.820 1834.870 879.880 ;
        RECT 2511.670 879.820 2511.990 879.880 ;
        RECT 1834.550 879.680 2511.990 879.820 ;
        RECT 1834.550 879.620 1834.870 879.680 ;
        RECT 2511.670 879.620 2511.990 879.680 ;
      LAYER via ;
        RECT 1830.900 1684.740 1831.160 1685.000 ;
        RECT 1834.580 1684.740 1834.840 1685.000 ;
        RECT 1834.580 879.620 1834.840 879.880 ;
        RECT 2511.700 879.620 2511.960 879.880 ;
      LAYER met2 ;
        RECT 1830.890 1700.000 1831.170 1704.000 ;
        RECT 1830.960 1685.030 1831.100 1700.000 ;
        RECT 1830.900 1684.710 1831.160 1685.030 ;
        RECT 1834.580 1684.710 1834.840 1685.030 ;
        RECT 1834.640 879.910 1834.780 1684.710 ;
        RECT 1834.580 879.590 1834.840 879.910 ;
        RECT 2511.700 879.590 2511.960 879.910 ;
        RECT 2511.760 17.410 2511.900 879.590 ;
        RECT 2511.760 17.270 2512.360 17.410 ;
        RECT 2512.220 2.400 2512.360 17.270 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1826.750 45.760 1827.030 46.040 ;
        RECT 2512.150 45.760 2512.430 46.040 ;
      LAYER met3 ;
        RECT 1826.725 46.050 1827.055 46.065 ;
        RECT 2512.125 46.050 2512.455 46.065 ;
        RECT 1826.725 45.750 2512.455 46.050 ;
        RECT 1826.725 45.735 1827.055 45.750 ;
        RECT 2512.125 45.735 2512.455 45.750 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 0.300 ;
=======
      LAYER met1 ;
        RECT 1835.930 1684.940 1836.250 1685.000 ;
        RECT 1841.450 1684.940 1841.770 1685.000 ;
        RECT 1835.930 1684.800 1841.770 1684.940 ;
        RECT 1835.930 1684.740 1836.250 1684.800 ;
        RECT 1841.450 1684.740 1841.770 1684.800 ;
        RECT 1841.450 1590.420 1841.770 1590.480 ;
        RECT 2525.470 1590.420 2525.790 1590.480 ;
        RECT 1841.450 1590.280 2525.790 1590.420 ;
        RECT 1841.450 1590.220 1841.770 1590.280 ;
        RECT 2525.470 1590.220 2525.790 1590.280 ;
        RECT 2525.470 62.120 2525.790 62.180 ;
        RECT 2530.070 62.120 2530.390 62.180 ;
        RECT 2525.470 61.980 2530.390 62.120 ;
        RECT 2525.470 61.920 2525.790 61.980 ;
        RECT 2530.070 61.920 2530.390 61.980 ;
      LAYER via ;
        RECT 1835.960 1684.740 1836.220 1685.000 ;
        RECT 1841.480 1684.740 1841.740 1685.000 ;
        RECT 1841.480 1590.220 1841.740 1590.480 ;
        RECT 2525.500 1590.220 2525.760 1590.480 ;
        RECT 2525.500 61.920 2525.760 62.180 ;
        RECT 2530.100 61.920 2530.360 62.180 ;
      LAYER met2 ;
        RECT 1835.950 1700.000 1836.230 1704.000 ;
        RECT 1836.020 1685.030 1836.160 1700.000 ;
        RECT 1835.960 1684.710 1836.220 1685.030 ;
        RECT 1841.480 1684.710 1841.740 1685.030 ;
        RECT 1841.540 1590.510 1841.680 1684.710 ;
        RECT 1841.480 1590.190 1841.740 1590.510 ;
        RECT 2525.500 1590.190 2525.760 1590.510 ;
        RECT 2525.560 62.210 2525.700 1590.190 ;
        RECT 2525.500 61.890 2525.760 62.210 ;
        RECT 2530.100 61.890 2530.360 62.210 ;
        RECT 2530.160 2.400 2530.300 61.890 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1832.730 45.080 1833.010 45.360 ;
        RECT 2530.090 45.080 2530.370 45.360 ;
      LAYER met3 ;
        RECT 1832.705 45.370 1833.035 45.385 ;
        RECT 2530.065 45.370 2530.395 45.385 ;
        RECT 1832.705 45.070 2530.395 45.370 ;
        RECT 1832.705 45.055 1833.035 45.070 ;
        RECT 2530.065 45.055 2530.395 45.070 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1837.770 1684.600 1838.090 1684.660 ;
        RECT 1840.990 1684.600 1841.310 1684.660 ;
        RECT 1837.770 1684.460 1841.310 1684.600 ;
        RECT 1837.770 1684.400 1838.090 1684.460 ;
        RECT 1840.990 1684.400 1841.310 1684.460 ;
        RECT 1840.990 36.620 1841.310 36.680 ;
        RECT 2548.010 36.620 2548.330 36.680 ;
        RECT 1840.990 36.480 2548.330 36.620 ;
        RECT 1840.990 36.420 1841.310 36.480 ;
        RECT 2548.010 36.420 2548.330 36.480 ;
      LAYER via ;
        RECT 1837.800 1684.400 1838.060 1684.660 ;
        RECT 1841.020 1684.400 1841.280 1684.660 ;
        RECT 1841.020 36.420 1841.280 36.680 ;
        RECT 2548.040 36.420 2548.300 36.680 ;
      LAYER met2 ;
        RECT 1837.790 1700.000 1838.070 1704.000 ;
        RECT 1837.860 1684.690 1838.000 1700.000 ;
        RECT 1837.800 1684.370 1838.060 1684.690 ;
        RECT 1841.020 1684.370 1841.280 1684.690 ;
        RECT 1841.080 36.710 1841.220 1684.370 ;
        RECT 1841.020 36.390 1841.280 36.710 ;
        RECT 2548.040 36.390 2548.300 36.710 ;
        RECT 2548.100 2.400 2548.240 36.390 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 2546.245 1538.925 2546.415 1587.035 ;
        RECT 2546.245 1442.025 2546.415 1490.475 ;
        RECT 2546.245 766.105 2546.415 814.215 ;
        RECT 2546.245 669.545 2546.415 717.655 ;
        RECT 2546.245 572.645 2546.415 620.755 ;
        RECT 2546.245 476.085 2546.415 524.195 ;
        RECT 2546.245 282.965 2546.415 331.075 ;
        RECT 2546.245 186.405 2546.415 234.515 ;
        RECT 2546.245 89.845 2546.415 137.955 ;
      LAYER mcon ;
        RECT 2546.245 1586.865 2546.415 1587.035 ;
        RECT 2546.245 1490.305 2546.415 1490.475 ;
        RECT 2546.245 814.045 2546.415 814.215 ;
        RECT 2546.245 717.485 2546.415 717.655 ;
        RECT 2546.245 620.585 2546.415 620.755 ;
        RECT 2546.245 524.025 2546.415 524.195 ;
        RECT 2546.245 330.905 2546.415 331.075 ;
        RECT 2546.245 234.345 2546.415 234.515 ;
        RECT 2546.245 137.785 2546.415 137.955 ;
      LAYER met1 ;
        RECT 1840.990 1597.220 1841.310 1597.280 ;
        RECT 2546.170 1597.220 2546.490 1597.280 ;
        RECT 1840.990 1597.080 2546.490 1597.220 ;
        RECT 1840.990 1597.020 1841.310 1597.080 ;
        RECT 2546.170 1597.020 2546.490 1597.080 ;
        RECT 2546.170 1587.020 2546.490 1587.080 ;
        RECT 2545.975 1586.880 2546.490 1587.020 ;
        RECT 2546.170 1586.820 2546.490 1586.880 ;
        RECT 2546.170 1539.080 2546.490 1539.140 ;
        RECT 2545.975 1538.940 2546.490 1539.080 ;
        RECT 2546.170 1538.880 2546.490 1538.940 ;
        RECT 2546.170 1490.460 2546.490 1490.520 ;
        RECT 2545.975 1490.320 2546.490 1490.460 ;
        RECT 2546.170 1490.260 2546.490 1490.320 ;
        RECT 2546.170 1442.180 2546.490 1442.240 ;
        RECT 2545.975 1442.040 2546.490 1442.180 ;
        RECT 2546.170 1441.980 2546.490 1442.040 ;
        RECT 2545.250 1345.620 2545.570 1345.680 ;
        RECT 2546.170 1345.620 2546.490 1345.680 ;
        RECT 2545.250 1345.480 2546.490 1345.620 ;
        RECT 2545.250 1345.420 2545.570 1345.480 ;
        RECT 2546.170 1345.420 2546.490 1345.480 ;
        RECT 2545.250 1249.060 2545.570 1249.120 ;
        RECT 2546.170 1249.060 2546.490 1249.120 ;
        RECT 2545.250 1248.920 2546.490 1249.060 ;
        RECT 2545.250 1248.860 2545.570 1248.920 ;
        RECT 2546.170 1248.860 2546.490 1248.920 ;
        RECT 2545.250 1152.500 2545.570 1152.560 ;
        RECT 2546.170 1152.500 2546.490 1152.560 ;
        RECT 2545.250 1152.360 2546.490 1152.500 ;
        RECT 2545.250 1152.300 2545.570 1152.360 ;
        RECT 2546.170 1152.300 2546.490 1152.360 ;
        RECT 2545.250 1007.320 2545.570 1007.380 ;
        RECT 2546.170 1007.320 2546.490 1007.380 ;
        RECT 2545.250 1007.180 2546.490 1007.320 ;
        RECT 2545.250 1007.120 2545.570 1007.180 ;
        RECT 2546.170 1007.120 2546.490 1007.180 ;
        RECT 2545.250 910.760 2545.570 910.820 ;
        RECT 2546.170 910.760 2546.490 910.820 ;
        RECT 2545.250 910.620 2546.490 910.760 ;
        RECT 2545.250 910.560 2545.570 910.620 ;
        RECT 2546.170 910.560 2546.490 910.620 ;
        RECT 2546.170 814.200 2546.490 814.260 ;
        RECT 2545.975 814.060 2546.490 814.200 ;
        RECT 2546.170 814.000 2546.490 814.060 ;
        RECT 2546.170 766.260 2546.490 766.320 ;
        RECT 2545.975 766.120 2546.490 766.260 ;
        RECT 2546.170 766.060 2546.490 766.120 ;
        RECT 2546.170 717.640 2546.490 717.700 ;
        RECT 2545.975 717.500 2546.490 717.640 ;
        RECT 2546.170 717.440 2546.490 717.500 ;
        RECT 2546.170 669.700 2546.490 669.760 ;
        RECT 2545.975 669.560 2546.490 669.700 ;
        RECT 2546.170 669.500 2546.490 669.560 ;
        RECT 2546.170 620.740 2546.490 620.800 ;
        RECT 2545.975 620.600 2546.490 620.740 ;
        RECT 2546.170 620.540 2546.490 620.600 ;
        RECT 2546.170 572.800 2546.490 572.860 ;
        RECT 2545.975 572.660 2546.490 572.800 ;
        RECT 2546.170 572.600 2546.490 572.660 ;
        RECT 2546.170 524.180 2546.490 524.240 ;
        RECT 2545.975 524.040 2546.490 524.180 ;
        RECT 2546.170 523.980 2546.490 524.040 ;
        RECT 2546.170 476.240 2546.490 476.300 ;
        RECT 2545.975 476.100 2546.490 476.240 ;
        RECT 2546.170 476.040 2546.490 476.100 ;
        RECT 2546.170 331.060 2546.490 331.120 ;
        RECT 2545.975 330.920 2546.490 331.060 ;
        RECT 2546.170 330.860 2546.490 330.920 ;
        RECT 2546.170 283.120 2546.490 283.180 ;
        RECT 2545.975 282.980 2546.490 283.120 ;
        RECT 2546.170 282.920 2546.490 282.980 ;
        RECT 2546.170 234.500 2546.490 234.560 ;
        RECT 2545.975 234.360 2546.490 234.500 ;
        RECT 2546.170 234.300 2546.490 234.360 ;
        RECT 2546.170 186.560 2546.490 186.620 ;
        RECT 2545.975 186.420 2546.490 186.560 ;
        RECT 2546.170 186.360 2546.490 186.420 ;
        RECT 2546.170 137.940 2546.490 138.000 ;
        RECT 2545.975 137.800 2546.490 137.940 ;
        RECT 2546.170 137.740 2546.490 137.800 ;
        RECT 2546.170 90.000 2546.490 90.060 ;
        RECT 2545.975 89.860 2546.490 90.000 ;
        RECT 2546.170 89.800 2546.490 89.860 ;
      LAYER via ;
        RECT 1841.020 1597.020 1841.280 1597.280 ;
        RECT 2546.200 1597.020 2546.460 1597.280 ;
        RECT 2546.200 1586.820 2546.460 1587.080 ;
        RECT 2546.200 1538.880 2546.460 1539.140 ;
        RECT 2546.200 1490.260 2546.460 1490.520 ;
        RECT 2546.200 1441.980 2546.460 1442.240 ;
        RECT 2545.280 1345.420 2545.540 1345.680 ;
        RECT 2546.200 1345.420 2546.460 1345.680 ;
        RECT 2545.280 1248.860 2545.540 1249.120 ;
        RECT 2546.200 1248.860 2546.460 1249.120 ;
        RECT 2545.280 1152.300 2545.540 1152.560 ;
        RECT 2546.200 1152.300 2546.460 1152.560 ;
        RECT 2545.280 1007.120 2545.540 1007.380 ;
        RECT 2546.200 1007.120 2546.460 1007.380 ;
        RECT 2545.280 910.560 2545.540 910.820 ;
        RECT 2546.200 910.560 2546.460 910.820 ;
        RECT 2546.200 814.000 2546.460 814.260 ;
        RECT 2546.200 766.060 2546.460 766.320 ;
        RECT 2546.200 717.440 2546.460 717.700 ;
        RECT 2546.200 669.500 2546.460 669.760 ;
        RECT 2546.200 620.540 2546.460 620.800 ;
        RECT 2546.200 572.600 2546.460 572.860 ;
        RECT 2546.200 523.980 2546.460 524.240 ;
        RECT 2546.200 476.040 2546.460 476.300 ;
        RECT 2546.200 330.860 2546.460 331.120 ;
        RECT 2546.200 282.920 2546.460 283.180 ;
        RECT 2546.200 234.300 2546.460 234.560 ;
        RECT 2546.200 186.360 2546.460 186.620 ;
        RECT 2546.200 137.740 2546.460 138.000 ;
        RECT 2546.200 89.800 2546.460 90.060 ;
      LAYER met2 ;
        RECT 1840.550 1700.410 1840.830 1704.000 ;
        RECT 1840.550 1700.270 1841.220 1700.410 ;
        RECT 1840.550 1700.000 1840.830 1700.270 ;
        RECT 1841.080 1597.310 1841.220 1700.270 ;
        RECT 1841.020 1596.990 1841.280 1597.310 ;
        RECT 2546.200 1596.990 2546.460 1597.310 ;
        RECT 2546.260 1587.110 2546.400 1596.990 ;
        RECT 2546.200 1586.790 2546.460 1587.110 ;
        RECT 2546.200 1538.850 2546.460 1539.170 ;
        RECT 2546.260 1490.550 2546.400 1538.850 ;
        RECT 2546.200 1490.230 2546.460 1490.550 ;
        RECT 2546.200 1441.950 2546.460 1442.270 ;
        RECT 2546.260 1393.845 2546.400 1441.950 ;
        RECT 2545.270 1393.475 2545.550 1393.845 ;
        RECT 2546.190 1393.475 2546.470 1393.845 ;
        RECT 2545.340 1345.710 2545.480 1393.475 ;
        RECT 2545.280 1345.390 2545.540 1345.710 ;
        RECT 2546.200 1345.390 2546.460 1345.710 ;
        RECT 2546.260 1297.285 2546.400 1345.390 ;
        RECT 2545.270 1296.915 2545.550 1297.285 ;
        RECT 2546.190 1296.915 2546.470 1297.285 ;
        RECT 2545.340 1249.150 2545.480 1296.915 ;
        RECT 2545.280 1248.830 2545.540 1249.150 ;
        RECT 2546.200 1248.830 2546.460 1249.150 ;
        RECT 2546.260 1200.725 2546.400 1248.830 ;
        RECT 2545.270 1200.355 2545.550 1200.725 ;
        RECT 2546.190 1200.355 2546.470 1200.725 ;
        RECT 2545.340 1152.590 2545.480 1200.355 ;
        RECT 2545.280 1152.270 2545.540 1152.590 ;
        RECT 2546.200 1152.270 2546.460 1152.590 ;
        RECT 2546.260 1104.165 2546.400 1152.270 ;
        RECT 2545.270 1103.795 2545.550 1104.165 ;
        RECT 2546.190 1103.795 2546.470 1104.165 ;
        RECT 2545.340 1055.885 2545.480 1103.795 ;
        RECT 2545.270 1055.515 2545.550 1055.885 ;
        RECT 2546.190 1055.515 2546.470 1055.885 ;
        RECT 2546.260 1007.410 2546.400 1055.515 ;
        RECT 2545.280 1007.090 2545.540 1007.410 ;
        RECT 2546.200 1007.090 2546.460 1007.410 ;
        RECT 2545.340 959.325 2545.480 1007.090 ;
        RECT 2545.270 958.955 2545.550 959.325 ;
        RECT 2546.190 958.955 2546.470 959.325 ;
        RECT 2546.260 910.850 2546.400 958.955 ;
        RECT 2545.280 910.530 2545.540 910.850 ;
        RECT 2546.200 910.530 2546.460 910.850 ;
        RECT 2545.340 862.765 2545.480 910.530 ;
        RECT 2545.270 862.395 2545.550 862.765 ;
        RECT 2546.190 862.395 2546.470 862.765 ;
        RECT 2546.260 814.290 2546.400 862.395 ;
        RECT 2546.200 813.970 2546.460 814.290 ;
        RECT 2546.200 766.030 2546.460 766.350 ;
        RECT 2546.260 717.730 2546.400 766.030 ;
        RECT 2546.200 717.410 2546.460 717.730 ;
        RECT 2546.200 669.470 2546.460 669.790 ;
        RECT 2546.260 620.830 2546.400 669.470 ;
        RECT 2546.200 620.510 2546.460 620.830 ;
        RECT 2546.200 572.570 2546.460 572.890 ;
        RECT 2546.260 524.270 2546.400 572.570 ;
        RECT 2546.200 523.950 2546.460 524.270 ;
        RECT 2546.200 476.010 2546.460 476.330 ;
        RECT 2546.260 331.150 2546.400 476.010 ;
        RECT 2546.200 330.830 2546.460 331.150 ;
        RECT 2546.200 282.890 2546.460 283.210 ;
        RECT 2546.260 234.590 2546.400 282.890 ;
        RECT 2546.200 234.270 2546.460 234.590 ;
        RECT 2546.200 186.330 2546.460 186.650 ;
        RECT 2546.260 138.030 2546.400 186.330 ;
        RECT 2546.200 137.710 2546.460 138.030 ;
        RECT 2546.200 89.770 2546.460 90.090 ;
        RECT 2546.260 72.490 2546.400 89.770 ;
        RECT 2546.260 72.350 2546.860 72.490 ;
        RECT 2546.720 61.610 2546.860 72.350 ;
        RECT 2546.720 61.470 2548.240 61.610 ;
        RECT 2548.100 2.400 2548.240 61.470 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
      LAYER via2 ;
        RECT 2545.270 1393.520 2545.550 1393.800 ;
        RECT 2546.190 1393.520 2546.470 1393.800 ;
        RECT 2545.270 1296.960 2545.550 1297.240 ;
        RECT 2546.190 1296.960 2546.470 1297.240 ;
        RECT 2545.270 1200.400 2545.550 1200.680 ;
        RECT 2546.190 1200.400 2546.470 1200.680 ;
        RECT 2545.270 1103.840 2545.550 1104.120 ;
        RECT 2546.190 1103.840 2546.470 1104.120 ;
        RECT 2545.270 1055.560 2545.550 1055.840 ;
        RECT 2546.190 1055.560 2546.470 1055.840 ;
        RECT 2545.270 959.000 2545.550 959.280 ;
        RECT 2546.190 959.000 2546.470 959.280 ;
        RECT 2545.270 862.440 2545.550 862.720 ;
        RECT 2546.190 862.440 2546.470 862.720 ;
      LAYER met3 ;
        RECT 2545.245 1393.810 2545.575 1393.825 ;
        RECT 2546.165 1393.810 2546.495 1393.825 ;
        RECT 2545.245 1393.510 2546.495 1393.810 ;
        RECT 2545.245 1393.495 2545.575 1393.510 ;
        RECT 2546.165 1393.495 2546.495 1393.510 ;
        RECT 2545.245 1297.250 2545.575 1297.265 ;
        RECT 2546.165 1297.250 2546.495 1297.265 ;
        RECT 2545.245 1296.950 2546.495 1297.250 ;
        RECT 2545.245 1296.935 2545.575 1296.950 ;
        RECT 2546.165 1296.935 2546.495 1296.950 ;
        RECT 2545.245 1200.690 2545.575 1200.705 ;
        RECT 2546.165 1200.690 2546.495 1200.705 ;
        RECT 2545.245 1200.390 2546.495 1200.690 ;
        RECT 2545.245 1200.375 2545.575 1200.390 ;
        RECT 2546.165 1200.375 2546.495 1200.390 ;
        RECT 2545.245 1104.130 2545.575 1104.145 ;
        RECT 2546.165 1104.130 2546.495 1104.145 ;
        RECT 2545.245 1103.830 2546.495 1104.130 ;
        RECT 2545.245 1103.815 2545.575 1103.830 ;
        RECT 2546.165 1103.815 2546.495 1103.830 ;
        RECT 2545.245 1055.850 2545.575 1055.865 ;
        RECT 2546.165 1055.850 2546.495 1055.865 ;
        RECT 2545.245 1055.550 2546.495 1055.850 ;
        RECT 2545.245 1055.535 2545.575 1055.550 ;
        RECT 2546.165 1055.535 2546.495 1055.550 ;
        RECT 2545.245 959.290 2545.575 959.305 ;
        RECT 2546.165 959.290 2546.495 959.305 ;
        RECT 2545.245 958.990 2546.495 959.290 ;
        RECT 2545.245 958.975 2545.575 958.990 ;
        RECT 2546.165 958.975 2546.495 958.990 ;
        RECT 2545.245 862.730 2545.575 862.745 ;
        RECT 2546.165 862.730 2546.495 862.745 ;
        RECT 2545.245 862.430 2546.495 862.730 ;
        RECT 2545.245 862.415 2545.575 862.430 ;
        RECT 2546.165 862.415 2546.495 862.430 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1845.590 1684.940 1845.910 1685.000 ;
        RECT 1846.970 1684.940 1847.290 1685.000 ;
        RECT 1845.590 1684.800 1847.290 1684.940 ;
        RECT 1845.590 1684.740 1845.910 1684.800 ;
        RECT 1846.970 1684.740 1847.290 1684.800 ;
        RECT 1846.970 1583.620 1847.290 1583.680 ;
        RECT 2559.970 1583.620 2560.290 1583.680 ;
        RECT 1846.970 1583.480 2560.290 1583.620 ;
        RECT 1846.970 1583.420 1847.290 1583.480 ;
        RECT 2559.970 1583.420 2560.290 1583.480 ;
        RECT 2559.970 35.940 2560.290 36.000 ;
        RECT 2565.950 35.940 2566.270 36.000 ;
        RECT 2559.970 35.800 2566.270 35.940 ;
        RECT 2559.970 35.740 2560.290 35.800 ;
        RECT 2565.950 35.740 2566.270 35.800 ;
      LAYER via ;
        RECT 1845.620 1684.740 1845.880 1685.000 ;
        RECT 1847.000 1684.740 1847.260 1685.000 ;
        RECT 1847.000 1583.420 1847.260 1583.680 ;
        RECT 2560.000 1583.420 2560.260 1583.680 ;
        RECT 2560.000 35.740 2560.260 36.000 ;
        RECT 2565.980 35.740 2566.240 36.000 ;
      LAYER met2 ;
        RECT 1845.610 1700.000 1845.890 1704.000 ;
        RECT 1845.680 1685.030 1845.820 1700.000 ;
        RECT 1845.620 1684.710 1845.880 1685.030 ;
        RECT 1847.000 1684.710 1847.260 1685.030 ;
        RECT 1847.060 1583.710 1847.200 1684.710 ;
        RECT 1847.000 1583.390 1847.260 1583.710 ;
        RECT 2560.000 1583.390 2560.260 1583.710 ;
        RECT 2560.060 36.030 2560.200 1583.390 ;
        RECT 2560.000 35.710 2560.260 36.030 ;
        RECT 2565.980 35.710 2566.240 36.030 ;
        RECT 2566.040 2.400 2566.180 35.710 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1847.890 37.300 1848.210 37.360 ;
        RECT 2583.890 37.300 2584.210 37.360 ;
        RECT 1847.890 37.160 2584.210 37.300 ;
        RECT 1847.890 37.100 1848.210 37.160 ;
        RECT 2583.890 37.100 2584.210 37.160 ;
      LAYER via ;
        RECT 1847.920 37.100 1848.180 37.360 ;
        RECT 2583.920 37.100 2584.180 37.360 ;
      LAYER met2 ;
        RECT 1847.450 1700.410 1847.730 1704.000 ;
        RECT 1847.450 1700.270 1848.120 1700.410 ;
        RECT 1847.450 1700.000 1847.730 1700.270 ;
        RECT 1847.980 37.390 1848.120 1700.270 ;
        RECT 1847.920 37.070 1848.180 37.390 ;
        RECT 2583.920 37.070 2584.180 37.390 ;
        RECT 2583.980 2.400 2584.120 37.070 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 2580.745 1538.925 2580.915 1576.495 ;
        RECT 2580.745 1442.025 2580.915 1490.475 ;
        RECT 2580.745 766.105 2580.915 814.215 ;
        RECT 2580.745 669.545 2580.915 717.655 ;
        RECT 2580.745 572.645 2580.915 620.755 ;
        RECT 2580.745 476.085 2580.915 524.195 ;
        RECT 2580.745 379.525 2580.915 427.635 ;
        RECT 2580.745 282.965 2580.915 331.075 ;
        RECT 2579.825 186.405 2579.995 234.515 ;
        RECT 2580.745 89.845 2580.915 137.955 ;
      LAYER mcon ;
        RECT 2580.745 1576.325 2580.915 1576.495 ;
        RECT 2580.745 1490.305 2580.915 1490.475 ;
        RECT 2580.745 814.045 2580.915 814.215 ;
        RECT 2580.745 717.485 2580.915 717.655 ;
        RECT 2580.745 620.585 2580.915 620.755 ;
        RECT 2580.745 524.025 2580.915 524.195 ;
        RECT 2580.745 427.465 2580.915 427.635 ;
        RECT 2580.745 330.905 2580.915 331.075 ;
        RECT 2579.825 234.345 2579.995 234.515 ;
        RECT 2580.745 137.785 2580.915 137.955 ;
      LAYER met1 ;
        RECT 1850.190 1683.920 1850.510 1683.980 ;
        RECT 1854.330 1683.920 1854.650 1683.980 ;
        RECT 1850.190 1683.780 1854.650 1683.920 ;
        RECT 1850.190 1683.720 1850.510 1683.780 ;
        RECT 1854.330 1683.720 1854.650 1683.780 ;
        RECT 1854.330 1576.480 1854.650 1576.540 ;
        RECT 2580.685 1576.480 2580.975 1576.525 ;
        RECT 1854.330 1576.340 2580.975 1576.480 ;
        RECT 1854.330 1576.280 1854.650 1576.340 ;
        RECT 2580.685 1576.295 2580.975 1576.340 ;
        RECT 2580.670 1539.080 2580.990 1539.140 ;
        RECT 2580.475 1538.940 2580.990 1539.080 ;
        RECT 2580.670 1538.880 2580.990 1538.940 ;
        RECT 2580.670 1490.460 2580.990 1490.520 ;
        RECT 2580.475 1490.320 2580.990 1490.460 ;
        RECT 2580.670 1490.260 2580.990 1490.320 ;
        RECT 2580.670 1442.180 2580.990 1442.240 ;
        RECT 2580.475 1442.040 2580.990 1442.180 ;
        RECT 2580.670 1441.980 2580.990 1442.040 ;
        RECT 2580.670 1345.620 2580.990 1345.680 ;
        RECT 2581.590 1345.620 2581.910 1345.680 ;
        RECT 2580.670 1345.480 2581.910 1345.620 ;
        RECT 2580.670 1345.420 2580.990 1345.480 ;
        RECT 2581.590 1345.420 2581.910 1345.480 ;
        RECT 2580.670 1249.060 2580.990 1249.120 ;
        RECT 2581.590 1249.060 2581.910 1249.120 ;
        RECT 2580.670 1248.920 2581.910 1249.060 ;
        RECT 2580.670 1248.860 2580.990 1248.920 ;
        RECT 2581.590 1248.860 2581.910 1248.920 ;
        RECT 2580.670 1152.500 2580.990 1152.560 ;
        RECT 2581.590 1152.500 2581.910 1152.560 ;
        RECT 2580.670 1152.360 2581.910 1152.500 ;
        RECT 2580.670 1152.300 2580.990 1152.360 ;
        RECT 2581.590 1152.300 2581.910 1152.360 ;
        RECT 2580.670 1007.320 2580.990 1007.380 ;
        RECT 2581.590 1007.320 2581.910 1007.380 ;
        RECT 2580.670 1007.180 2581.910 1007.320 ;
        RECT 2580.670 1007.120 2580.990 1007.180 ;
        RECT 2581.590 1007.120 2581.910 1007.180 ;
        RECT 2580.670 910.760 2580.990 910.820 ;
        RECT 2581.590 910.760 2581.910 910.820 ;
        RECT 2580.670 910.620 2581.910 910.760 ;
        RECT 2580.670 910.560 2580.990 910.620 ;
        RECT 2581.590 910.560 2581.910 910.620 ;
        RECT 2580.670 814.200 2580.990 814.260 ;
        RECT 2580.475 814.060 2580.990 814.200 ;
        RECT 2580.670 814.000 2580.990 814.060 ;
        RECT 2580.670 766.260 2580.990 766.320 ;
        RECT 2580.475 766.120 2580.990 766.260 ;
        RECT 2580.670 766.060 2580.990 766.120 ;
        RECT 2580.670 717.640 2580.990 717.700 ;
        RECT 2580.475 717.500 2580.990 717.640 ;
        RECT 2580.670 717.440 2580.990 717.500 ;
        RECT 2580.670 669.700 2580.990 669.760 ;
        RECT 2580.475 669.560 2580.990 669.700 ;
        RECT 2580.670 669.500 2580.990 669.560 ;
        RECT 2580.670 620.740 2580.990 620.800 ;
        RECT 2580.475 620.600 2580.990 620.740 ;
        RECT 2580.670 620.540 2580.990 620.600 ;
        RECT 2580.670 572.800 2580.990 572.860 ;
        RECT 2580.475 572.660 2580.990 572.800 ;
        RECT 2580.670 572.600 2580.990 572.660 ;
        RECT 2580.670 524.180 2580.990 524.240 ;
        RECT 2580.475 524.040 2580.990 524.180 ;
        RECT 2580.670 523.980 2580.990 524.040 ;
        RECT 2580.670 476.240 2580.990 476.300 ;
        RECT 2580.475 476.100 2580.990 476.240 ;
        RECT 2580.670 476.040 2580.990 476.100 ;
        RECT 2580.670 427.620 2580.990 427.680 ;
        RECT 2580.475 427.480 2580.990 427.620 ;
        RECT 2580.670 427.420 2580.990 427.480 ;
        RECT 2580.670 379.680 2580.990 379.740 ;
        RECT 2580.475 379.540 2580.990 379.680 ;
        RECT 2580.670 379.480 2580.990 379.540 ;
        RECT 2580.670 331.060 2580.990 331.120 ;
        RECT 2580.475 330.920 2580.990 331.060 ;
        RECT 2580.670 330.860 2580.990 330.920 ;
        RECT 2580.670 283.120 2580.990 283.180 ;
        RECT 2580.475 282.980 2580.990 283.120 ;
        RECT 2580.670 282.920 2580.990 282.980 ;
        RECT 2579.765 234.500 2580.055 234.545 ;
        RECT 2580.670 234.500 2580.990 234.560 ;
        RECT 2579.765 234.360 2580.990 234.500 ;
        RECT 2579.765 234.315 2580.055 234.360 ;
        RECT 2580.670 234.300 2580.990 234.360 ;
        RECT 2579.750 186.560 2580.070 186.620 ;
        RECT 2579.555 186.420 2580.070 186.560 ;
        RECT 2579.750 186.360 2580.070 186.420 ;
        RECT 2580.670 137.940 2580.990 138.000 ;
        RECT 2580.475 137.800 2580.990 137.940 ;
        RECT 2580.670 137.740 2580.990 137.800 ;
        RECT 2580.670 90.000 2580.990 90.060 ;
        RECT 2580.475 89.860 2580.990 90.000 ;
        RECT 2580.670 89.800 2580.990 89.860 ;
        RECT 2580.670 62.260 2580.990 62.520 ;
        RECT 2580.760 62.120 2580.900 62.260 ;
        RECT 2583.890 62.120 2584.210 62.180 ;
        RECT 2580.760 61.980 2584.210 62.120 ;
        RECT 2583.890 61.920 2584.210 61.980 ;
        RECT 2583.890 47.980 2584.210 48.240 ;
        RECT 2583.980 47.560 2584.120 47.980 ;
        RECT 2583.890 47.300 2584.210 47.560 ;
      LAYER via ;
        RECT 1850.220 1683.720 1850.480 1683.980 ;
        RECT 1854.360 1683.720 1854.620 1683.980 ;
        RECT 1854.360 1576.280 1854.620 1576.540 ;
        RECT 2580.700 1538.880 2580.960 1539.140 ;
        RECT 2580.700 1490.260 2580.960 1490.520 ;
        RECT 2580.700 1441.980 2580.960 1442.240 ;
        RECT 2580.700 1345.420 2580.960 1345.680 ;
        RECT 2581.620 1345.420 2581.880 1345.680 ;
        RECT 2580.700 1248.860 2580.960 1249.120 ;
        RECT 2581.620 1248.860 2581.880 1249.120 ;
        RECT 2580.700 1152.300 2580.960 1152.560 ;
        RECT 2581.620 1152.300 2581.880 1152.560 ;
        RECT 2580.700 1007.120 2580.960 1007.380 ;
        RECT 2581.620 1007.120 2581.880 1007.380 ;
        RECT 2580.700 910.560 2580.960 910.820 ;
        RECT 2581.620 910.560 2581.880 910.820 ;
        RECT 2580.700 814.000 2580.960 814.260 ;
        RECT 2580.700 766.060 2580.960 766.320 ;
        RECT 2580.700 717.440 2580.960 717.700 ;
        RECT 2580.700 669.500 2580.960 669.760 ;
        RECT 2580.700 620.540 2580.960 620.800 ;
        RECT 2580.700 572.600 2580.960 572.860 ;
        RECT 2580.700 523.980 2580.960 524.240 ;
        RECT 2580.700 476.040 2580.960 476.300 ;
        RECT 2580.700 427.420 2580.960 427.680 ;
        RECT 2580.700 379.480 2580.960 379.740 ;
        RECT 2580.700 330.860 2580.960 331.120 ;
        RECT 2580.700 282.920 2580.960 283.180 ;
        RECT 2580.700 234.300 2580.960 234.560 ;
        RECT 2579.780 186.360 2580.040 186.620 ;
        RECT 2580.700 137.740 2580.960 138.000 ;
        RECT 2580.700 89.800 2580.960 90.060 ;
        RECT 2580.700 62.260 2580.960 62.520 ;
        RECT 2583.920 61.920 2584.180 62.180 ;
        RECT 2583.920 47.980 2584.180 48.240 ;
        RECT 2583.920 47.300 2584.180 47.560 ;
      LAYER met2 ;
        RECT 1850.210 1700.000 1850.490 1704.000 ;
        RECT 1850.280 1684.010 1850.420 1700.000 ;
        RECT 1850.220 1683.690 1850.480 1684.010 ;
        RECT 1854.360 1683.690 1854.620 1684.010 ;
        RECT 1854.420 1576.570 1854.560 1683.690 ;
        RECT 1854.360 1576.250 1854.620 1576.570 ;
        RECT 2580.700 1538.850 2580.960 1539.170 ;
        RECT 2580.760 1490.550 2580.900 1538.850 ;
        RECT 2580.700 1490.230 2580.960 1490.550 ;
        RECT 2580.700 1441.950 2580.960 1442.270 ;
        RECT 2580.760 1393.845 2580.900 1441.950 ;
        RECT 2580.690 1393.475 2580.970 1393.845 ;
        RECT 2581.610 1393.475 2581.890 1393.845 ;
        RECT 2581.680 1345.710 2581.820 1393.475 ;
        RECT 2580.700 1345.390 2580.960 1345.710 ;
        RECT 2581.620 1345.390 2581.880 1345.710 ;
        RECT 2580.760 1297.285 2580.900 1345.390 ;
        RECT 2580.690 1296.915 2580.970 1297.285 ;
        RECT 2581.610 1296.915 2581.890 1297.285 ;
        RECT 2581.680 1249.150 2581.820 1296.915 ;
        RECT 2580.700 1248.830 2580.960 1249.150 ;
        RECT 2581.620 1248.830 2581.880 1249.150 ;
        RECT 2580.760 1208.885 2580.900 1248.830 ;
        RECT 2580.690 1208.515 2580.970 1208.885 ;
        RECT 2580.690 1207.835 2580.970 1208.205 ;
        RECT 2580.760 1200.725 2580.900 1207.835 ;
        RECT 2580.690 1200.355 2580.970 1200.725 ;
        RECT 2581.610 1200.355 2581.890 1200.725 ;
        RECT 2581.680 1152.590 2581.820 1200.355 ;
        RECT 2580.700 1152.270 2580.960 1152.590 ;
        RECT 2581.620 1152.270 2581.880 1152.590 ;
        RECT 2580.760 1104.165 2580.900 1152.270 ;
        RECT 2580.690 1103.795 2580.970 1104.165 ;
        RECT 2581.610 1103.795 2581.890 1104.165 ;
        RECT 2581.680 1055.885 2581.820 1103.795 ;
        RECT 2580.690 1055.515 2580.970 1055.885 ;
        RECT 2581.610 1055.515 2581.890 1055.885 ;
        RECT 2580.760 1007.410 2580.900 1055.515 ;
        RECT 2580.700 1007.090 2580.960 1007.410 ;
        RECT 2581.620 1007.090 2581.880 1007.410 ;
        RECT 2581.680 959.325 2581.820 1007.090 ;
        RECT 2580.690 958.955 2580.970 959.325 ;
        RECT 2581.610 958.955 2581.890 959.325 ;
        RECT 2580.760 910.850 2580.900 958.955 ;
        RECT 2580.700 910.530 2580.960 910.850 ;
        RECT 2581.620 910.530 2581.880 910.850 ;
        RECT 2581.680 862.765 2581.820 910.530 ;
        RECT 2580.690 862.395 2580.970 862.765 ;
        RECT 2581.610 862.395 2581.890 862.765 ;
        RECT 2580.760 821.965 2580.900 862.395 ;
        RECT 2580.690 821.595 2580.970 821.965 ;
        RECT 2580.690 820.915 2580.970 821.285 ;
        RECT 2580.760 814.290 2580.900 820.915 ;
        RECT 2580.700 813.970 2580.960 814.290 ;
        RECT 2580.700 766.030 2580.960 766.350 ;
        RECT 2580.760 717.730 2580.900 766.030 ;
        RECT 2580.700 717.410 2580.960 717.730 ;
        RECT 2580.700 669.470 2580.960 669.790 ;
        RECT 2580.760 620.830 2580.900 669.470 ;
        RECT 2580.700 620.510 2580.960 620.830 ;
        RECT 2580.700 572.570 2580.960 572.890 ;
        RECT 2580.760 524.270 2580.900 572.570 ;
        RECT 2580.700 523.950 2580.960 524.270 ;
        RECT 2580.700 476.010 2580.960 476.330 ;
        RECT 2580.760 427.710 2580.900 476.010 ;
        RECT 2580.700 427.390 2580.960 427.710 ;
        RECT 2580.700 379.450 2580.960 379.770 ;
        RECT 2580.760 331.150 2580.900 379.450 ;
        RECT 2580.700 330.830 2580.960 331.150 ;
        RECT 2580.700 282.890 2580.960 283.210 ;
        RECT 2580.760 234.590 2580.900 282.890 ;
        RECT 2580.700 234.270 2580.960 234.590 ;
        RECT 2579.780 186.330 2580.040 186.650 ;
        RECT 2579.840 145.365 2579.980 186.330 ;
        RECT 2579.770 144.995 2580.050 145.365 ;
        RECT 2580.690 144.995 2580.970 145.365 ;
        RECT 2580.760 138.030 2580.900 144.995 ;
        RECT 2580.700 137.710 2580.960 138.030 ;
        RECT 2580.700 89.770 2580.960 90.090 ;
        RECT 2580.760 62.550 2580.900 89.770 ;
        RECT 2580.700 62.230 2580.960 62.550 ;
        RECT 2583.920 61.890 2584.180 62.210 ;
        RECT 2583.980 48.270 2584.120 61.890 ;
        RECT 2583.920 47.950 2584.180 48.270 ;
        RECT 2583.920 47.270 2584.180 47.590 ;
        RECT 2583.980 2.400 2584.120 47.270 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
      LAYER via2 ;
        RECT 2580.690 1393.520 2580.970 1393.800 ;
        RECT 2581.610 1393.520 2581.890 1393.800 ;
        RECT 2580.690 1296.960 2580.970 1297.240 ;
        RECT 2581.610 1296.960 2581.890 1297.240 ;
        RECT 2580.690 1208.560 2580.970 1208.840 ;
        RECT 2580.690 1207.880 2580.970 1208.160 ;
        RECT 2580.690 1200.400 2580.970 1200.680 ;
        RECT 2581.610 1200.400 2581.890 1200.680 ;
        RECT 2580.690 1103.840 2580.970 1104.120 ;
        RECT 2581.610 1103.840 2581.890 1104.120 ;
        RECT 2580.690 1055.560 2580.970 1055.840 ;
        RECT 2581.610 1055.560 2581.890 1055.840 ;
        RECT 2580.690 959.000 2580.970 959.280 ;
        RECT 2581.610 959.000 2581.890 959.280 ;
        RECT 2580.690 862.440 2580.970 862.720 ;
        RECT 2581.610 862.440 2581.890 862.720 ;
        RECT 2580.690 821.640 2580.970 821.920 ;
        RECT 2580.690 820.960 2580.970 821.240 ;
        RECT 2579.770 145.040 2580.050 145.320 ;
        RECT 2580.690 145.040 2580.970 145.320 ;
      LAYER met3 ;
        RECT 2580.665 1393.810 2580.995 1393.825 ;
        RECT 2581.585 1393.810 2581.915 1393.825 ;
        RECT 2580.665 1393.510 2581.915 1393.810 ;
        RECT 2580.665 1393.495 2580.995 1393.510 ;
        RECT 2581.585 1393.495 2581.915 1393.510 ;
        RECT 2580.665 1297.250 2580.995 1297.265 ;
        RECT 2581.585 1297.250 2581.915 1297.265 ;
        RECT 2580.665 1296.950 2581.915 1297.250 ;
        RECT 2580.665 1296.935 2580.995 1296.950 ;
        RECT 2581.585 1296.935 2581.915 1296.950 ;
        RECT 2580.665 1208.850 2580.995 1208.865 ;
        RECT 2579.990 1208.550 2580.995 1208.850 ;
        RECT 2579.990 1208.170 2580.290 1208.550 ;
        RECT 2580.665 1208.535 2580.995 1208.550 ;
        RECT 2580.665 1208.170 2580.995 1208.185 ;
        RECT 2579.990 1207.870 2580.995 1208.170 ;
        RECT 2580.665 1207.855 2580.995 1207.870 ;
        RECT 2580.665 1200.690 2580.995 1200.705 ;
        RECT 2581.585 1200.690 2581.915 1200.705 ;
        RECT 2580.665 1200.390 2581.915 1200.690 ;
        RECT 2580.665 1200.375 2580.995 1200.390 ;
        RECT 2581.585 1200.375 2581.915 1200.390 ;
        RECT 2580.665 1104.130 2580.995 1104.145 ;
        RECT 2581.585 1104.130 2581.915 1104.145 ;
        RECT 2580.665 1103.830 2581.915 1104.130 ;
        RECT 2580.665 1103.815 2580.995 1103.830 ;
        RECT 2581.585 1103.815 2581.915 1103.830 ;
        RECT 2580.665 1055.850 2580.995 1055.865 ;
        RECT 2581.585 1055.850 2581.915 1055.865 ;
        RECT 2580.665 1055.550 2581.915 1055.850 ;
        RECT 2580.665 1055.535 2580.995 1055.550 ;
        RECT 2581.585 1055.535 2581.915 1055.550 ;
        RECT 2580.665 959.290 2580.995 959.305 ;
        RECT 2581.585 959.290 2581.915 959.305 ;
        RECT 2580.665 958.990 2581.915 959.290 ;
        RECT 2580.665 958.975 2580.995 958.990 ;
        RECT 2581.585 958.975 2581.915 958.990 ;
        RECT 2580.665 862.730 2580.995 862.745 ;
        RECT 2581.585 862.730 2581.915 862.745 ;
        RECT 2580.665 862.430 2581.915 862.730 ;
        RECT 2580.665 862.415 2580.995 862.430 ;
        RECT 2581.585 862.415 2581.915 862.430 ;
        RECT 2580.665 821.930 2580.995 821.945 ;
        RECT 2579.990 821.630 2580.995 821.930 ;
        RECT 2579.990 821.250 2580.290 821.630 ;
        RECT 2580.665 821.615 2580.995 821.630 ;
        RECT 2580.665 821.250 2580.995 821.265 ;
        RECT 2579.990 820.950 2580.995 821.250 ;
        RECT 2580.665 820.935 2580.995 820.950 ;
        RECT 2579.745 145.330 2580.075 145.345 ;
        RECT 2580.665 145.330 2580.995 145.345 ;
        RECT 2579.745 145.030 2580.995 145.330 ;
        RECT 2579.745 145.015 2580.075 145.030 ;
        RECT 2580.665 145.015 2580.995 145.030 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1366.270 1678.140 1366.590 1678.200 ;
        RECT 1369.030 1678.140 1369.350 1678.200 ;
        RECT 1366.270 1678.000 1369.350 1678.140 ;
        RECT 1366.270 1677.940 1366.590 1678.000 ;
        RECT 1369.030 1677.940 1369.350 1678.000 ;
        RECT 817.490 31.860 817.810 31.920 ;
        RECT 1366.270 31.860 1366.590 31.920 ;
        RECT 817.490 31.720 1366.590 31.860 ;
        RECT 817.490 31.660 817.810 31.720 ;
        RECT 1366.270 31.660 1366.590 31.720 ;
      LAYER via ;
        RECT 1366.300 1677.940 1366.560 1678.200 ;
        RECT 1369.060 1677.940 1369.320 1678.200 ;
        RECT 817.520 31.660 817.780 31.920 ;
        RECT 1366.300 31.660 1366.560 31.920 ;
      LAYER met2 ;
        RECT 1370.430 1700.410 1370.710 1704.000 ;
        RECT 1369.120 1700.270 1370.710 1700.410 ;
        RECT 1369.120 1678.230 1369.260 1700.270 ;
        RECT 1370.430 1700.000 1370.710 1700.270 ;
        RECT 1366.300 1677.910 1366.560 1678.230 ;
        RECT 1369.060 1677.910 1369.320 1678.230 ;
        RECT 1366.360 31.950 1366.500 1677.910 ;
        RECT 817.520 31.630 817.780 31.950 ;
        RECT 1366.300 31.630 1366.560 31.950 ;
        RECT 817.580 2.400 817.720 31.630 ;
=======
      LAYER li1 ;
        RECT 1368.185 1497.785 1368.355 1555.755 ;
        RECT 1368.185 1400.885 1368.355 1490.475 ;
        RECT 1368.185 1297.185 1368.355 1345.295 ;
        RECT 1368.185 1041.165 1368.355 1083.155 ;
        RECT 1368.645 848.725 1368.815 882.555 ;
        RECT 1369.105 752.165 1369.275 800.275 ;
        RECT 1368.185 614.125 1368.355 662.235 ;
        RECT 1368.185 565.505 1368.355 590.155 ;
        RECT 1368.645 476.085 1368.815 517.735 ;
        RECT 1368.645 343.485 1368.815 386.155 ;
        RECT 1368.645 276.505 1368.815 292.315 ;
        RECT 1368.185 227.885 1368.355 275.995 ;
        RECT 1368.185 138.125 1368.355 186.235 ;
        RECT 1368.185 89.845 1368.355 113.815 ;
      LAYER mcon ;
        RECT 1368.185 1555.585 1368.355 1555.755 ;
        RECT 1368.185 1490.305 1368.355 1490.475 ;
        RECT 1368.185 1345.125 1368.355 1345.295 ;
        RECT 1368.185 1082.985 1368.355 1083.155 ;
        RECT 1368.645 882.385 1368.815 882.555 ;
        RECT 1369.105 800.105 1369.275 800.275 ;
        RECT 1368.185 662.065 1368.355 662.235 ;
        RECT 1368.185 589.985 1368.355 590.155 ;
        RECT 1368.645 517.565 1368.815 517.735 ;
        RECT 1368.645 385.985 1368.815 386.155 ;
        RECT 1368.645 292.145 1368.815 292.315 ;
        RECT 1368.185 275.825 1368.355 275.995 ;
        RECT 1368.185 186.065 1368.355 186.235 ;
        RECT 1368.185 113.645 1368.355 113.815 ;
      LAYER met1 ;
        RECT 1368.125 1555.740 1368.415 1555.785 ;
        RECT 1368.570 1555.740 1368.890 1555.800 ;
        RECT 1368.125 1555.600 1368.890 1555.740 ;
        RECT 1368.125 1555.555 1368.415 1555.600 ;
        RECT 1368.570 1555.540 1368.890 1555.600 ;
        RECT 1368.110 1497.940 1368.430 1498.000 ;
        RECT 1367.915 1497.800 1368.430 1497.940 ;
        RECT 1368.110 1497.740 1368.430 1497.800 ;
        RECT 1368.110 1490.460 1368.430 1490.520 ;
        RECT 1367.915 1490.320 1368.430 1490.460 ;
        RECT 1368.110 1490.260 1368.430 1490.320 ;
        RECT 1368.110 1401.040 1368.430 1401.100 ;
        RECT 1367.915 1400.900 1368.430 1401.040 ;
        RECT 1368.110 1400.840 1368.430 1400.900 ;
        RECT 1368.110 1352.760 1368.430 1352.820 ;
        RECT 1368.570 1352.760 1368.890 1352.820 ;
        RECT 1368.110 1352.620 1368.890 1352.760 ;
        RECT 1368.110 1352.560 1368.430 1352.620 ;
        RECT 1368.570 1352.560 1368.890 1352.620 ;
        RECT 1368.125 1345.280 1368.415 1345.325 ;
        RECT 1368.570 1345.280 1368.890 1345.340 ;
        RECT 1368.125 1345.140 1368.890 1345.280 ;
        RECT 1368.125 1345.095 1368.415 1345.140 ;
        RECT 1368.570 1345.080 1368.890 1345.140 ;
        RECT 1368.110 1297.340 1368.430 1297.400 ;
        RECT 1367.915 1297.200 1368.430 1297.340 ;
        RECT 1368.110 1297.140 1368.430 1297.200 ;
        RECT 1368.110 1273.680 1368.430 1273.940 ;
        RECT 1368.200 1273.260 1368.340 1273.680 ;
        RECT 1368.110 1273.000 1368.430 1273.260 ;
        RECT 1368.110 1201.260 1368.430 1201.520 ;
        RECT 1368.200 1200.840 1368.340 1201.260 ;
        RECT 1368.110 1200.580 1368.430 1200.840 ;
        RECT 1368.110 1145.500 1368.430 1145.760 ;
        RECT 1368.200 1145.080 1368.340 1145.500 ;
        RECT 1368.110 1144.820 1368.430 1145.080 ;
        RECT 1368.110 1083.140 1368.430 1083.200 ;
        RECT 1367.915 1083.000 1368.430 1083.140 ;
        RECT 1368.110 1082.940 1368.430 1083.000 ;
        RECT 1368.125 1041.320 1368.415 1041.365 ;
        RECT 1369.030 1041.320 1369.350 1041.380 ;
        RECT 1368.125 1041.180 1369.350 1041.320 ;
        RECT 1368.125 1041.135 1368.415 1041.180 ;
        RECT 1369.030 1041.120 1369.350 1041.180 ;
        RECT 1368.110 979.920 1368.430 980.180 ;
        RECT 1368.200 979.440 1368.340 979.920 ;
        RECT 1368.570 979.440 1368.890 979.500 ;
        RECT 1368.200 979.300 1368.890 979.440 ;
        RECT 1368.570 979.240 1368.890 979.300 ;
        RECT 1368.570 938.100 1368.890 938.360 ;
        RECT 1368.660 937.960 1368.800 938.100 ;
        RECT 1369.030 937.960 1369.350 938.020 ;
        RECT 1368.660 937.820 1369.350 937.960 ;
        RECT 1369.030 937.760 1369.350 937.820 ;
        RECT 1368.585 882.540 1368.875 882.585 ;
        RECT 1369.030 882.540 1369.350 882.600 ;
        RECT 1368.585 882.400 1369.350 882.540 ;
        RECT 1368.585 882.355 1368.875 882.400 ;
        RECT 1369.030 882.340 1369.350 882.400 ;
        RECT 1368.570 848.880 1368.890 848.940 ;
        RECT 1368.375 848.740 1368.890 848.880 ;
        RECT 1368.570 848.680 1368.890 848.740 ;
        RECT 1368.570 800.260 1368.890 800.320 ;
        RECT 1369.045 800.260 1369.335 800.305 ;
        RECT 1368.570 800.120 1369.335 800.260 ;
        RECT 1368.570 800.060 1368.890 800.120 ;
        RECT 1369.045 800.075 1369.335 800.120 ;
        RECT 1368.570 752.320 1368.890 752.380 ;
        RECT 1369.045 752.320 1369.335 752.365 ;
        RECT 1368.570 752.180 1369.335 752.320 ;
        RECT 1368.570 752.120 1368.890 752.180 ;
        RECT 1369.045 752.135 1369.335 752.180 ;
        RECT 1368.125 662.220 1368.415 662.265 ;
        RECT 1368.570 662.220 1368.890 662.280 ;
        RECT 1368.125 662.080 1368.890 662.220 ;
        RECT 1368.125 662.035 1368.415 662.080 ;
        RECT 1368.570 662.020 1368.890 662.080 ;
        RECT 1368.110 614.280 1368.430 614.340 ;
        RECT 1367.915 614.140 1368.430 614.280 ;
        RECT 1368.110 614.080 1368.430 614.140 ;
        RECT 1368.125 590.140 1368.415 590.185 ;
        RECT 1368.570 590.140 1368.890 590.200 ;
        RECT 1368.125 590.000 1368.890 590.140 ;
        RECT 1368.125 589.955 1368.415 590.000 ;
        RECT 1368.570 589.940 1368.890 590.000 ;
        RECT 1368.110 565.660 1368.430 565.720 ;
        RECT 1367.915 565.520 1368.430 565.660 ;
        RECT 1368.110 565.460 1368.430 565.520 ;
        RECT 1368.110 518.060 1368.430 518.120 ;
        RECT 1368.110 517.920 1368.800 518.060 ;
        RECT 1368.110 517.860 1368.430 517.920 ;
        RECT 1368.660 517.765 1368.800 517.920 ;
        RECT 1368.585 517.535 1368.875 517.765 ;
        RECT 1368.570 476.240 1368.890 476.300 ;
        RECT 1368.375 476.100 1368.890 476.240 ;
        RECT 1368.570 476.040 1368.890 476.100 ;
        RECT 1368.570 386.140 1368.890 386.200 ;
        RECT 1368.375 386.000 1368.890 386.140 ;
        RECT 1368.570 385.940 1368.890 386.000 ;
        RECT 1368.570 343.640 1368.890 343.700 ;
        RECT 1368.375 343.500 1368.890 343.640 ;
        RECT 1368.570 343.440 1368.890 343.500 ;
        RECT 1368.570 292.300 1368.890 292.360 ;
        RECT 1368.375 292.160 1368.890 292.300 ;
        RECT 1368.570 292.100 1368.890 292.160 ;
        RECT 1368.570 276.660 1368.890 276.720 ;
        RECT 1368.375 276.520 1368.890 276.660 ;
        RECT 1368.570 276.460 1368.890 276.520 ;
        RECT 1368.110 275.980 1368.430 276.040 ;
        RECT 1367.915 275.840 1368.430 275.980 ;
        RECT 1368.110 275.780 1368.430 275.840 ;
        RECT 1368.110 228.040 1368.430 228.100 ;
        RECT 1367.915 227.900 1368.430 228.040 ;
        RECT 1368.110 227.840 1368.430 227.900 ;
        RECT 1368.125 186.220 1368.415 186.265 ;
        RECT 1368.570 186.220 1368.890 186.280 ;
        RECT 1368.125 186.080 1368.890 186.220 ;
        RECT 1368.125 186.035 1368.415 186.080 ;
        RECT 1368.570 186.020 1368.890 186.080 ;
        RECT 1368.110 138.280 1368.430 138.340 ;
        RECT 1367.915 138.140 1368.430 138.280 ;
        RECT 1368.110 138.080 1368.430 138.140 ;
        RECT 1368.110 113.800 1368.430 113.860 ;
        RECT 1367.915 113.660 1368.430 113.800 ;
        RECT 1368.110 113.600 1368.430 113.660 ;
        RECT 1368.125 90.000 1368.415 90.045 ;
        RECT 1368.570 90.000 1368.890 90.060 ;
        RECT 1368.125 89.860 1368.890 90.000 ;
        RECT 1368.125 89.815 1368.415 89.860 ;
        RECT 1368.570 89.800 1368.890 89.860 ;
        RECT 817.490 32.200 817.810 32.260 ;
        RECT 1368.570 32.200 1368.890 32.260 ;
        RECT 817.490 32.060 1368.890 32.200 ;
        RECT 817.490 32.000 817.810 32.060 ;
        RECT 1368.570 32.000 1368.890 32.060 ;
      LAYER via ;
        RECT 1368.600 1555.540 1368.860 1555.800 ;
        RECT 1368.140 1497.740 1368.400 1498.000 ;
        RECT 1368.140 1490.260 1368.400 1490.520 ;
        RECT 1368.140 1400.840 1368.400 1401.100 ;
        RECT 1368.140 1352.560 1368.400 1352.820 ;
        RECT 1368.600 1352.560 1368.860 1352.820 ;
        RECT 1368.600 1345.080 1368.860 1345.340 ;
        RECT 1368.140 1297.140 1368.400 1297.400 ;
        RECT 1368.140 1273.680 1368.400 1273.940 ;
        RECT 1368.140 1273.000 1368.400 1273.260 ;
        RECT 1368.140 1201.260 1368.400 1201.520 ;
        RECT 1368.140 1200.580 1368.400 1200.840 ;
        RECT 1368.140 1145.500 1368.400 1145.760 ;
        RECT 1368.140 1144.820 1368.400 1145.080 ;
        RECT 1368.140 1082.940 1368.400 1083.200 ;
        RECT 1369.060 1041.120 1369.320 1041.380 ;
        RECT 1368.140 979.920 1368.400 980.180 ;
        RECT 1368.600 979.240 1368.860 979.500 ;
        RECT 1368.600 938.100 1368.860 938.360 ;
        RECT 1369.060 937.760 1369.320 938.020 ;
        RECT 1369.060 882.340 1369.320 882.600 ;
        RECT 1368.600 848.680 1368.860 848.940 ;
        RECT 1368.600 800.060 1368.860 800.320 ;
        RECT 1368.600 752.120 1368.860 752.380 ;
        RECT 1368.600 662.020 1368.860 662.280 ;
        RECT 1368.140 614.080 1368.400 614.340 ;
        RECT 1368.600 589.940 1368.860 590.200 ;
        RECT 1368.140 565.460 1368.400 565.720 ;
        RECT 1368.140 517.860 1368.400 518.120 ;
        RECT 1368.600 476.040 1368.860 476.300 ;
        RECT 1368.600 385.940 1368.860 386.200 ;
        RECT 1368.600 343.440 1368.860 343.700 ;
        RECT 1368.600 292.100 1368.860 292.360 ;
        RECT 1368.600 276.460 1368.860 276.720 ;
        RECT 1368.140 275.780 1368.400 276.040 ;
        RECT 1368.140 227.840 1368.400 228.100 ;
        RECT 1368.600 186.020 1368.860 186.280 ;
        RECT 1368.140 138.080 1368.400 138.340 ;
        RECT 1368.140 113.600 1368.400 113.860 ;
        RECT 1368.600 89.800 1368.860 90.060 ;
        RECT 817.520 32.000 817.780 32.260 ;
        RECT 1368.600 32.000 1368.860 32.260 ;
      LAYER met2 ;
        RECT 1371.350 1700.410 1371.630 1704.000 ;
        RECT 1370.040 1700.270 1371.630 1700.410 ;
        RECT 1370.040 1678.140 1370.180 1700.270 ;
        RECT 1371.350 1700.000 1371.630 1700.270 ;
        RECT 1368.660 1678.000 1370.180 1678.140 ;
        RECT 1368.660 1555.830 1368.800 1678.000 ;
        RECT 1368.600 1555.510 1368.860 1555.830 ;
        RECT 1368.140 1497.710 1368.400 1498.030 ;
        RECT 1368.200 1490.550 1368.340 1497.710 ;
        RECT 1368.140 1490.230 1368.400 1490.550 ;
        RECT 1368.140 1400.810 1368.400 1401.130 ;
        RECT 1368.200 1352.850 1368.340 1400.810 ;
        RECT 1368.140 1352.530 1368.400 1352.850 ;
        RECT 1368.600 1352.530 1368.860 1352.850 ;
        RECT 1368.660 1345.370 1368.800 1352.530 ;
        RECT 1368.600 1345.050 1368.860 1345.370 ;
        RECT 1368.140 1297.110 1368.400 1297.430 ;
        RECT 1368.200 1273.970 1368.340 1297.110 ;
        RECT 1368.140 1273.650 1368.400 1273.970 ;
        RECT 1368.140 1272.970 1368.400 1273.290 ;
        RECT 1368.200 1201.550 1368.340 1272.970 ;
        RECT 1368.140 1201.230 1368.400 1201.550 ;
        RECT 1368.140 1200.550 1368.400 1200.870 ;
        RECT 1368.200 1145.790 1368.340 1200.550 ;
        RECT 1368.140 1145.470 1368.400 1145.790 ;
        RECT 1368.140 1144.790 1368.400 1145.110 ;
        RECT 1368.200 1083.230 1368.340 1144.790 ;
        RECT 1368.140 1082.910 1368.400 1083.230 ;
        RECT 1369.060 1041.090 1369.320 1041.410 ;
        RECT 1369.120 1017.690 1369.260 1041.090 ;
        RECT 1368.200 1017.550 1369.260 1017.690 ;
        RECT 1368.200 980.210 1368.340 1017.550 ;
        RECT 1368.140 979.890 1368.400 980.210 ;
        RECT 1368.600 979.210 1368.860 979.530 ;
        RECT 1368.660 938.390 1368.800 979.210 ;
        RECT 1368.600 938.070 1368.860 938.390 ;
        RECT 1369.060 937.730 1369.320 938.050 ;
        RECT 1369.120 882.630 1369.260 937.730 ;
        RECT 1369.060 882.310 1369.320 882.630 ;
        RECT 1368.600 848.650 1368.860 848.970 ;
        RECT 1368.660 800.350 1368.800 848.650 ;
        RECT 1368.600 800.030 1368.860 800.350 ;
        RECT 1368.600 752.090 1368.860 752.410 ;
        RECT 1368.660 734.810 1368.800 752.090 ;
        RECT 1368.200 734.670 1368.800 734.810 ;
        RECT 1368.200 686.530 1368.340 734.670 ;
        RECT 1368.200 686.390 1368.800 686.530 ;
        RECT 1368.660 662.310 1368.800 686.390 ;
        RECT 1368.600 661.990 1368.860 662.310 ;
        RECT 1368.140 614.050 1368.400 614.370 ;
        RECT 1368.200 613.770 1368.340 614.050 ;
        RECT 1368.200 613.630 1368.800 613.770 ;
        RECT 1368.660 590.230 1368.800 613.630 ;
        RECT 1368.600 589.910 1368.860 590.230 ;
        RECT 1368.140 565.430 1368.400 565.750 ;
        RECT 1368.200 518.150 1368.340 565.430 ;
        RECT 1368.140 517.830 1368.400 518.150 ;
        RECT 1368.600 476.010 1368.860 476.330 ;
        RECT 1368.660 386.230 1368.800 476.010 ;
        RECT 1368.600 385.910 1368.860 386.230 ;
        RECT 1368.600 343.410 1368.860 343.730 ;
        RECT 1368.660 292.390 1368.800 343.410 ;
        RECT 1368.600 292.070 1368.860 292.390 ;
        RECT 1368.600 276.490 1368.860 276.750 ;
        RECT 1368.200 276.430 1368.860 276.490 ;
        RECT 1368.200 276.350 1368.800 276.430 ;
        RECT 1368.200 276.070 1368.340 276.350 ;
        RECT 1368.140 275.750 1368.400 276.070 ;
        RECT 1368.140 227.810 1368.400 228.130 ;
        RECT 1368.200 209.170 1368.340 227.810 ;
        RECT 1368.200 209.030 1368.800 209.170 ;
        RECT 1368.660 186.310 1368.800 209.030 ;
        RECT 1368.600 185.990 1368.860 186.310 ;
        RECT 1368.140 138.050 1368.400 138.370 ;
        RECT 1368.200 113.890 1368.340 138.050 ;
        RECT 1368.140 113.570 1368.400 113.890 ;
        RECT 1368.600 89.770 1368.860 90.090 ;
        RECT 1368.660 32.290 1368.800 89.770 ;
        RECT 817.520 31.970 817.780 32.290 ;
        RECT 1368.600 31.970 1368.860 32.290 ;
        RECT 817.580 2.400 817.720 31.970 ;
>>>>>>> re-updated local openlane
        RECT 817.370 -4.800 817.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1854.790 1569.680 1855.110 1569.740 ;
        RECT 2601.830 1569.680 2602.150 1569.740 ;
        RECT 1854.790 1569.540 2602.150 1569.680 ;
        RECT 1854.790 1569.480 1855.110 1569.540 ;
        RECT 2601.830 1569.480 2602.150 1569.540 ;
      LAYER via ;
        RECT 1854.820 1569.480 1855.080 1569.740 ;
        RECT 2601.860 1569.480 2602.120 1569.740 ;
      LAYER met2 ;
        RECT 1855.270 1700.410 1855.550 1704.000 ;
        RECT 1854.880 1700.270 1855.550 1700.410 ;
        RECT 1854.880 1569.770 1855.020 1700.270 ;
        RECT 1855.270 1700.000 1855.550 1700.270 ;
        RECT 1854.820 1569.450 1855.080 1569.770 ;
        RECT 2601.860 1569.450 2602.120 1569.770 ;
        RECT 2601.920 7.210 2602.060 1569.450 ;
        RECT 2601.460 7.070 2602.060 7.210 ;
        RECT 2601.460 2.400 2601.600 7.070 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1862.150 36.280 1862.470 36.340 ;
        RECT 1862.150 36.140 2596.540 36.280 ;
        RECT 1862.150 36.080 1862.470 36.140 ;
        RECT 2596.400 35.600 2596.540 36.140 ;
        RECT 2619.310 35.600 2619.630 35.660 ;
        RECT 2596.400 35.460 2619.630 35.600 ;
        RECT 2619.310 35.400 2619.630 35.460 ;
      LAYER via ;
        RECT 1862.180 36.080 1862.440 36.340 ;
        RECT 2619.340 35.400 2619.600 35.660 ;
      LAYER met2 ;
        RECT 1859.870 1700.410 1860.150 1704.000 ;
        RECT 1859.870 1700.270 1861.460 1700.410 ;
        RECT 1859.870 1700.000 1860.150 1700.270 ;
        RECT 1861.320 1677.970 1861.460 1700.270 ;
        RECT 1861.320 1677.830 1862.380 1677.970 ;
        RECT 1862.240 36.370 1862.380 1677.830 ;
        RECT 1862.180 36.050 1862.440 36.370 ;
        RECT 2619.340 35.370 2619.600 35.690 ;
        RECT 2619.400 2.400 2619.540 35.370 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1864.910 1683.920 1865.230 1683.980 ;
        RECT 1868.130 1683.920 1868.450 1683.980 ;
        RECT 1864.910 1683.780 1868.450 1683.920 ;
        RECT 1864.910 1683.720 1865.230 1683.780 ;
        RECT 1868.130 1683.720 1868.450 1683.780 ;
        RECT 1868.130 36.620 1868.450 36.680 ;
        RECT 2637.250 36.620 2637.570 36.680 ;
        RECT 1868.130 36.480 2637.570 36.620 ;
        RECT 1868.130 36.420 1868.450 36.480 ;
        RECT 2637.250 36.420 2637.570 36.480 ;
      LAYER via ;
        RECT 1864.940 1683.720 1865.200 1683.980 ;
        RECT 1868.160 1683.720 1868.420 1683.980 ;
        RECT 1868.160 36.420 1868.420 36.680 ;
        RECT 2637.280 36.420 2637.540 36.680 ;
      LAYER met2 ;
        RECT 1864.930 1700.000 1865.210 1704.000 ;
        RECT 1865.000 1684.010 1865.140 1700.000 ;
        RECT 1864.940 1683.690 1865.200 1684.010 ;
        RECT 1868.160 1683.690 1868.420 1684.010 ;
        RECT 1868.220 36.710 1868.360 1683.690 ;
        RECT 1868.160 36.390 1868.420 36.710 ;
        RECT 2637.280 36.390 2637.540 36.710 ;
        RECT 2637.340 2.400 2637.480 36.390 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 0.300 ;
=======
      LAYER met1 ;
        RECT 1868.590 36.960 1868.910 37.020 ;
        RECT 2655.190 36.960 2655.510 37.020 ;
        RECT 1868.590 36.820 2655.510 36.960 ;
        RECT 1868.590 36.760 1868.910 36.820 ;
        RECT 2655.190 36.760 2655.510 36.820 ;
      LAYER via ;
        RECT 1868.620 36.760 1868.880 37.020 ;
        RECT 2655.220 36.760 2655.480 37.020 ;
      LAYER met2 ;
        RECT 1869.530 1700.410 1869.810 1704.000 ;
        RECT 1868.680 1700.270 1869.810 1700.410 ;
        RECT 1868.680 37.050 1868.820 1700.270 ;
        RECT 1869.530 1700.000 1869.810 1700.270 ;
        RECT 1868.620 36.730 1868.880 37.050 ;
        RECT 2655.220 36.730 2655.480 37.050 ;
        RECT 2655.280 2.400 2655.420 36.730 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1874.570 1684.600 1874.890 1684.660 ;
        RECT 1875.950 1684.600 1876.270 1684.660 ;
        RECT 1874.570 1684.460 1876.270 1684.600 ;
        RECT 1874.570 1684.400 1874.890 1684.460 ;
        RECT 1875.950 1684.400 1876.270 1684.460 ;
        RECT 1875.950 37.300 1876.270 37.360 ;
        RECT 2672.670 37.300 2672.990 37.360 ;
        RECT 1875.950 37.160 2672.990 37.300 ;
        RECT 1875.950 37.100 1876.270 37.160 ;
        RECT 2672.670 37.100 2672.990 37.160 ;
      LAYER via ;
        RECT 1874.600 1684.400 1874.860 1684.660 ;
        RECT 1875.980 1684.400 1876.240 1684.660 ;
        RECT 1875.980 37.100 1876.240 37.360 ;
        RECT 2672.700 37.100 2672.960 37.360 ;
      LAYER met2 ;
        RECT 1874.590 1700.000 1874.870 1704.000 ;
        RECT 1874.660 1684.690 1874.800 1700.000 ;
        RECT 1874.600 1684.370 1874.860 1684.690 ;
        RECT 1875.980 1684.370 1876.240 1684.690 ;
        RECT 1876.040 37.390 1876.180 1684.370 ;
        RECT 1875.980 37.070 1876.240 37.390 ;
        RECT 2672.700 37.070 2672.960 37.390 ;
        RECT 2672.760 2.400 2672.900 37.070 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1879.170 1683.920 1879.490 1683.980 ;
        RECT 1882.390 1683.920 1882.710 1683.980 ;
        RECT 1879.170 1683.780 1882.710 1683.920 ;
        RECT 1879.170 1683.720 1879.490 1683.780 ;
        RECT 1882.390 1683.720 1882.710 1683.780 ;
        RECT 1882.390 37.640 1882.710 37.700 ;
        RECT 2690.610 37.640 2690.930 37.700 ;
        RECT 1882.390 37.500 2690.930 37.640 ;
        RECT 1882.390 37.440 1882.710 37.500 ;
        RECT 2690.610 37.440 2690.930 37.500 ;
      LAYER via ;
        RECT 1879.200 1683.720 1879.460 1683.980 ;
        RECT 1882.420 1683.720 1882.680 1683.980 ;
        RECT 1882.420 37.440 1882.680 37.700 ;
        RECT 2690.640 37.440 2690.900 37.700 ;
      LAYER met2 ;
        RECT 1879.190 1700.000 1879.470 1704.000 ;
        RECT 1879.260 1684.010 1879.400 1700.000 ;
        RECT 1879.200 1683.690 1879.460 1684.010 ;
        RECT 1882.420 1683.690 1882.680 1684.010 ;
        RECT 1882.480 37.730 1882.620 1683.690 ;
        RECT 1882.420 37.410 1882.680 37.730 ;
        RECT 2690.640 37.410 2690.900 37.730 ;
        RECT 2690.700 2.400 2690.840 37.410 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1884.230 1684.600 1884.550 1684.660 ;
        RECT 1889.290 1684.600 1889.610 1684.660 ;
        RECT 1884.230 1684.460 1889.610 1684.600 ;
        RECT 1884.230 1684.400 1884.550 1684.460 ;
        RECT 1889.290 1684.400 1889.610 1684.460 ;
        RECT 1889.290 41.380 1889.610 41.440 ;
        RECT 2708.550 41.380 2708.870 41.440 ;
        RECT 1889.290 41.240 2708.870 41.380 ;
        RECT 1889.290 41.180 1889.610 41.240 ;
        RECT 2708.550 41.180 2708.870 41.240 ;
      LAYER via ;
        RECT 1884.260 1684.400 1884.520 1684.660 ;
        RECT 1889.320 1684.400 1889.580 1684.660 ;
        RECT 1889.320 41.180 1889.580 41.440 ;
        RECT 2708.580 41.180 2708.840 41.440 ;
      LAYER met2 ;
        RECT 1884.250 1700.000 1884.530 1704.000 ;
        RECT 1884.320 1684.690 1884.460 1700.000 ;
        RECT 1884.260 1684.370 1884.520 1684.690 ;
        RECT 1889.320 1684.370 1889.580 1684.690 ;
        RECT 1889.380 41.470 1889.520 1684.370 ;
        RECT 1889.320 41.150 1889.580 41.470 ;
        RECT 2708.580 41.150 2708.840 41.470 ;
        RECT 2708.640 2.400 2708.780 41.150 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1888.830 41.040 1889.150 41.100 ;
        RECT 2726.490 41.040 2726.810 41.100 ;
        RECT 1888.830 40.900 2726.810 41.040 ;
        RECT 1888.830 40.840 1889.150 40.900 ;
        RECT 2726.490 40.840 2726.810 40.900 ;
      LAYER via ;
        RECT 1888.860 40.840 1889.120 41.100 ;
        RECT 2726.520 40.840 2726.780 41.100 ;
      LAYER met2 ;
        RECT 1888.850 1700.000 1889.130 1704.000 ;
        RECT 1888.920 41.130 1889.060 1700.000 ;
        RECT 1888.860 40.810 1889.120 41.130 ;
        RECT 2726.520 40.810 2726.780 41.130 ;
        RECT 2726.580 2.400 2726.720 40.810 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 0.300 ;
=======
      LAYER met1 ;
        RECT 1895.270 40.700 1895.590 40.760 ;
        RECT 2744.430 40.700 2744.750 40.760 ;
        RECT 1895.270 40.560 2744.750 40.700 ;
        RECT 1895.270 40.500 1895.590 40.560 ;
        RECT 2744.430 40.500 2744.750 40.560 ;
      LAYER via ;
        RECT 1895.300 40.500 1895.560 40.760 ;
        RECT 2744.460 40.500 2744.720 40.760 ;
      LAYER met2 ;
        RECT 1893.910 1700.410 1894.190 1704.000 ;
        RECT 1893.910 1700.270 1894.580 1700.410 ;
        RECT 1893.910 1700.000 1894.190 1700.270 ;
        RECT 1894.440 1656.210 1894.580 1700.270 ;
        RECT 1894.440 1656.070 1895.500 1656.210 ;
        RECT 1895.360 40.790 1895.500 1656.070 ;
        RECT 1895.300 40.470 1895.560 40.790 ;
        RECT 2744.460 40.470 2744.720 40.790 ;
        RECT 2744.520 2.400 2744.660 40.470 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1898.490 1683.920 1898.810 1683.980 ;
        RECT 1902.630 1683.920 1902.950 1683.980 ;
        RECT 1898.490 1683.780 1902.950 1683.920 ;
        RECT 1898.490 1683.720 1898.810 1683.780 ;
        RECT 1902.630 1683.720 1902.950 1683.780 ;
        RECT 1902.630 40.360 1902.950 40.420 ;
        RECT 2761.910 40.360 2762.230 40.420 ;
        RECT 1902.630 40.220 2762.230 40.360 ;
        RECT 1902.630 40.160 1902.950 40.220 ;
        RECT 2761.910 40.160 2762.230 40.220 ;
      LAYER via ;
        RECT 1898.520 1683.720 1898.780 1683.980 ;
        RECT 1902.660 1683.720 1902.920 1683.980 ;
        RECT 1902.660 40.160 1902.920 40.420 ;
        RECT 2761.940 40.160 2762.200 40.420 ;
      LAYER met2 ;
        RECT 1898.510 1700.000 1898.790 1704.000 ;
        RECT 1898.580 1684.010 1898.720 1700.000 ;
        RECT 1898.520 1683.690 1898.780 1684.010 ;
        RECT 1902.660 1683.690 1902.920 1684.010 ;
        RECT 1902.720 40.450 1902.860 1683.690 ;
        RECT 1902.660 40.130 1902.920 40.450 ;
        RECT 2761.940 40.130 2762.200 40.450 ;
        RECT 2762.000 2.400 2762.140 40.130 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 0.300 ;
=======
      LAYER met1 ;
        RECT 835.430 32.540 835.750 32.600 ;
        RECT 1375.010 32.540 1375.330 32.600 ;
        RECT 835.430 32.400 1375.330 32.540 ;
        RECT 835.430 32.340 835.750 32.400 ;
        RECT 1375.010 32.340 1375.330 32.400 ;
      LAYER via ;
        RECT 835.460 32.340 835.720 32.600 ;
        RECT 1375.040 32.340 1375.300 32.600 ;
      LAYER met2 ;
        RECT 1375.950 1700.410 1376.230 1704.000 ;
        RECT 1375.100 1700.270 1376.230 1700.410 ;
        RECT 1375.100 32.630 1375.240 1700.270 ;
        RECT 1375.950 1700.000 1376.230 1700.270 ;
        RECT 835.460 32.310 835.720 32.630 ;
        RECT 1375.040 32.310 1375.300 32.630 ;
        RECT 835.520 2.400 835.660 32.310 ;
        RECT 835.310 -4.800 835.870 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1903.090 40.020 1903.410 40.080 ;
        RECT 2779.850 40.020 2780.170 40.080 ;
        RECT 1903.090 39.880 2780.170 40.020 ;
        RECT 1903.090 39.820 1903.410 39.880 ;
        RECT 2779.850 39.820 2780.170 39.880 ;
      LAYER via ;
        RECT 1903.120 39.820 1903.380 40.080 ;
        RECT 2779.880 39.820 2780.140 40.080 ;
      LAYER met2 ;
        RECT 1903.570 1700.410 1903.850 1704.000 ;
        RECT 1903.180 1700.270 1903.850 1700.410 ;
        RECT 1903.180 40.110 1903.320 1700.270 ;
        RECT 1903.570 1700.000 1903.850 1700.270 ;
        RECT 1903.120 39.790 1903.380 40.110 ;
        RECT 2779.880 39.790 2780.140 40.110 ;
        RECT 2779.940 2.400 2780.080 39.790 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 0.300 ;
=======
      LAYER met1 ;
        RECT 1909.530 39.680 1909.850 39.740 ;
        RECT 2797.790 39.680 2798.110 39.740 ;
        RECT 1909.530 39.540 2798.110 39.680 ;
        RECT 1909.530 39.480 1909.850 39.540 ;
        RECT 2797.790 39.480 2798.110 39.540 ;
      LAYER via ;
        RECT 1909.560 39.480 1909.820 39.740 ;
        RECT 2797.820 39.480 2798.080 39.740 ;
      LAYER met2 ;
        RECT 1908.170 1700.410 1908.450 1704.000 ;
        RECT 1908.170 1700.270 1909.760 1700.410 ;
        RECT 1908.170 1700.000 1908.450 1700.270 ;
        RECT 1909.620 39.770 1909.760 1700.270 ;
        RECT 1909.560 39.450 1909.820 39.770 ;
        RECT 2797.820 39.450 2798.080 39.770 ;
        RECT 2797.880 2.400 2798.020 39.450 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1913.210 1683.920 1913.530 1683.980 ;
        RECT 1916.430 1683.920 1916.750 1683.980 ;
        RECT 1913.210 1683.780 1916.750 1683.920 ;
        RECT 1913.210 1683.720 1913.530 1683.780 ;
        RECT 1916.430 1683.720 1916.750 1683.780 ;
        RECT 1916.430 39.340 1916.750 39.400 ;
        RECT 2815.730 39.340 2816.050 39.400 ;
        RECT 1916.430 39.200 2816.050 39.340 ;
        RECT 1916.430 39.140 1916.750 39.200 ;
        RECT 2815.730 39.140 2816.050 39.200 ;
      LAYER via ;
        RECT 1913.240 1683.720 1913.500 1683.980 ;
        RECT 1916.460 1683.720 1916.720 1683.980 ;
        RECT 1916.460 39.140 1916.720 39.400 ;
        RECT 2815.760 39.140 2816.020 39.400 ;
      LAYER met2 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2815.610 -4.800 2816.170 0.300 ;
=======
        RECT 1910.010 1700.000 1910.290 1704.000 ;
        RECT 1910.080 41.325 1910.220 1700.000 ;
        RECT 1910.010 40.955 1910.290 41.325 ;
        RECT 2815.750 40.955 2816.030 41.325 ;
        RECT 2815.820 2.400 2815.960 40.955 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
      LAYER via2 ;
        RECT 1910.010 41.000 1910.290 41.280 ;
        RECT 2815.750 41.000 2816.030 41.280 ;
      LAYER met3 ;
        RECT 1909.985 41.290 1910.315 41.305 ;
        RECT 2815.725 41.290 2816.055 41.305 ;
        RECT 1909.985 40.990 2816.055 41.290 ;
        RECT 1909.985 40.975 1910.315 40.990 ;
        RECT 2815.725 40.975 2816.055 40.990 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1913.230 1700.000 1913.510 1704.000 ;
        RECT 1913.300 1684.010 1913.440 1700.000 ;
        RECT 1913.240 1683.690 1913.500 1684.010 ;
        RECT 1916.460 1683.690 1916.720 1684.010 ;
        RECT 1916.520 39.430 1916.660 1683.690 ;
        RECT 1916.460 39.110 1916.720 39.430 ;
        RECT 2815.760 39.110 2816.020 39.430 ;
        RECT 2815.820 2.400 2815.960 39.110 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1915.970 1684.260 1916.290 1684.320 ;
        RECT 1917.810 1684.260 1918.130 1684.320 ;
        RECT 1915.970 1684.120 1918.130 1684.260 ;
        RECT 1915.970 1684.060 1916.290 1684.120 ;
        RECT 1917.810 1684.060 1918.130 1684.120 ;
        RECT 1915.970 39.000 1916.290 39.060 ;
        RECT 2833.670 39.000 2833.990 39.060 ;
        RECT 1915.970 38.860 2833.990 39.000 ;
        RECT 1915.970 38.800 1916.290 38.860 ;
        RECT 2833.670 38.800 2833.990 38.860 ;
      LAYER via ;
        RECT 1916.000 1684.060 1916.260 1684.320 ;
        RECT 1917.840 1684.060 1918.100 1684.320 ;
        RECT 1916.000 38.800 1916.260 39.060 ;
        RECT 2833.700 38.800 2833.960 39.060 ;
      LAYER met2 ;
        RECT 1917.830 1700.000 1918.110 1704.000 ;
        RECT 1917.900 1684.350 1918.040 1700.000 ;
        RECT 1916.000 1684.030 1916.260 1684.350 ;
        RECT 1917.840 1684.030 1918.100 1684.350 ;
        RECT 1916.060 39.090 1916.200 1684.030 ;
        RECT 1916.000 38.770 1916.260 39.090 ;
        RECT 2833.700 38.770 2833.960 39.090 ;
        RECT 2833.760 2.400 2833.900 38.770 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1917.370 40.320 1917.650 40.600 ;
        RECT 2833.690 40.320 2833.970 40.600 ;
      LAYER met3 ;
        RECT 1917.345 40.610 1917.675 40.625 ;
        RECT 2833.665 40.610 2833.995 40.625 ;
        RECT 1917.345 40.310 2833.995 40.610 ;
        RECT 1917.345 40.295 1917.675 40.310 ;
        RECT 2833.665 40.295 2833.995 40.310 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1923.330 38.660 1923.650 38.720 ;
        RECT 2851.150 38.660 2851.470 38.720 ;
        RECT 1923.330 38.520 2851.470 38.660 ;
        RECT 1923.330 38.460 1923.650 38.520 ;
        RECT 2851.150 38.460 2851.470 38.520 ;
      LAYER via ;
        RECT 1923.360 38.460 1923.620 38.720 ;
        RECT 2851.180 38.460 2851.440 38.720 ;
      LAYER met2 ;
        RECT 1922.890 1700.410 1923.170 1704.000 ;
        RECT 1922.890 1700.270 1923.560 1700.410 ;
        RECT 1922.890 1700.000 1923.170 1700.270 ;
        RECT 1923.420 38.750 1923.560 1700.270 ;
        RECT 1923.360 38.430 1923.620 38.750 ;
        RECT 2851.180 38.430 2851.440 38.750 ;
        RECT 2851.240 2.400 2851.380 38.430 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1923.350 39.640 1923.630 39.920 ;
        RECT 2851.170 39.640 2851.450 39.920 ;
      LAYER met3 ;
        RECT 1923.325 39.930 1923.655 39.945 ;
        RECT 2851.145 39.930 2851.475 39.945 ;
        RECT 1923.325 39.630 2851.475 39.930 ;
        RECT 1923.325 39.615 1923.655 39.630 ;
        RECT 2851.145 39.615 2851.475 39.630 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2868.970 -4.800 2869.530 0.300 ;
=======
        RECT 1924.730 1700.410 1925.010 1704.000 ;
        RECT 1923.420 1700.270 1925.010 1700.410 ;
        RECT 1923.420 1677.970 1923.560 1700.270 ;
        RECT 1924.730 1700.000 1925.010 1700.270 ;
        RECT 1922.960 1677.830 1923.560 1677.970 ;
        RECT 1922.960 39.285 1923.100 1677.830 ;
        RECT 1922.890 38.915 1923.170 39.285 ;
        RECT 2869.110 38.915 2869.390 39.285 ;
        RECT 2869.180 2.400 2869.320 38.915 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
      LAYER via2 ;
        RECT 1922.890 38.960 1923.170 39.240 ;
        RECT 2869.110 38.960 2869.390 39.240 ;
      LAYER met3 ;
        RECT 1922.865 39.250 1923.195 39.265 ;
        RECT 2869.085 39.250 2869.415 39.265 ;
        RECT 1922.865 38.950 2869.415 39.250 ;
        RECT 1922.865 38.935 1923.195 38.950 ;
        RECT 2869.085 38.935 2869.415 38.950 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1927.470 1685.280 1927.790 1685.340 ;
        RECT 1930.230 1685.280 1930.550 1685.340 ;
        RECT 1927.470 1685.140 1930.550 1685.280 ;
        RECT 1927.470 1685.080 1927.790 1685.140 ;
        RECT 1930.230 1685.080 1930.550 1685.140 ;
        RECT 1930.230 38.320 1930.550 38.380 ;
        RECT 2869.090 38.320 2869.410 38.380 ;
        RECT 1930.230 38.180 2869.410 38.320 ;
        RECT 1930.230 38.120 1930.550 38.180 ;
        RECT 2869.090 38.120 2869.410 38.180 ;
      LAYER via ;
        RECT 1927.500 1685.080 1927.760 1685.340 ;
        RECT 1930.260 1685.080 1930.520 1685.340 ;
        RECT 1930.260 38.120 1930.520 38.380 ;
        RECT 2869.120 38.120 2869.380 38.380 ;
      LAYER met2 ;
        RECT 1927.490 1700.000 1927.770 1704.000 ;
        RECT 1927.560 1685.370 1927.700 1700.000 ;
        RECT 1927.500 1685.050 1927.760 1685.370 ;
        RECT 1930.260 1685.050 1930.520 1685.370 ;
        RECT 1930.320 38.410 1930.460 1685.050 ;
        RECT 1930.260 38.090 1930.520 38.410 ;
        RECT 2869.120 38.090 2869.380 38.410 ;
        RECT 2869.180 2.400 2869.320 38.090 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1932.530 1684.260 1932.850 1684.320 ;
        RECT 1937.130 1684.260 1937.450 1684.320 ;
        RECT 1932.530 1684.120 1937.450 1684.260 ;
        RECT 1932.530 1684.060 1932.850 1684.120 ;
        RECT 1937.130 1684.060 1937.450 1684.120 ;
        RECT 1937.130 37.980 1937.450 38.040 ;
        RECT 2887.030 37.980 2887.350 38.040 ;
        RECT 1937.130 37.840 2887.350 37.980 ;
        RECT 1937.130 37.780 1937.450 37.840 ;
        RECT 2887.030 37.780 2887.350 37.840 ;
      LAYER via ;
        RECT 1932.560 1684.060 1932.820 1684.320 ;
        RECT 1937.160 1684.060 1937.420 1684.320 ;
        RECT 1937.160 37.780 1937.420 38.040 ;
        RECT 2887.060 37.780 2887.320 38.040 ;
      LAYER met2 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 2886.910 -4.800 2887.470 0.300 ;
=======
        RECT 1929.330 1700.410 1929.610 1704.000 ;
        RECT 1929.330 1700.270 1930.920 1700.410 ;
        RECT 1929.330 1700.000 1929.610 1700.270 ;
        RECT 1930.780 38.605 1930.920 1700.270 ;
        RECT 1930.710 38.235 1930.990 38.605 ;
        RECT 2887.050 38.235 2887.330 38.605 ;
        RECT 2887.120 2.400 2887.260 38.235 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
      LAYER via2 ;
        RECT 1930.710 38.280 1930.990 38.560 ;
        RECT 2887.050 38.280 2887.330 38.560 ;
      LAYER met3 ;
        RECT 1930.685 38.570 1931.015 38.585 ;
        RECT 2887.025 38.570 2887.355 38.585 ;
        RECT 1930.685 38.270 2887.355 38.570 ;
        RECT 1930.685 38.255 1931.015 38.270 ;
        RECT 2887.025 38.255 2887.355 38.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1932.550 1700.000 1932.830 1704.000 ;
        RECT 1932.620 1684.350 1932.760 1700.000 ;
        RECT 1932.560 1684.030 1932.820 1684.350 ;
        RECT 1937.160 1684.030 1937.420 1684.350 ;
        RECT 1937.220 38.070 1937.360 1684.030 ;
        RECT 1937.160 37.750 1937.420 38.070 ;
        RECT 2887.060 37.750 2887.320 38.070 ;
        RECT 2887.120 2.400 2887.260 37.750 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1934.370 1684.260 1934.690 1684.320 ;
        RECT 1938.050 1684.260 1938.370 1684.320 ;
        RECT 1934.370 1684.120 1938.370 1684.260 ;
        RECT 1934.370 1684.060 1934.690 1684.120 ;
        RECT 1938.050 1684.060 1938.370 1684.120 ;
      LAYER via ;
        RECT 1934.400 1684.060 1934.660 1684.320 ;
        RECT 1938.080 1684.060 1938.340 1684.320 ;
=======
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1937.150 1700.410 1937.430 1704.000 ;
        RECT 1937.150 1700.270 1937.820 1700.410 ;
        RECT 1937.150 1700.000 1937.430 1700.270 ;
        RECT 1937.680 37.925 1937.820 1700.270 ;
        RECT 1937.610 37.555 1937.890 37.925 ;
        RECT 2904.990 37.555 2905.270 37.925 ;
        RECT 2905.060 2.400 2905.200 37.555 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 1937.610 37.600 1937.890 37.880 ;
        RECT 2904.990 37.600 2905.270 37.880 ;
      LAYER met3 ;
        RECT 1937.585 37.890 1937.915 37.905 ;
        RECT 2904.965 37.890 2905.295 37.905 ;
        RECT 1937.585 37.590 2905.295 37.890 ;
        RECT 1937.585 37.575 1937.915 37.590 ;
        RECT 2904.965 37.575 2905.295 37.590 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 0.300 ;
=======
      LAYER met1 ;
        RECT 852.910 32.880 853.230 32.940 ;
        RECT 1380.530 32.880 1380.850 32.940 ;
        RECT 852.910 32.740 1380.850 32.880 ;
        RECT 852.910 32.680 853.230 32.740 ;
        RECT 1380.530 32.680 1380.850 32.740 ;
      LAYER via ;
        RECT 852.940 32.680 853.200 32.940 ;
        RECT 1380.560 32.680 1380.820 32.940 ;
      LAYER met2 ;
        RECT 1381.010 1700.410 1381.290 1704.000 ;
        RECT 1380.620 1700.270 1381.290 1700.410 ;
        RECT 1380.620 32.970 1380.760 1700.270 ;
        RECT 1381.010 1700.000 1381.290 1700.270 ;
        RECT 852.940 32.650 853.200 32.970 ;
        RECT 1380.560 32.650 1380.820 32.970 ;
        RECT 853.000 2.400 853.140 32.650 ;
        RECT 852.790 -4.800 853.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1380.070 1678.480 1380.390 1678.540 ;
        RECT 1384.670 1678.480 1384.990 1678.540 ;
        RECT 1380.070 1678.340 1384.990 1678.480 ;
        RECT 1380.070 1678.280 1380.390 1678.340 ;
        RECT 1384.670 1678.280 1384.990 1678.340 ;
        RECT 870.850 33.220 871.170 33.280 ;
        RECT 1380.070 33.220 1380.390 33.280 ;
        RECT 870.850 33.080 1380.390 33.220 ;
        RECT 870.850 33.020 871.170 33.080 ;
        RECT 1380.070 33.020 1380.390 33.080 ;
      LAYER via ;
        RECT 1380.100 1678.280 1380.360 1678.540 ;
        RECT 1384.700 1678.280 1384.960 1678.540 ;
        RECT 870.880 33.020 871.140 33.280 ;
        RECT 1380.100 33.020 1380.360 33.280 ;
      LAYER met2 ;
        RECT 1385.610 1700.410 1385.890 1704.000 ;
        RECT 1384.760 1700.270 1385.890 1700.410 ;
        RECT 1384.760 1678.570 1384.900 1700.270 ;
        RECT 1385.610 1700.000 1385.890 1700.270 ;
        RECT 1380.100 1678.250 1380.360 1678.570 ;
        RECT 1384.700 1678.250 1384.960 1678.570 ;
        RECT 1380.160 33.310 1380.300 1678.250 ;
        RECT 870.880 32.990 871.140 33.310 ;
        RECT 1380.100 32.990 1380.360 33.310 ;
        RECT 870.940 2.400 871.080 32.990 ;
        RECT 870.730 -4.800 871.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 0.300 ;
=======
      LAYER met1 ;
        RECT 888.790 33.220 889.110 33.280 ;
        RECT 1388.810 33.220 1389.130 33.280 ;
        RECT 888.790 33.080 1389.130 33.220 ;
        RECT 888.790 33.020 889.110 33.080 ;
        RECT 1388.810 33.020 1389.130 33.080 ;
      LAYER via ;
        RECT 888.820 33.020 889.080 33.280 ;
        RECT 1388.840 33.020 1389.100 33.280 ;
      LAYER met2 ;
        RECT 1389.750 1700.410 1390.030 1704.000 ;
        RECT 1388.900 1700.270 1390.030 1700.410 ;
        RECT 1388.900 33.310 1389.040 1700.270 ;
        RECT 1389.750 1700.000 1390.030 1700.270 ;
        RECT 888.820 32.990 889.080 33.310 ;
        RECT 1388.840 32.990 1389.100 33.310 ;
        RECT 888.880 2.400 889.020 32.990 ;
        RECT 888.670 -4.800 889.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1388.425 1442.025 1388.595 1506.115 ;
        RECT 1388.885 1228.165 1389.055 1235.475 ;
        RECT 1387.965 952.085 1388.135 986.595 ;
        RECT 1388.425 476.085 1388.595 524.195 ;
        RECT 1388.885 434.945 1389.055 449.055 ;
        RECT 1388.425 331.245 1388.595 379.355 ;
      LAYER mcon ;
        RECT 1388.425 1505.945 1388.595 1506.115 ;
        RECT 1388.885 1235.305 1389.055 1235.475 ;
        RECT 1387.965 986.425 1388.135 986.595 ;
        RECT 1388.425 524.025 1388.595 524.195 ;
        RECT 1388.885 448.885 1389.055 449.055 ;
        RECT 1388.425 379.185 1388.595 379.355 ;
      LAYER met1 ;
        RECT 1388.350 1607.900 1388.670 1608.160 ;
        RECT 1388.440 1607.420 1388.580 1607.900 ;
        RECT 1388.810 1607.420 1389.130 1607.480 ;
        RECT 1388.440 1607.280 1389.130 1607.420 ;
        RECT 1388.810 1607.220 1389.130 1607.280 ;
        RECT 1388.365 1506.100 1388.655 1506.145 ;
        RECT 1388.810 1506.100 1389.130 1506.160 ;
        RECT 1388.365 1505.960 1389.130 1506.100 ;
        RECT 1388.365 1505.915 1388.655 1505.960 ;
        RECT 1388.810 1505.900 1389.130 1505.960 ;
        RECT 1388.350 1442.180 1388.670 1442.240 ;
        RECT 1388.155 1442.040 1388.670 1442.180 ;
        RECT 1388.350 1441.980 1388.670 1442.040 ;
        RECT 1388.350 1352.760 1388.670 1352.820 ;
        RECT 1388.810 1352.760 1389.130 1352.820 ;
        RECT 1388.350 1352.620 1389.130 1352.760 ;
        RECT 1388.350 1352.560 1388.670 1352.620 ;
        RECT 1388.810 1352.560 1389.130 1352.620 ;
        RECT 1388.810 1235.460 1389.130 1235.520 ;
        RECT 1388.615 1235.320 1389.130 1235.460 ;
        RECT 1388.810 1235.260 1389.130 1235.320 ;
        RECT 1388.810 1228.320 1389.130 1228.380 ;
        RECT 1388.615 1228.180 1389.130 1228.320 ;
        RECT 1388.810 1228.120 1389.130 1228.180 ;
        RECT 1388.810 1179.700 1389.130 1179.760 ;
        RECT 1389.270 1179.700 1389.590 1179.760 ;
        RECT 1388.810 1179.560 1389.590 1179.700 ;
        RECT 1388.810 1179.500 1389.130 1179.560 ;
        RECT 1389.270 1179.500 1389.590 1179.560 ;
        RECT 1387.905 986.580 1388.195 986.625 ;
        RECT 1388.350 986.580 1388.670 986.640 ;
        RECT 1387.905 986.440 1388.670 986.580 ;
        RECT 1387.905 986.395 1388.195 986.440 ;
        RECT 1388.350 986.380 1388.670 986.440 ;
        RECT 1387.905 952.240 1388.195 952.285 ;
        RECT 1388.350 952.240 1388.670 952.300 ;
        RECT 1387.905 952.100 1388.670 952.240 ;
        RECT 1387.905 952.055 1388.195 952.100 ;
        RECT 1388.350 952.040 1388.670 952.100 ;
        RECT 1388.350 926.740 1388.670 926.800 ;
        RECT 1389.730 926.740 1390.050 926.800 ;
        RECT 1388.350 926.600 1390.050 926.740 ;
        RECT 1388.350 926.540 1388.670 926.600 ;
        RECT 1389.730 926.540 1390.050 926.600 ;
        RECT 1386.970 758.440 1387.290 758.500 ;
        RECT 1388.810 758.440 1389.130 758.500 ;
        RECT 1386.970 758.300 1389.130 758.440 ;
        RECT 1386.970 758.240 1387.290 758.300 ;
        RECT 1388.810 758.240 1389.130 758.300 ;
        RECT 1386.970 704.040 1387.290 704.100 ;
        RECT 1388.350 704.040 1388.670 704.100 ;
        RECT 1386.970 703.900 1388.670 704.040 ;
        RECT 1386.970 703.840 1387.290 703.900 ;
        RECT 1388.350 703.840 1388.670 703.900 ;
        RECT 1388.350 524.180 1388.670 524.240 ;
        RECT 1388.155 524.040 1388.670 524.180 ;
        RECT 1388.350 523.980 1388.670 524.040 ;
        RECT 1388.365 476.240 1388.655 476.285 ;
        RECT 1388.810 476.240 1389.130 476.300 ;
        RECT 1388.365 476.100 1389.130 476.240 ;
        RECT 1388.365 476.055 1388.655 476.100 ;
        RECT 1388.810 476.040 1389.130 476.100 ;
        RECT 1388.810 449.040 1389.130 449.100 ;
        RECT 1388.615 448.900 1389.130 449.040 ;
        RECT 1388.810 448.840 1389.130 448.900 ;
        RECT 1388.810 435.100 1389.130 435.160 ;
        RECT 1388.615 434.960 1389.130 435.100 ;
        RECT 1388.810 434.900 1389.130 434.960 ;
        RECT 1388.365 379.340 1388.655 379.385 ;
        RECT 1388.810 379.340 1389.130 379.400 ;
        RECT 1388.365 379.200 1389.130 379.340 ;
        RECT 1388.365 379.155 1388.655 379.200 ;
        RECT 1388.810 379.140 1389.130 379.200 ;
        RECT 1388.350 331.400 1388.670 331.460 ;
        RECT 1388.155 331.260 1388.670 331.400 ;
        RECT 1388.350 331.200 1388.670 331.260 ;
        RECT 1388.350 303.660 1388.670 303.920 ;
        RECT 1388.440 303.520 1388.580 303.660 ;
        RECT 1388.810 303.520 1389.130 303.580 ;
        RECT 1388.440 303.380 1389.130 303.520 ;
        RECT 1388.810 303.320 1389.130 303.380 ;
        RECT 1388.810 255.580 1389.130 255.640 ;
        RECT 1388.440 255.440 1389.130 255.580 ;
        RECT 1388.440 255.300 1388.580 255.440 ;
        RECT 1388.810 255.380 1389.130 255.440 ;
        RECT 1388.350 255.040 1388.670 255.300 ;
        RECT 1388.350 193.500 1388.670 193.760 ;
        RECT 1388.440 193.080 1388.580 193.500 ;
        RECT 1388.350 192.820 1388.670 193.080 ;
        RECT 888.790 33.560 889.110 33.620 ;
        RECT 1388.810 33.560 1389.130 33.620 ;
        RECT 888.790 33.420 1389.130 33.560 ;
        RECT 888.790 33.360 889.110 33.420 ;
        RECT 1388.810 33.360 1389.130 33.420 ;
      LAYER via ;
        RECT 1388.380 1607.900 1388.640 1608.160 ;
        RECT 1388.840 1607.220 1389.100 1607.480 ;
        RECT 1388.840 1505.900 1389.100 1506.160 ;
        RECT 1388.380 1441.980 1388.640 1442.240 ;
        RECT 1388.380 1352.560 1388.640 1352.820 ;
        RECT 1388.840 1352.560 1389.100 1352.820 ;
        RECT 1388.840 1235.260 1389.100 1235.520 ;
        RECT 1388.840 1228.120 1389.100 1228.380 ;
        RECT 1388.840 1179.500 1389.100 1179.760 ;
        RECT 1389.300 1179.500 1389.560 1179.760 ;
        RECT 1388.380 986.380 1388.640 986.640 ;
        RECT 1388.380 952.040 1388.640 952.300 ;
        RECT 1388.380 926.540 1388.640 926.800 ;
        RECT 1389.760 926.540 1390.020 926.800 ;
        RECT 1387.000 758.240 1387.260 758.500 ;
        RECT 1388.840 758.240 1389.100 758.500 ;
        RECT 1387.000 703.840 1387.260 704.100 ;
        RECT 1388.380 703.840 1388.640 704.100 ;
        RECT 1388.380 523.980 1388.640 524.240 ;
        RECT 1388.840 476.040 1389.100 476.300 ;
        RECT 1388.840 448.840 1389.100 449.100 ;
        RECT 1388.840 434.900 1389.100 435.160 ;
        RECT 1388.840 379.140 1389.100 379.400 ;
        RECT 1388.380 331.200 1388.640 331.460 ;
        RECT 1388.380 303.660 1388.640 303.920 ;
        RECT 1388.840 303.320 1389.100 303.580 ;
        RECT 1388.840 255.380 1389.100 255.640 ;
        RECT 1388.380 255.040 1388.640 255.300 ;
        RECT 1388.380 193.500 1388.640 193.760 ;
        RECT 1388.380 192.820 1388.640 193.080 ;
        RECT 888.820 33.360 889.080 33.620 ;
        RECT 1388.840 33.360 1389.100 33.620 ;
      LAYER met2 ;
        RECT 1390.670 1700.410 1390.950 1704.000 ;
        RECT 1389.360 1700.270 1390.950 1700.410 ;
        RECT 1389.360 1678.140 1389.500 1700.270 ;
        RECT 1390.670 1700.000 1390.950 1700.270 ;
        RECT 1388.440 1678.000 1389.500 1678.140 ;
        RECT 1388.440 1608.190 1388.580 1678.000 ;
        RECT 1388.380 1607.870 1388.640 1608.190 ;
        RECT 1388.840 1607.190 1389.100 1607.510 ;
        RECT 1388.900 1573.365 1389.040 1607.190 ;
        RECT 1388.830 1572.995 1389.110 1573.365 ;
        RECT 1389.750 1572.995 1390.030 1573.365 ;
        RECT 1389.820 1525.085 1389.960 1572.995 ;
        RECT 1388.830 1524.715 1389.110 1525.085 ;
        RECT 1389.750 1524.715 1390.030 1525.085 ;
        RECT 1388.900 1506.190 1389.040 1524.715 ;
        RECT 1388.840 1505.870 1389.100 1506.190 ;
        RECT 1388.380 1441.950 1388.640 1442.270 ;
        RECT 1388.440 1352.850 1388.580 1441.950 ;
        RECT 1388.380 1352.530 1388.640 1352.850 ;
        RECT 1388.840 1352.530 1389.100 1352.850 ;
        RECT 1388.900 1235.550 1389.040 1352.530 ;
        RECT 1388.840 1235.230 1389.100 1235.550 ;
        RECT 1388.840 1228.090 1389.100 1228.410 ;
        RECT 1388.900 1179.790 1389.040 1228.090 ;
        RECT 1388.840 1179.470 1389.100 1179.790 ;
        RECT 1389.300 1179.470 1389.560 1179.790 ;
        RECT 1389.360 1072.770 1389.500 1179.470 ;
        RECT 1388.900 1072.630 1389.500 1072.770 ;
        RECT 1388.900 1017.690 1389.040 1072.630 ;
        RECT 1388.440 1017.550 1389.040 1017.690 ;
        RECT 1388.440 986.670 1388.580 1017.550 ;
        RECT 1388.380 986.350 1388.640 986.670 ;
        RECT 1388.380 952.010 1388.640 952.330 ;
        RECT 1388.440 926.830 1388.580 952.010 ;
        RECT 1388.380 926.510 1388.640 926.830 ;
        RECT 1389.760 926.510 1390.020 926.830 ;
        RECT 1389.820 808.365 1389.960 926.510 ;
        RECT 1389.750 807.995 1390.030 808.365 ;
        RECT 1388.370 807.315 1388.650 807.685 ;
        RECT 1388.440 759.290 1388.580 807.315 ;
        RECT 1388.440 759.150 1389.040 759.290 ;
        RECT 1388.900 758.530 1389.040 759.150 ;
        RECT 1387.000 758.210 1387.260 758.530 ;
        RECT 1388.840 758.210 1389.100 758.530 ;
        RECT 1387.060 704.130 1387.200 758.210 ;
        RECT 1387.000 703.810 1387.260 704.130 ;
        RECT 1388.380 703.810 1388.640 704.130 ;
        RECT 1388.440 703.530 1388.580 703.810 ;
        RECT 1388.440 703.390 1389.500 703.530 ;
        RECT 1389.360 689.930 1389.500 703.390 ;
        RECT 1388.900 689.790 1389.500 689.930 ;
        RECT 1388.900 643.010 1389.040 689.790 ;
        RECT 1388.900 642.870 1389.500 643.010 ;
        RECT 1389.360 641.650 1389.500 642.870 ;
        RECT 1388.900 641.510 1389.500 641.650 ;
        RECT 1388.900 572.970 1389.040 641.510 ;
        RECT 1388.440 572.830 1389.040 572.970 ;
        RECT 1388.440 524.270 1388.580 572.830 ;
        RECT 1388.380 523.950 1388.640 524.270 ;
        RECT 1388.840 476.010 1389.100 476.330 ;
        RECT 1388.900 449.130 1389.040 476.010 ;
        RECT 1388.840 448.810 1389.100 449.130 ;
        RECT 1388.840 434.870 1389.100 435.190 ;
        RECT 1388.900 381.210 1389.040 434.870 ;
        RECT 1388.440 381.070 1389.040 381.210 ;
        RECT 1388.440 379.850 1388.580 381.070 ;
        RECT 1388.440 379.710 1389.040 379.850 ;
        RECT 1388.900 379.430 1389.040 379.710 ;
        RECT 1388.840 379.110 1389.100 379.430 ;
        RECT 1388.380 331.170 1388.640 331.490 ;
        RECT 1388.440 303.950 1388.580 331.170 ;
        RECT 1388.380 303.630 1388.640 303.950 ;
        RECT 1388.840 303.290 1389.100 303.610 ;
        RECT 1388.900 255.670 1389.040 303.290 ;
        RECT 1388.840 255.350 1389.100 255.670 ;
        RECT 1388.380 255.010 1388.640 255.330 ;
        RECT 1388.440 193.790 1388.580 255.010 ;
        RECT 1388.380 193.470 1388.640 193.790 ;
        RECT 1388.380 192.790 1388.640 193.110 ;
        RECT 1388.440 144.685 1388.580 192.790 ;
        RECT 1388.370 144.315 1388.650 144.685 ;
        RECT 1388.830 143.635 1389.110 144.005 ;
        RECT 1388.900 33.650 1389.040 143.635 ;
        RECT 888.820 33.330 889.080 33.650 ;
        RECT 1388.840 33.330 1389.100 33.650 ;
        RECT 888.880 2.400 889.020 33.330 ;
        RECT 888.670 -4.800 889.230 2.400 ;
      LAYER via2 ;
        RECT 1388.830 1573.040 1389.110 1573.320 ;
        RECT 1389.750 1573.040 1390.030 1573.320 ;
        RECT 1388.830 1524.760 1389.110 1525.040 ;
        RECT 1389.750 1524.760 1390.030 1525.040 ;
        RECT 1389.750 808.040 1390.030 808.320 ;
        RECT 1388.370 807.360 1388.650 807.640 ;
        RECT 1388.370 144.360 1388.650 144.640 ;
        RECT 1388.830 143.680 1389.110 143.960 ;
      LAYER met3 ;
        RECT 1388.805 1573.330 1389.135 1573.345 ;
        RECT 1389.725 1573.330 1390.055 1573.345 ;
        RECT 1388.805 1573.030 1390.055 1573.330 ;
        RECT 1388.805 1573.015 1389.135 1573.030 ;
        RECT 1389.725 1573.015 1390.055 1573.030 ;
        RECT 1388.805 1525.050 1389.135 1525.065 ;
        RECT 1389.725 1525.050 1390.055 1525.065 ;
        RECT 1388.805 1524.750 1390.055 1525.050 ;
        RECT 1388.805 1524.735 1389.135 1524.750 ;
        RECT 1389.725 1524.735 1390.055 1524.750 ;
        RECT 1389.725 808.330 1390.055 808.345 ;
        RECT 1387.670 808.030 1390.055 808.330 ;
        RECT 1387.670 807.650 1387.970 808.030 ;
        RECT 1389.725 808.015 1390.055 808.030 ;
        RECT 1388.345 807.650 1388.675 807.665 ;
        RECT 1387.670 807.350 1388.675 807.650 ;
        RECT 1388.345 807.335 1388.675 807.350 ;
        RECT 1388.345 144.650 1388.675 144.665 ;
        RECT 1387.670 144.350 1388.675 144.650 ;
        RECT 1387.670 143.970 1387.970 144.350 ;
        RECT 1388.345 144.335 1388.675 144.350 ;
        RECT 1388.805 143.970 1389.135 143.985 ;
        RECT 1387.670 143.670 1389.135 143.970 ;
        RECT 1388.805 143.655 1389.135 143.670 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 0.300 ;
=======
      LAYER met1 ;
        RECT 906.730 33.900 907.050 33.960 ;
        RECT 1394.330 33.900 1394.650 33.960 ;
        RECT 906.730 33.760 1394.650 33.900 ;
        RECT 906.730 33.700 907.050 33.760 ;
        RECT 1394.330 33.700 1394.650 33.760 ;
      LAYER via ;
        RECT 906.760 33.700 907.020 33.960 ;
        RECT 1394.360 33.700 1394.620 33.960 ;
      LAYER met2 ;
        RECT 1395.270 1700.410 1395.550 1704.000 ;
        RECT 1394.420 1700.270 1395.550 1700.410 ;
        RECT 1394.420 33.990 1394.560 1700.270 ;
        RECT 1395.270 1700.000 1395.550 1700.270 ;
        RECT 906.760 33.670 907.020 33.990 ;
        RECT 1394.360 33.670 1394.620 33.990 ;
        RECT 906.820 2.400 906.960 33.670 ;
        RECT 906.610 -4.800 907.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1395.710 1677.460 1396.030 1677.520 ;
        RECT 1398.930 1677.460 1399.250 1677.520 ;
        RECT 1395.710 1677.320 1399.250 1677.460 ;
        RECT 1395.710 1677.260 1396.030 1677.320 ;
        RECT 1398.930 1677.260 1399.250 1677.320 ;
        RECT 924.210 34.240 924.530 34.300 ;
        RECT 1395.710 34.240 1396.030 34.300 ;
        RECT 924.210 34.100 1396.030 34.240 ;
        RECT 924.210 34.040 924.530 34.100 ;
        RECT 1395.710 34.040 1396.030 34.100 ;
      LAYER via ;
        RECT 1395.740 1677.260 1396.000 1677.520 ;
        RECT 1398.960 1677.260 1399.220 1677.520 ;
        RECT 924.240 34.040 924.500 34.300 ;
        RECT 1395.740 34.040 1396.000 34.300 ;
      LAYER met2 ;
        RECT 1400.330 1700.410 1400.610 1704.000 ;
        RECT 1399.020 1700.270 1400.610 1700.410 ;
        RECT 1399.020 1677.550 1399.160 1700.270 ;
        RECT 1400.330 1700.000 1400.610 1700.270 ;
        RECT 1395.740 1677.230 1396.000 1677.550 ;
        RECT 1398.960 1677.230 1399.220 1677.550 ;
        RECT 1395.800 34.330 1395.940 1677.230 ;
        RECT 924.240 34.010 924.500 34.330 ;
        RECT 1395.740 34.010 1396.000 34.330 ;
        RECT 924.300 2.400 924.440 34.010 ;
        RECT 924.090 -4.800 924.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1401.230 1678.820 1401.550 1678.880 ;
        RECT 1403.990 1678.820 1404.310 1678.880 ;
        RECT 1401.230 1678.680 1404.310 1678.820 ;
        RECT 1401.230 1678.620 1401.550 1678.680 ;
        RECT 1403.990 1678.620 1404.310 1678.680 ;
        RECT 942.150 30.500 942.470 30.560 ;
        RECT 1401.230 30.500 1401.550 30.560 ;
        RECT 942.150 30.360 1401.550 30.500 ;
        RECT 942.150 30.300 942.470 30.360 ;
        RECT 1401.230 30.300 1401.550 30.360 ;
      LAYER via ;
        RECT 1401.260 1678.620 1401.520 1678.880 ;
        RECT 1404.020 1678.620 1404.280 1678.880 ;
        RECT 942.180 30.300 942.440 30.560 ;
        RECT 1401.260 30.300 1401.520 30.560 ;
      LAYER met2 ;
        RECT 1404.930 1700.410 1405.210 1704.000 ;
        RECT 1404.080 1700.270 1405.210 1700.410 ;
        RECT 1404.080 1678.910 1404.220 1700.270 ;
        RECT 1404.930 1700.000 1405.210 1700.270 ;
        RECT 1401.260 1678.590 1401.520 1678.910 ;
        RECT 1404.020 1678.590 1404.280 1678.910 ;
        RECT 1401.320 30.590 1401.460 1678.590 ;
        RECT 942.180 30.270 942.440 30.590 ;
        RECT 1401.260 30.270 1401.520 30.590 ;
        RECT 942.240 2.400 942.380 30.270 ;
        RECT 942.030 -4.800 942.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 0.300 ;
=======
      LAYER met1 ;
        RECT 960.090 30.160 960.410 30.220 ;
        RECT 1408.590 30.160 1408.910 30.220 ;
        RECT 960.090 30.020 1408.910 30.160 ;
        RECT 960.090 29.960 960.410 30.020 ;
        RECT 1408.590 29.960 1408.910 30.020 ;
      LAYER via ;
        RECT 960.120 29.960 960.380 30.220 ;
        RECT 1408.620 29.960 1408.880 30.220 ;
      LAYER met2 ;
        RECT 1409.990 1700.410 1410.270 1704.000 ;
        RECT 1408.680 1700.270 1410.270 1700.410 ;
        RECT 1408.680 30.250 1408.820 1700.270 ;
        RECT 1409.990 1700.000 1410.270 1700.270 ;
        RECT 960.120 29.930 960.380 30.250 ;
        RECT 1408.620 29.930 1408.880 30.250 ;
        RECT 960.180 2.400 960.320 29.930 ;
        RECT 959.970 -4.800 960.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 0.300 ;
=======
      LAYER met1 ;
        RECT 978.030 29.820 978.350 29.880 ;
        RECT 1415.490 29.820 1415.810 29.880 ;
        RECT 978.030 29.680 1415.810 29.820 ;
        RECT 978.030 29.620 978.350 29.680 ;
        RECT 1415.490 29.620 1415.810 29.680 ;
      LAYER via ;
        RECT 978.060 29.620 978.320 29.880 ;
        RECT 1415.520 29.620 1415.780 29.880 ;
      LAYER met2 ;
        RECT 1414.590 1700.410 1414.870 1704.000 ;
        RECT 1414.590 1700.270 1415.720 1700.410 ;
        RECT 1414.590 1700.000 1414.870 1700.270 ;
        RECT 1415.580 29.910 1415.720 1700.270 ;
        RECT 978.060 29.590 978.320 29.910 ;
        RECT 1415.520 29.590 1415.780 29.910 ;
        RECT 978.120 2.400 978.260 29.590 ;
        RECT 977.910 -4.800 978.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 656.830 -4.800 657.390 0.300 ;
=======
        RECT 1327.190 1700.410 1327.470 1704.000 ;
        RECT 1325.880 1700.270 1327.470 1700.410 ;
        RECT 1325.880 33.845 1326.020 1700.270 ;
        RECT 1327.190 1700.000 1327.470 1700.270 ;
        RECT 656.970 33.475 657.250 33.845 ;
        RECT 1325.810 33.475 1326.090 33.845 ;
        RECT 657.040 2.400 657.180 33.475 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 656.970 33.520 657.250 33.800 ;
        RECT 1325.810 33.520 1326.090 33.800 ;
      LAYER met3 ;
        RECT 656.945 33.810 657.275 33.825 ;
        RECT 1325.785 33.810 1326.115 33.825 ;
        RECT 656.945 33.510 1326.115 33.810 ;
        RECT 656.945 33.495 657.275 33.510 ;
        RECT 1325.785 33.495 1326.115 33.510 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 656.950 31.860 657.270 31.920 ;
        RECT 1325.790 31.860 1326.110 31.920 ;
        RECT 656.950 31.720 1326.110 31.860 ;
        RECT 656.950 31.660 657.270 31.720 ;
        RECT 1325.790 31.660 1326.110 31.720 ;
      LAYER via ;
        RECT 656.980 31.660 657.240 31.920 ;
        RECT 1325.820 31.660 1326.080 31.920 ;
      LAYER met2 ;
        RECT 1327.650 1700.410 1327.930 1704.000 ;
        RECT 1326.800 1700.270 1327.930 1700.410 ;
        RECT 1326.800 1677.970 1326.940 1700.270 ;
        RECT 1327.650 1700.000 1327.930 1700.270 ;
        RECT 1325.880 1677.830 1326.940 1677.970 ;
        RECT 1325.880 31.950 1326.020 1677.830 ;
        RECT 656.980 31.630 657.240 31.950 ;
        RECT 1325.820 31.630 1326.080 31.950 ;
        RECT 657.040 2.400 657.180 31.630 ;
        RECT 656.830 -4.800 657.390 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1415.030 1678.140 1415.350 1678.200 ;
        RECT 1418.710 1678.140 1419.030 1678.200 ;
        RECT 1415.030 1678.000 1419.030 1678.140 ;
        RECT 1415.030 1677.940 1415.350 1678.000 ;
        RECT 1418.710 1677.940 1419.030 1678.000 ;
        RECT 995.970 29.480 996.290 29.540 ;
        RECT 1415.030 29.480 1415.350 29.540 ;
        RECT 995.970 29.340 1415.350 29.480 ;
        RECT 995.970 29.280 996.290 29.340 ;
        RECT 1415.030 29.280 1415.350 29.340 ;
      LAYER via ;
        RECT 1415.060 1677.940 1415.320 1678.200 ;
        RECT 1418.740 1677.940 1419.000 1678.200 ;
        RECT 996.000 29.280 996.260 29.540 ;
        RECT 1415.060 29.280 1415.320 29.540 ;
      LAYER met2 ;
        RECT 1419.650 1700.410 1419.930 1704.000 ;
        RECT 1418.800 1700.270 1419.930 1700.410 ;
        RECT 1418.800 1678.230 1418.940 1700.270 ;
        RECT 1419.650 1700.000 1419.930 1700.270 ;
        RECT 1415.060 1677.910 1415.320 1678.230 ;
        RECT 1418.740 1677.910 1419.000 1678.230 ;
        RECT 1415.120 29.570 1415.260 1677.910 ;
        RECT 996.000 29.250 996.260 29.570 ;
        RECT 1415.060 29.250 1415.320 29.570 ;
        RECT 996.060 2.400 996.200 29.250 ;
        RECT 995.850 -4.800 996.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 0.300 ;
=======
      LAYER met1 ;
        RECT 1013.450 29.140 1013.770 29.200 ;
        RECT 1422.390 29.140 1422.710 29.200 ;
        RECT 1013.450 29.000 1422.710 29.140 ;
        RECT 1013.450 28.940 1013.770 29.000 ;
        RECT 1422.390 28.940 1422.710 29.000 ;
      LAYER via ;
        RECT 1013.480 28.940 1013.740 29.200 ;
        RECT 1422.420 28.940 1422.680 29.200 ;
      LAYER met2 ;
        RECT 1424.710 1700.410 1424.990 1704.000 ;
        RECT 1423.400 1700.270 1424.990 1700.410 ;
        RECT 1423.400 1659.610 1423.540 1700.270 ;
        RECT 1424.710 1700.000 1424.990 1700.270 ;
        RECT 1422.480 1659.470 1423.540 1659.610 ;
        RECT 1422.480 29.230 1422.620 1659.470 ;
        RECT 1013.480 28.910 1013.740 29.230 ;
        RECT 1422.420 28.910 1422.680 29.230 ;
        RECT 1013.540 2.400 1013.680 28.910 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 0.300 ;
=======
      LAYER met1 ;
        RECT 1031.390 29.140 1031.710 29.200 ;
        RECT 1429.290 29.140 1429.610 29.200 ;
        RECT 1031.390 29.000 1429.610 29.140 ;
        RECT 1031.390 28.940 1031.710 29.000 ;
        RECT 1429.290 28.940 1429.610 29.000 ;
=======
      LAYER li1 ;
        RECT 1428.905 1283.585 1429.075 1352.435 ;
        RECT 1428.905 1041.845 1429.075 1077.035 ;
        RECT 1429.365 428.145 1429.535 475.915 ;
        RECT 1427.985 372.725 1428.155 420.835 ;
      LAYER mcon ;
        RECT 1428.905 1352.265 1429.075 1352.435 ;
        RECT 1428.905 1076.865 1429.075 1077.035 ;
        RECT 1429.365 475.745 1429.535 475.915 ;
        RECT 1427.985 420.665 1428.155 420.835 ;
      LAYER met1 ;
        RECT 1428.830 1559.280 1429.150 1559.540 ;
        RECT 1428.920 1559.140 1429.060 1559.280 ;
        RECT 1429.290 1559.140 1429.610 1559.200 ;
        RECT 1428.920 1559.000 1429.610 1559.140 ;
        RECT 1429.290 1558.940 1429.610 1559.000 ;
        RECT 1428.830 1497.600 1429.150 1497.660 ;
        RECT 1429.290 1497.600 1429.610 1497.660 ;
        RECT 1428.830 1497.460 1429.610 1497.600 ;
        RECT 1428.830 1497.400 1429.150 1497.460 ;
        RECT 1429.290 1497.400 1429.610 1497.460 ;
        RECT 1428.845 1352.420 1429.135 1352.465 ;
        RECT 1429.290 1352.420 1429.610 1352.480 ;
        RECT 1428.845 1352.280 1429.610 1352.420 ;
        RECT 1428.845 1352.235 1429.135 1352.280 ;
        RECT 1429.290 1352.220 1429.610 1352.280 ;
        RECT 1428.845 1283.740 1429.135 1283.785 ;
        RECT 1429.290 1283.740 1429.610 1283.800 ;
        RECT 1428.845 1283.600 1429.610 1283.740 ;
        RECT 1428.845 1283.555 1429.135 1283.600 ;
        RECT 1429.290 1283.540 1429.610 1283.600 ;
        RECT 1428.830 1077.020 1429.150 1077.080 ;
        RECT 1428.635 1076.880 1429.150 1077.020 ;
        RECT 1428.830 1076.820 1429.150 1076.880 ;
        RECT 1428.845 1042.000 1429.135 1042.045 ;
        RECT 1429.290 1042.000 1429.610 1042.060 ;
        RECT 1428.845 1041.860 1429.610 1042.000 ;
        RECT 1428.845 1041.815 1429.135 1041.860 ;
        RECT 1429.290 1041.800 1429.610 1041.860 ;
        RECT 1428.830 966.180 1429.150 966.240 ;
        RECT 1429.290 966.180 1429.610 966.240 ;
        RECT 1428.830 966.040 1429.610 966.180 ;
        RECT 1428.830 965.980 1429.150 966.040 ;
        RECT 1429.290 965.980 1429.610 966.040 ;
        RECT 1428.830 910.760 1429.150 910.820 ;
        RECT 1429.290 910.760 1429.610 910.820 ;
        RECT 1428.830 910.620 1429.610 910.760 ;
        RECT 1428.830 910.560 1429.150 910.620 ;
        RECT 1429.290 910.560 1429.610 910.620 ;
        RECT 1429.290 856.020 1429.610 856.080 ;
        RECT 1428.920 855.880 1429.610 856.020 ;
        RECT 1428.920 855.740 1429.060 855.880 ;
        RECT 1429.290 855.820 1429.610 855.880 ;
        RECT 1428.830 855.480 1429.150 855.740 ;
        RECT 1429.290 693.500 1429.610 693.560 ;
        RECT 1430.210 693.500 1430.530 693.560 ;
        RECT 1429.290 693.360 1430.530 693.500 ;
        RECT 1429.290 693.300 1429.610 693.360 ;
        RECT 1430.210 693.300 1430.530 693.360 ;
        RECT 1429.290 475.900 1429.610 475.960 ;
        RECT 1429.095 475.760 1429.610 475.900 ;
        RECT 1429.290 475.700 1429.610 475.760 ;
        RECT 1429.290 428.300 1429.610 428.360 ;
        RECT 1429.095 428.160 1429.610 428.300 ;
        RECT 1429.290 428.100 1429.610 428.160 ;
        RECT 1427.925 420.820 1428.215 420.865 ;
        RECT 1429.290 420.820 1429.610 420.880 ;
        RECT 1427.925 420.680 1429.610 420.820 ;
        RECT 1427.925 420.635 1428.215 420.680 ;
        RECT 1429.290 420.620 1429.610 420.680 ;
        RECT 1427.925 372.880 1428.215 372.925 ;
        RECT 1428.370 372.880 1428.690 372.940 ;
        RECT 1427.925 372.740 1428.690 372.880 ;
        RECT 1427.925 372.695 1428.215 372.740 ;
        RECT 1428.370 372.680 1428.690 372.740 ;
        RECT 1428.830 203.560 1429.150 203.620 ;
        RECT 1430.210 203.560 1430.530 203.620 ;
        RECT 1428.830 203.420 1430.530 203.560 ;
        RECT 1428.830 203.360 1429.150 203.420 ;
        RECT 1430.210 203.360 1430.530 203.420 ;
        RECT 1428.370 141.680 1428.690 141.740 ;
        RECT 1430.210 141.680 1430.530 141.740 ;
        RECT 1428.370 141.540 1430.530 141.680 ;
        RECT 1428.370 141.480 1428.690 141.540 ;
        RECT 1430.210 141.480 1430.530 141.540 ;
        RECT 1428.370 83.200 1428.690 83.260 ;
        RECT 1428.830 83.200 1429.150 83.260 ;
        RECT 1428.370 83.060 1429.150 83.200 ;
        RECT 1428.370 83.000 1428.690 83.060 ;
        RECT 1428.830 83.000 1429.150 83.060 ;
        RECT 1031.390 28.800 1031.710 28.860 ;
        RECT 1428.830 28.800 1429.150 28.860 ;
        RECT 1031.390 28.660 1429.150 28.800 ;
        RECT 1031.390 28.600 1031.710 28.660 ;
        RECT 1428.830 28.600 1429.150 28.660 ;
>>>>>>> re-updated local openlane
      LAYER via ;
        RECT 1428.860 1559.280 1429.120 1559.540 ;
        RECT 1429.320 1558.940 1429.580 1559.200 ;
        RECT 1428.860 1497.400 1429.120 1497.660 ;
        RECT 1429.320 1497.400 1429.580 1497.660 ;
        RECT 1429.320 1352.220 1429.580 1352.480 ;
        RECT 1429.320 1283.540 1429.580 1283.800 ;
        RECT 1428.860 1076.820 1429.120 1077.080 ;
        RECT 1429.320 1041.800 1429.580 1042.060 ;
        RECT 1428.860 965.980 1429.120 966.240 ;
        RECT 1429.320 965.980 1429.580 966.240 ;
        RECT 1428.860 910.560 1429.120 910.820 ;
        RECT 1429.320 910.560 1429.580 910.820 ;
        RECT 1429.320 855.820 1429.580 856.080 ;
        RECT 1428.860 855.480 1429.120 855.740 ;
        RECT 1429.320 693.300 1429.580 693.560 ;
        RECT 1430.240 693.300 1430.500 693.560 ;
        RECT 1429.320 475.700 1429.580 475.960 ;
        RECT 1429.320 428.100 1429.580 428.360 ;
        RECT 1429.320 420.620 1429.580 420.880 ;
        RECT 1428.400 372.680 1428.660 372.940 ;
        RECT 1428.860 203.360 1429.120 203.620 ;
        RECT 1430.240 203.360 1430.500 203.620 ;
        RECT 1428.400 141.480 1428.660 141.740 ;
        RECT 1430.240 141.480 1430.500 141.740 ;
        RECT 1428.400 83.000 1428.660 83.260 ;
        RECT 1428.860 83.000 1429.120 83.260 ;
        RECT 1031.420 28.600 1031.680 28.860 ;
        RECT 1428.860 28.600 1429.120 28.860 ;
      LAYER met2 ;
        RECT 1429.310 1700.000 1429.590 1704.000 ;
        RECT 1429.380 1618.130 1429.520 1700.000 ;
        RECT 1428.920 1617.990 1429.520 1618.130 ;
        RECT 1428.920 1559.570 1429.060 1617.990 ;
        RECT 1428.860 1559.250 1429.120 1559.570 ;
        RECT 1429.320 1558.910 1429.580 1559.230 ;
        RECT 1429.380 1497.690 1429.520 1558.910 ;
        RECT 1428.860 1497.370 1429.120 1497.690 ;
        RECT 1429.320 1497.370 1429.580 1497.690 ;
        RECT 1428.920 1460.370 1429.060 1497.370 ;
        RECT 1428.920 1460.230 1429.520 1460.370 ;
        RECT 1429.380 1352.510 1429.520 1460.230 ;
        RECT 1429.320 1352.190 1429.580 1352.510 ;
        RECT 1429.320 1283.510 1429.580 1283.830 ;
        RECT 1429.380 1208.090 1429.520 1283.510 ;
        RECT 1428.920 1207.950 1429.520 1208.090 ;
        RECT 1428.920 1077.110 1429.060 1207.950 ;
        RECT 1428.860 1076.790 1429.120 1077.110 ;
        RECT 1429.320 1041.770 1429.580 1042.090 ;
        RECT 1429.380 1024.490 1429.520 1041.770 ;
        RECT 1428.920 1024.350 1429.520 1024.490 ;
        RECT 1428.920 966.270 1429.060 1024.350 ;
        RECT 1428.860 966.010 1429.120 966.270 ;
        RECT 1429.320 966.010 1429.580 966.270 ;
        RECT 1428.860 965.950 1429.580 966.010 ;
        RECT 1428.920 965.870 1429.520 965.950 ;
        RECT 1428.920 910.850 1429.060 965.870 ;
        RECT 1428.860 910.530 1429.120 910.850 ;
        RECT 1429.320 910.530 1429.580 910.850 ;
        RECT 1429.380 856.110 1429.520 910.530 ;
        RECT 1429.320 855.790 1429.580 856.110 ;
        RECT 1428.860 855.450 1429.120 855.770 ;
        RECT 1428.920 806.890 1429.060 855.450 ;
        RECT 1428.920 806.750 1429.520 806.890 ;
        RECT 1429.380 693.590 1429.520 806.750 ;
        RECT 1429.320 693.270 1429.580 693.590 ;
        RECT 1430.240 693.270 1430.500 693.590 ;
        RECT 1430.300 579.885 1430.440 693.270 ;
        RECT 1429.310 579.515 1429.590 579.885 ;
        RECT 1430.230 579.515 1430.510 579.885 ;
        RECT 1429.380 555.290 1429.520 579.515 ;
        RECT 1428.920 555.150 1429.520 555.290 ;
        RECT 1428.920 500.210 1429.060 555.150 ;
        RECT 1428.920 500.070 1429.520 500.210 ;
        RECT 1429.380 475.990 1429.520 500.070 ;
        RECT 1429.320 475.670 1429.580 475.990 ;
        RECT 1429.320 428.070 1429.580 428.390 ;
        RECT 1429.380 420.910 1429.520 428.070 ;
        RECT 1429.320 420.590 1429.580 420.910 ;
        RECT 1428.400 372.650 1428.660 372.970 ;
        RECT 1428.460 354.690 1428.600 372.650 ;
        RECT 1428.460 354.550 1429.520 354.690 ;
        RECT 1429.380 258.810 1429.520 354.550 ;
        RECT 1428.920 258.670 1429.520 258.810 ;
        RECT 1428.920 203.650 1429.060 258.670 ;
        RECT 1428.860 203.330 1429.120 203.650 ;
        RECT 1430.240 203.330 1430.500 203.650 ;
        RECT 1430.300 141.770 1430.440 203.330 ;
        RECT 1428.400 141.450 1428.660 141.770 ;
        RECT 1430.240 141.450 1430.500 141.770 ;
        RECT 1428.460 83.290 1428.600 141.450 ;
        RECT 1428.400 82.970 1428.660 83.290 ;
        RECT 1428.860 82.970 1429.120 83.290 ;
        RECT 1428.920 28.890 1429.060 82.970 ;
        RECT 1031.420 28.570 1031.680 28.890 ;
        RECT 1428.860 28.570 1429.120 28.890 ;
        RECT 1031.480 2.400 1031.620 28.570 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 1429.310 579.560 1429.590 579.840 ;
        RECT 1430.230 579.560 1430.510 579.840 ;
      LAYER met3 ;
        RECT 1429.285 579.850 1429.615 579.865 ;
        RECT 1430.205 579.850 1430.535 579.865 ;
        RECT 1429.285 579.550 1430.535 579.850 ;
        RECT 1429.285 579.535 1429.615 579.550 ;
        RECT 1430.205 579.535 1430.535 579.550 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1428.830 1678.480 1429.150 1678.540 ;
        RECT 1432.050 1678.480 1432.370 1678.540 ;
        RECT 1428.830 1678.340 1432.370 1678.480 ;
        RECT 1428.830 1678.280 1429.150 1678.340 ;
        RECT 1432.050 1678.280 1432.370 1678.340 ;
        RECT 1049.330 28.800 1049.650 28.860 ;
        RECT 1428.830 28.800 1429.150 28.860 ;
        RECT 1049.330 28.660 1429.150 28.800 ;
        RECT 1049.330 28.600 1049.650 28.660 ;
        RECT 1428.830 28.600 1429.150 28.660 ;
      LAYER via ;
        RECT 1428.860 1678.280 1429.120 1678.540 ;
        RECT 1432.080 1678.280 1432.340 1678.540 ;
        RECT 1049.360 28.600 1049.620 28.860 ;
        RECT 1428.860 28.600 1429.120 28.860 ;
      LAYER met2 ;
        RECT 1432.990 1700.410 1433.270 1704.000 ;
        RECT 1432.140 1700.270 1433.270 1700.410 ;
        RECT 1432.140 1678.570 1432.280 1700.270 ;
        RECT 1432.990 1700.000 1433.270 1700.270 ;
        RECT 1428.860 1678.250 1429.120 1678.570 ;
        RECT 1432.080 1678.250 1432.340 1678.570 ;
        RECT 1428.920 28.890 1429.060 1678.250 ;
        RECT 1049.360 28.570 1049.620 28.890 ;
        RECT 1428.860 28.570 1429.120 28.890 ;
        RECT 1049.420 2.400 1049.560 28.570 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1430.745 1531.445 1430.915 1539.435 ;
      LAYER mcon ;
        RECT 1430.745 1539.265 1430.915 1539.435 ;
      LAYER met1 ;
        RECT 1430.670 1573.420 1430.990 1573.480 ;
        RECT 1431.590 1573.420 1431.910 1573.480 ;
        RECT 1430.670 1573.280 1431.910 1573.420 ;
        RECT 1430.670 1573.220 1430.990 1573.280 ;
        RECT 1431.590 1573.220 1431.910 1573.280 ;
        RECT 1430.670 1539.420 1430.990 1539.480 ;
        RECT 1430.475 1539.280 1430.990 1539.420 ;
        RECT 1430.670 1539.220 1430.990 1539.280 ;
        RECT 1430.670 1531.600 1430.990 1531.660 ;
        RECT 1430.475 1531.460 1430.990 1531.600 ;
        RECT 1430.670 1531.400 1430.990 1531.460 ;
        RECT 1430.670 1449.320 1430.990 1449.380 ;
        RECT 1430.670 1449.180 1431.360 1449.320 ;
        RECT 1430.670 1449.120 1430.990 1449.180 ;
        RECT 1431.220 1449.040 1431.360 1449.180 ;
        RECT 1431.130 1448.780 1431.450 1449.040 ;
        RECT 1430.210 1363.100 1430.530 1363.360 ;
        RECT 1430.300 1362.680 1430.440 1363.100 ;
        RECT 1430.210 1362.420 1430.530 1362.680 ;
        RECT 1430.210 1304.480 1430.530 1304.540 ;
        RECT 1430.670 1304.480 1430.990 1304.540 ;
        RECT 1430.210 1304.340 1430.990 1304.480 ;
        RECT 1430.210 1304.280 1430.530 1304.340 ;
        RECT 1430.670 1304.280 1430.990 1304.340 ;
        RECT 1430.670 966.180 1430.990 966.240 ;
        RECT 1431.130 966.180 1431.450 966.240 ;
        RECT 1430.670 966.040 1431.450 966.180 ;
        RECT 1430.670 965.980 1430.990 966.040 ;
        RECT 1431.130 965.980 1431.450 966.040 ;
        RECT 1430.670 717.640 1430.990 717.700 ;
        RECT 1431.130 717.640 1431.450 717.700 ;
        RECT 1430.670 717.500 1431.450 717.640 ;
        RECT 1430.670 717.440 1430.990 717.500 ;
        RECT 1431.130 717.440 1431.450 717.500 ;
        RECT 1430.670 289.920 1430.990 289.980 ;
        RECT 1431.130 289.920 1431.450 289.980 ;
        RECT 1430.670 289.780 1431.450 289.920 ;
        RECT 1430.670 289.720 1430.990 289.780 ;
        RECT 1431.130 289.720 1431.450 289.780 ;
        RECT 1430.670 62.460 1430.990 62.520 ;
        RECT 1430.300 62.320 1430.990 62.460 ;
        RECT 1430.300 62.180 1430.440 62.320 ;
        RECT 1430.670 62.260 1430.990 62.320 ;
        RECT 1430.210 61.920 1430.530 62.180 ;
        RECT 1049.330 28.460 1049.650 28.520 ;
        RECT 1430.210 28.460 1430.530 28.520 ;
        RECT 1049.330 28.320 1430.530 28.460 ;
        RECT 1049.330 28.260 1049.650 28.320 ;
        RECT 1430.210 28.260 1430.530 28.320 ;
      LAYER via ;
        RECT 1430.700 1573.220 1430.960 1573.480 ;
        RECT 1431.620 1573.220 1431.880 1573.480 ;
        RECT 1430.700 1539.220 1430.960 1539.480 ;
        RECT 1430.700 1531.400 1430.960 1531.660 ;
        RECT 1430.700 1449.120 1430.960 1449.380 ;
        RECT 1431.160 1448.780 1431.420 1449.040 ;
        RECT 1430.240 1363.100 1430.500 1363.360 ;
        RECT 1430.240 1362.420 1430.500 1362.680 ;
        RECT 1430.240 1304.280 1430.500 1304.540 ;
        RECT 1430.700 1304.280 1430.960 1304.540 ;
        RECT 1430.700 965.980 1430.960 966.240 ;
        RECT 1431.160 965.980 1431.420 966.240 ;
        RECT 1430.700 717.440 1430.960 717.700 ;
        RECT 1431.160 717.440 1431.420 717.700 ;
        RECT 1430.700 289.720 1430.960 289.980 ;
        RECT 1431.160 289.720 1431.420 289.980 ;
        RECT 1430.700 62.260 1430.960 62.520 ;
        RECT 1430.240 61.920 1430.500 62.180 ;
        RECT 1049.360 28.260 1049.620 28.520 ;
        RECT 1430.240 28.260 1430.500 28.520 ;
      LAYER met2 ;
        RECT 1434.370 1700.410 1434.650 1704.000 ;
        RECT 1433.060 1700.270 1434.650 1700.410 ;
        RECT 1433.060 1669.925 1433.200 1700.270 ;
        RECT 1434.370 1700.000 1434.650 1700.270 ;
        RECT 1432.070 1669.555 1432.350 1669.925 ;
        RECT 1432.990 1669.555 1433.270 1669.925 ;
        RECT 1432.140 1627.650 1432.280 1669.555 ;
        RECT 1430.760 1627.510 1432.280 1627.650 ;
        RECT 1430.760 1621.645 1430.900 1627.510 ;
        RECT 1430.690 1621.275 1430.970 1621.645 ;
        RECT 1431.610 1621.275 1431.890 1621.645 ;
        RECT 1431.680 1573.510 1431.820 1621.275 ;
        RECT 1430.700 1573.190 1430.960 1573.510 ;
        RECT 1431.620 1573.190 1431.880 1573.510 ;
        RECT 1430.760 1539.510 1430.900 1573.190 ;
        RECT 1430.700 1539.190 1430.960 1539.510 ;
        RECT 1430.700 1531.370 1430.960 1531.690 ;
        RECT 1430.760 1507.970 1430.900 1531.370 ;
        RECT 1430.760 1507.830 1431.360 1507.970 ;
        RECT 1431.220 1483.490 1431.360 1507.830 ;
        RECT 1430.760 1483.350 1431.360 1483.490 ;
        RECT 1430.760 1449.410 1430.900 1483.350 ;
        RECT 1430.700 1449.090 1430.960 1449.410 ;
        RECT 1431.160 1448.750 1431.420 1449.070 ;
        RECT 1431.220 1387.045 1431.360 1448.750 ;
        RECT 1430.230 1386.675 1430.510 1387.045 ;
        RECT 1431.150 1386.675 1431.430 1387.045 ;
        RECT 1430.300 1363.390 1430.440 1386.675 ;
        RECT 1430.240 1363.070 1430.500 1363.390 ;
        RECT 1430.240 1362.390 1430.500 1362.710 ;
        RECT 1430.300 1304.570 1430.440 1362.390 ;
        RECT 1430.240 1304.250 1430.500 1304.570 ;
        RECT 1430.700 1304.250 1430.960 1304.570 ;
        RECT 1430.760 1303.970 1430.900 1304.250 ;
        RECT 1430.760 1303.830 1431.360 1303.970 ;
        RECT 1431.220 1173.410 1431.360 1303.830 ;
        RECT 1430.760 1173.270 1431.360 1173.410 ;
        RECT 1430.760 1152.330 1430.900 1173.270 ;
        RECT 1430.760 1152.190 1431.820 1152.330 ;
        RECT 1431.680 1080.250 1431.820 1152.190 ;
        RECT 1431.220 1080.110 1431.820 1080.250 ;
        RECT 1431.220 966.270 1431.360 1080.110 ;
        RECT 1430.700 965.950 1430.960 966.270 ;
        RECT 1431.160 965.950 1431.420 966.270 ;
        RECT 1430.760 910.930 1430.900 965.950 ;
        RECT 1430.760 910.790 1431.360 910.930 ;
        RECT 1431.220 787.170 1431.360 910.790 ;
        RECT 1430.760 787.030 1431.360 787.170 ;
        RECT 1430.760 742.290 1430.900 787.030 ;
        RECT 1430.760 742.150 1431.360 742.290 ;
        RECT 1431.220 717.730 1431.360 742.150 ;
        RECT 1430.700 717.410 1430.960 717.730 ;
        RECT 1431.160 717.410 1431.420 717.730 ;
        RECT 1430.760 641.650 1430.900 717.410 ;
        RECT 1430.760 641.510 1431.360 641.650 ;
        RECT 1431.220 497.490 1431.360 641.510 ;
        RECT 1430.760 497.350 1431.360 497.490 ;
        RECT 1430.760 448.530 1430.900 497.350 ;
        RECT 1430.760 448.390 1431.360 448.530 ;
        RECT 1431.220 290.010 1431.360 448.390 ;
        RECT 1430.700 289.690 1430.960 290.010 ;
        RECT 1431.160 289.690 1431.420 290.010 ;
        RECT 1430.760 254.730 1430.900 289.690 ;
        RECT 1430.760 254.590 1431.360 254.730 ;
        RECT 1431.220 110.570 1431.360 254.590 ;
        RECT 1430.760 110.430 1431.360 110.570 ;
        RECT 1430.760 62.550 1430.900 110.430 ;
        RECT 1430.700 62.230 1430.960 62.550 ;
        RECT 1430.240 61.890 1430.500 62.210 ;
        RECT 1430.300 28.550 1430.440 61.890 ;
        RECT 1049.360 28.230 1049.620 28.550 ;
        RECT 1430.240 28.230 1430.500 28.550 ;
        RECT 1049.420 2.400 1049.560 28.230 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
      LAYER via2 ;
        RECT 1432.070 1669.600 1432.350 1669.880 ;
        RECT 1432.990 1669.600 1433.270 1669.880 ;
        RECT 1430.690 1621.320 1430.970 1621.600 ;
        RECT 1431.610 1621.320 1431.890 1621.600 ;
        RECT 1430.230 1386.720 1430.510 1387.000 ;
        RECT 1431.150 1386.720 1431.430 1387.000 ;
      LAYER met3 ;
        RECT 1432.045 1669.890 1432.375 1669.905 ;
        RECT 1432.965 1669.890 1433.295 1669.905 ;
        RECT 1432.045 1669.590 1433.295 1669.890 ;
        RECT 1432.045 1669.575 1432.375 1669.590 ;
        RECT 1432.965 1669.575 1433.295 1669.590 ;
        RECT 1430.665 1621.610 1430.995 1621.625 ;
        RECT 1431.585 1621.610 1431.915 1621.625 ;
        RECT 1430.665 1621.310 1431.915 1621.610 ;
        RECT 1430.665 1621.295 1430.995 1621.310 ;
        RECT 1431.585 1621.295 1431.915 1621.310 ;
        RECT 1430.205 1387.010 1430.535 1387.025 ;
        RECT 1431.125 1387.010 1431.455 1387.025 ;
        RECT 1430.205 1386.710 1431.455 1387.010 ;
        RECT 1430.205 1386.695 1430.535 1386.710 ;
        RECT 1431.125 1386.695 1431.455 1386.710 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 0.300 ;
=======
      LAYER met1 ;
        RECT 1067.270 28.460 1067.590 28.520 ;
        RECT 1437.110 28.460 1437.430 28.520 ;
        RECT 1067.270 28.320 1437.430 28.460 ;
        RECT 1067.270 28.260 1067.590 28.320 ;
        RECT 1437.110 28.260 1437.430 28.320 ;
      LAYER via ;
        RECT 1067.300 28.260 1067.560 28.520 ;
        RECT 1437.140 28.260 1437.400 28.520 ;
      LAYER met2 ;
        RECT 1438.050 1700.410 1438.330 1704.000 ;
        RECT 1437.200 1700.270 1438.330 1700.410 ;
        RECT 1437.200 28.550 1437.340 1700.270 ;
        RECT 1438.050 1700.000 1438.330 1700.270 ;
        RECT 1067.300 28.230 1067.560 28.550 ;
        RECT 1437.140 28.230 1437.400 28.550 ;
        RECT 1067.360 2.400 1067.500 28.230 ;
=======
      LAYER li1 ;
        RECT 1437.645 227.885 1437.815 275.995 ;
      LAYER mcon ;
        RECT 1437.645 275.825 1437.815 275.995 ;
      LAYER met1 ;
        RECT 1437.570 593.340 1437.890 593.600 ;
        RECT 1437.660 592.920 1437.800 593.340 ;
        RECT 1437.570 592.660 1437.890 592.920 ;
        RECT 1437.570 386.140 1437.890 386.200 ;
        RECT 1438.030 386.140 1438.350 386.200 ;
        RECT 1437.570 386.000 1438.350 386.140 ;
        RECT 1437.570 385.940 1437.890 386.000 ;
        RECT 1438.030 385.940 1438.350 386.000 ;
        RECT 1437.585 275.980 1437.875 276.025 ;
        RECT 1438.030 275.980 1438.350 276.040 ;
        RECT 1437.585 275.840 1438.350 275.980 ;
        RECT 1437.585 275.795 1437.875 275.840 ;
        RECT 1438.030 275.780 1438.350 275.840 ;
        RECT 1437.570 228.040 1437.890 228.100 ;
        RECT 1437.375 227.900 1437.890 228.040 ;
        RECT 1437.570 227.840 1437.890 227.900 ;
        RECT 1437.570 159.020 1437.890 159.080 ;
        RECT 1437.200 158.880 1437.890 159.020 ;
        RECT 1437.200 158.740 1437.340 158.880 ;
        RECT 1437.570 158.820 1437.890 158.880 ;
        RECT 1437.110 158.480 1437.430 158.740 ;
        RECT 1437.110 137.940 1437.430 138.000 ;
        RECT 1438.030 137.940 1438.350 138.000 ;
        RECT 1437.110 137.800 1438.350 137.940 ;
        RECT 1437.110 137.740 1437.430 137.800 ;
        RECT 1438.030 137.740 1438.350 137.800 ;
        RECT 1437.110 48.520 1437.430 48.580 ;
        RECT 1438.030 48.520 1438.350 48.580 ;
        RECT 1437.110 48.380 1438.350 48.520 ;
        RECT 1437.110 48.320 1437.430 48.380 ;
        RECT 1438.030 48.320 1438.350 48.380 ;
        RECT 1067.270 28.120 1067.590 28.180 ;
        RECT 1437.110 28.120 1437.430 28.180 ;
        RECT 1067.270 27.980 1437.430 28.120 ;
        RECT 1067.270 27.920 1067.590 27.980 ;
        RECT 1437.110 27.920 1437.430 27.980 ;
      LAYER via ;
        RECT 1437.600 593.340 1437.860 593.600 ;
        RECT 1437.600 592.660 1437.860 592.920 ;
        RECT 1437.600 385.940 1437.860 386.200 ;
        RECT 1438.060 385.940 1438.320 386.200 ;
        RECT 1438.060 275.780 1438.320 276.040 ;
        RECT 1437.600 227.840 1437.860 228.100 ;
        RECT 1437.600 158.820 1437.860 159.080 ;
        RECT 1437.140 158.480 1437.400 158.740 ;
        RECT 1437.140 137.740 1437.400 138.000 ;
        RECT 1438.060 137.740 1438.320 138.000 ;
        RECT 1437.140 48.320 1437.400 48.580 ;
        RECT 1438.060 48.320 1438.320 48.580 ;
        RECT 1067.300 27.920 1067.560 28.180 ;
        RECT 1437.140 27.920 1437.400 28.180 ;
      LAYER met2 ;
        RECT 1438.970 1700.410 1439.250 1704.000 ;
        RECT 1438.120 1700.270 1439.250 1700.410 ;
        RECT 1438.120 1656.210 1438.260 1700.270 ;
        RECT 1438.970 1700.000 1439.250 1700.270 ;
        RECT 1437.660 1656.070 1438.260 1656.210 ;
        RECT 1437.660 787.170 1437.800 1656.070 ;
        RECT 1437.200 787.030 1437.800 787.170 ;
        RECT 1437.200 786.490 1437.340 787.030 ;
        RECT 1437.200 786.350 1437.800 786.490 ;
        RECT 1437.660 593.630 1437.800 786.350 ;
        RECT 1437.600 593.310 1437.860 593.630 ;
        RECT 1437.600 592.630 1437.860 592.950 ;
        RECT 1437.660 497.490 1437.800 592.630 ;
        RECT 1437.200 497.350 1437.800 497.490 ;
        RECT 1437.200 496.810 1437.340 497.350 ;
        RECT 1437.200 496.670 1437.800 496.810 ;
        RECT 1437.660 386.230 1437.800 496.670 ;
        RECT 1437.600 385.910 1437.860 386.230 ;
        RECT 1438.060 385.910 1438.320 386.230 ;
        RECT 1438.120 276.070 1438.260 385.910 ;
        RECT 1438.060 275.750 1438.320 276.070 ;
        RECT 1437.600 227.810 1437.860 228.130 ;
        RECT 1437.660 159.110 1437.800 227.810 ;
        RECT 1437.600 158.790 1437.860 159.110 ;
        RECT 1437.140 158.450 1437.400 158.770 ;
        RECT 1437.200 138.030 1437.340 158.450 ;
        RECT 1437.140 137.710 1437.400 138.030 ;
        RECT 1438.060 137.710 1438.320 138.030 ;
        RECT 1438.120 48.610 1438.260 137.710 ;
        RECT 1437.140 48.290 1437.400 48.610 ;
        RECT 1438.060 48.290 1438.320 48.610 ;
        RECT 1437.200 28.210 1437.340 48.290 ;
        RECT 1067.300 27.890 1067.560 28.210 ;
        RECT 1437.140 27.890 1437.400 28.210 ;
        RECT 1067.360 2.400 1067.500 27.890 ;
>>>>>>> re-updated local openlane
        RECT 1067.150 -4.800 1067.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1085.210 27.780 1085.530 27.840 ;
        RECT 1443.090 27.780 1443.410 27.840 ;
        RECT 1085.210 27.640 1443.410 27.780 ;
        RECT 1085.210 27.580 1085.530 27.640 ;
        RECT 1443.090 27.580 1443.410 27.640 ;
      LAYER via ;
        RECT 1085.240 27.580 1085.500 27.840 ;
        RECT 1443.120 27.580 1443.380 27.840 ;
      LAYER met2 ;
        RECT 1444.030 1700.410 1444.310 1704.000 ;
        RECT 1443.180 1700.270 1444.310 1700.410 ;
        RECT 1443.180 27.870 1443.320 1700.270 ;
        RECT 1444.030 1700.000 1444.310 1700.270 ;
        RECT 1085.240 27.550 1085.500 27.870 ;
        RECT 1443.120 27.550 1443.380 27.870 ;
        RECT 1085.300 2.400 1085.440 27.550 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 0.300 ;
=======
      LAYER li1 ;
        RECT 1445.005 1545.045 1445.175 1587.035 ;
        RECT 1446.845 1048.645 1447.015 1089.955 ;
        RECT 1445.005 783.105 1445.175 807.075 ;
        RECT 1444.545 620.925 1444.715 628.235 ;
        RECT 1444.545 434.265 1444.715 475.915 ;
        RECT 1444.545 227.885 1444.715 275.995 ;
        RECT 1445.005 131.325 1445.175 159.035 ;
        RECT 1444.085 27.625 1444.255 36.295 ;
      LAYER mcon ;
        RECT 1445.005 1586.865 1445.175 1587.035 ;
        RECT 1446.845 1089.785 1447.015 1089.955 ;
        RECT 1445.005 806.905 1445.175 807.075 ;
        RECT 1444.545 628.065 1444.715 628.235 ;
        RECT 1444.545 475.745 1444.715 475.915 ;
        RECT 1444.545 275.825 1444.715 275.995 ;
        RECT 1445.005 158.865 1445.175 159.035 ;
        RECT 1444.085 36.125 1444.255 36.295 ;
      LAYER met1 ;
        RECT 1444.930 1587.020 1445.250 1587.080 ;
        RECT 1444.735 1586.880 1445.250 1587.020 ;
        RECT 1444.930 1586.820 1445.250 1586.880 ;
        RECT 1444.945 1545.200 1445.235 1545.245 ;
        RECT 1445.390 1545.200 1445.710 1545.260 ;
        RECT 1444.945 1545.060 1445.710 1545.200 ;
        RECT 1444.945 1545.015 1445.235 1545.060 ;
        RECT 1445.390 1545.000 1445.710 1545.060 ;
        RECT 1444.930 1497.600 1445.250 1497.660 ;
        RECT 1445.390 1497.600 1445.710 1497.660 ;
        RECT 1444.930 1497.460 1445.710 1497.600 ;
        RECT 1444.930 1497.400 1445.250 1497.460 ;
        RECT 1445.390 1497.400 1445.710 1497.460 ;
        RECT 1444.930 1463.260 1445.250 1463.320 ;
        RECT 1444.560 1463.120 1445.250 1463.260 ;
        RECT 1444.560 1462.640 1444.700 1463.120 ;
        RECT 1444.930 1463.060 1445.250 1463.120 ;
        RECT 1444.470 1462.380 1444.790 1462.640 ;
        RECT 1444.470 1400.700 1444.790 1400.760 ;
        RECT 1444.930 1400.700 1445.250 1400.760 ;
        RECT 1444.470 1400.560 1445.250 1400.700 ;
        RECT 1444.470 1400.500 1444.790 1400.560 ;
        RECT 1444.930 1400.500 1445.250 1400.560 ;
        RECT 1444.470 1352.560 1444.790 1352.820 ;
        RECT 1444.560 1352.080 1444.700 1352.560 ;
        RECT 1444.930 1352.080 1445.250 1352.140 ;
        RECT 1444.560 1351.940 1445.250 1352.080 ;
        RECT 1444.930 1351.880 1445.250 1351.940 ;
        RECT 1444.470 1249.060 1444.790 1249.120 ;
        RECT 1444.930 1249.060 1445.250 1249.120 ;
        RECT 1444.470 1248.920 1445.250 1249.060 ;
        RECT 1444.470 1248.860 1444.790 1248.920 ;
        RECT 1444.930 1248.860 1445.250 1248.920 ;
        RECT 1444.930 1159.640 1445.250 1159.700 ;
        RECT 1444.560 1159.500 1445.250 1159.640 ;
        RECT 1444.560 1159.360 1444.700 1159.500 ;
        RECT 1444.930 1159.440 1445.250 1159.500 ;
        RECT 1444.470 1159.100 1444.790 1159.360 ;
        RECT 1444.010 1145.360 1444.330 1145.420 ;
        RECT 1444.470 1145.360 1444.790 1145.420 ;
        RECT 1444.010 1145.220 1444.790 1145.360 ;
        RECT 1444.010 1145.160 1444.330 1145.220 ;
        RECT 1444.470 1145.160 1444.790 1145.220 ;
        RECT 1444.930 1097.080 1445.250 1097.140 ;
        RECT 1446.770 1097.080 1447.090 1097.140 ;
        RECT 1444.930 1096.940 1447.090 1097.080 ;
        RECT 1444.930 1096.880 1445.250 1096.940 ;
        RECT 1446.770 1096.880 1447.090 1096.940 ;
        RECT 1446.770 1089.940 1447.090 1090.000 ;
        RECT 1446.575 1089.800 1447.090 1089.940 ;
        RECT 1446.770 1089.740 1447.090 1089.800 ;
        RECT 1446.770 1048.800 1447.090 1048.860 ;
        RECT 1446.575 1048.660 1447.090 1048.800 ;
        RECT 1446.770 1048.600 1447.090 1048.660 ;
        RECT 1444.470 862.820 1444.790 862.880 ;
        RECT 1445.390 862.820 1445.710 862.880 ;
        RECT 1444.470 862.680 1445.710 862.820 ;
        RECT 1444.470 862.620 1444.790 862.680 ;
        RECT 1445.390 862.620 1445.710 862.680 ;
        RECT 1444.930 807.060 1445.250 807.120 ;
        RECT 1444.735 806.920 1445.250 807.060 ;
        RECT 1444.930 806.860 1445.250 806.920 ;
        RECT 1444.930 783.260 1445.250 783.320 ;
        RECT 1444.735 783.120 1445.250 783.260 ;
        RECT 1444.930 783.060 1445.250 783.120 ;
        RECT 1444.930 724.440 1445.250 724.500 ;
        RECT 1445.390 724.440 1445.710 724.500 ;
        RECT 1444.930 724.300 1445.710 724.440 ;
        RECT 1444.930 724.240 1445.250 724.300 ;
        RECT 1445.390 724.240 1445.710 724.300 ;
        RECT 1444.470 676.160 1444.790 676.220 ;
        RECT 1445.390 676.160 1445.710 676.220 ;
        RECT 1444.470 676.020 1445.710 676.160 ;
        RECT 1444.470 675.960 1444.790 676.020 ;
        RECT 1445.390 675.960 1445.710 676.020 ;
        RECT 1444.485 628.220 1444.775 628.265 ;
        RECT 1445.390 628.220 1445.710 628.280 ;
        RECT 1444.485 628.080 1445.710 628.220 ;
        RECT 1444.485 628.035 1444.775 628.080 ;
        RECT 1445.390 628.020 1445.710 628.080 ;
        RECT 1444.470 621.080 1444.790 621.140 ;
        RECT 1444.275 620.940 1444.790 621.080 ;
        RECT 1444.470 620.880 1444.790 620.940 ;
        RECT 1444.470 572.800 1444.790 572.860 ;
        RECT 1445.390 572.800 1445.710 572.860 ;
        RECT 1444.470 572.660 1445.710 572.800 ;
        RECT 1444.470 572.600 1444.790 572.660 ;
        RECT 1445.390 572.600 1445.710 572.660 ;
        RECT 1444.470 475.900 1444.790 475.960 ;
        RECT 1444.275 475.760 1444.790 475.900 ;
        RECT 1444.470 475.700 1444.790 475.760 ;
        RECT 1444.485 434.420 1444.775 434.465 ;
        RECT 1444.930 434.420 1445.250 434.480 ;
        RECT 1444.485 434.280 1445.250 434.420 ;
        RECT 1444.485 434.235 1444.775 434.280 ;
        RECT 1444.930 434.220 1445.250 434.280 ;
        RECT 1444.470 379.680 1444.790 379.740 ;
        RECT 1444.930 379.680 1445.250 379.740 ;
        RECT 1444.470 379.540 1445.250 379.680 ;
        RECT 1444.470 379.480 1444.790 379.540 ;
        RECT 1444.930 379.480 1445.250 379.540 ;
        RECT 1444.470 275.980 1444.790 276.040 ;
        RECT 1444.275 275.840 1444.790 275.980 ;
        RECT 1444.470 275.780 1444.790 275.840 ;
        RECT 1444.470 228.040 1444.790 228.100 ;
        RECT 1444.275 227.900 1444.790 228.040 ;
        RECT 1444.470 227.840 1444.790 227.900 ;
        RECT 1444.930 159.020 1445.250 159.080 ;
        RECT 1444.735 158.880 1445.250 159.020 ;
        RECT 1444.930 158.820 1445.250 158.880 ;
        RECT 1444.930 131.480 1445.250 131.540 ;
        RECT 1444.735 131.340 1445.250 131.480 ;
        RECT 1444.930 131.280 1445.250 131.340 ;
        RECT 1444.010 83.200 1444.330 83.260 ;
        RECT 1444.930 83.200 1445.250 83.260 ;
        RECT 1444.010 83.060 1445.250 83.200 ;
        RECT 1444.010 83.000 1444.330 83.060 ;
        RECT 1444.930 83.000 1445.250 83.060 ;
        RECT 1444.010 36.280 1444.330 36.340 ;
        RECT 1443.815 36.140 1444.330 36.280 ;
        RECT 1444.010 36.080 1444.330 36.140 ;
        RECT 1102.690 27.780 1103.010 27.840 ;
        RECT 1444.025 27.780 1444.315 27.825 ;
        RECT 1102.690 27.640 1444.315 27.780 ;
        RECT 1102.690 27.580 1103.010 27.640 ;
        RECT 1444.025 27.595 1444.315 27.640 ;
      LAYER via ;
        RECT 1444.960 1586.820 1445.220 1587.080 ;
        RECT 1445.420 1545.000 1445.680 1545.260 ;
        RECT 1444.960 1497.400 1445.220 1497.660 ;
        RECT 1445.420 1497.400 1445.680 1497.660 ;
        RECT 1444.960 1463.060 1445.220 1463.320 ;
        RECT 1444.500 1462.380 1444.760 1462.640 ;
        RECT 1444.500 1400.500 1444.760 1400.760 ;
        RECT 1444.960 1400.500 1445.220 1400.760 ;
        RECT 1444.500 1352.560 1444.760 1352.820 ;
        RECT 1444.960 1351.880 1445.220 1352.140 ;
        RECT 1444.500 1248.860 1444.760 1249.120 ;
        RECT 1444.960 1248.860 1445.220 1249.120 ;
        RECT 1444.960 1159.440 1445.220 1159.700 ;
        RECT 1444.500 1159.100 1444.760 1159.360 ;
        RECT 1444.040 1145.160 1444.300 1145.420 ;
        RECT 1444.500 1145.160 1444.760 1145.420 ;
        RECT 1444.960 1096.880 1445.220 1097.140 ;
        RECT 1446.800 1096.880 1447.060 1097.140 ;
        RECT 1446.800 1089.740 1447.060 1090.000 ;
        RECT 1446.800 1048.600 1447.060 1048.860 ;
        RECT 1444.500 862.620 1444.760 862.880 ;
        RECT 1445.420 862.620 1445.680 862.880 ;
        RECT 1444.960 806.860 1445.220 807.120 ;
        RECT 1444.960 783.060 1445.220 783.320 ;
        RECT 1444.960 724.240 1445.220 724.500 ;
        RECT 1445.420 724.240 1445.680 724.500 ;
        RECT 1444.500 675.960 1444.760 676.220 ;
        RECT 1445.420 675.960 1445.680 676.220 ;
        RECT 1445.420 628.020 1445.680 628.280 ;
        RECT 1444.500 620.880 1444.760 621.140 ;
        RECT 1444.500 572.600 1444.760 572.860 ;
        RECT 1445.420 572.600 1445.680 572.860 ;
        RECT 1444.500 475.700 1444.760 475.960 ;
        RECT 1444.960 434.220 1445.220 434.480 ;
        RECT 1444.500 379.480 1444.760 379.740 ;
        RECT 1444.960 379.480 1445.220 379.740 ;
        RECT 1444.500 275.780 1444.760 276.040 ;
        RECT 1444.500 227.840 1444.760 228.100 ;
        RECT 1444.960 158.820 1445.220 159.080 ;
        RECT 1444.960 131.280 1445.220 131.540 ;
        RECT 1444.040 83.000 1444.300 83.260 ;
        RECT 1444.960 83.000 1445.220 83.260 ;
        RECT 1444.040 36.080 1444.300 36.340 ;
        RECT 1102.720 27.580 1102.980 27.840 ;
      LAYER met2 ;
        RECT 1447.710 1700.410 1447.990 1704.000 ;
        RECT 1446.860 1700.270 1447.990 1700.410 ;
        RECT 1446.860 1656.210 1447.000 1700.270 ;
        RECT 1447.710 1700.000 1447.990 1700.270 ;
        RECT 1445.020 1656.070 1447.000 1656.210 ;
        RECT 1445.020 1587.110 1445.160 1656.070 ;
        RECT 1444.960 1586.790 1445.220 1587.110 ;
        RECT 1445.420 1544.970 1445.680 1545.290 ;
        RECT 1445.480 1497.690 1445.620 1544.970 ;
        RECT 1444.960 1497.370 1445.220 1497.690 ;
        RECT 1445.420 1497.370 1445.680 1497.690 ;
        RECT 1445.020 1463.350 1445.160 1497.370 ;
        RECT 1444.960 1463.030 1445.220 1463.350 ;
        RECT 1444.500 1462.350 1444.760 1462.670 ;
        RECT 1444.560 1425.010 1444.700 1462.350 ;
        RECT 1444.560 1424.870 1445.160 1425.010 ;
        RECT 1445.020 1400.790 1445.160 1424.870 ;
        RECT 1444.500 1400.470 1444.760 1400.790 ;
        RECT 1444.960 1400.470 1445.220 1400.790 ;
        RECT 1444.560 1352.850 1444.700 1400.470 ;
        RECT 1444.500 1352.530 1444.760 1352.850 ;
        RECT 1444.960 1351.850 1445.220 1352.170 ;
        RECT 1445.020 1304.650 1445.160 1351.850 ;
        RECT 1444.560 1304.510 1445.160 1304.650 ;
        RECT 1444.560 1249.150 1444.700 1304.510 ;
        RECT 1444.500 1248.830 1444.760 1249.150 ;
        RECT 1444.960 1248.830 1445.220 1249.150 ;
        RECT 1445.020 1159.730 1445.160 1248.830 ;
        RECT 1444.960 1159.410 1445.220 1159.730 ;
        RECT 1444.500 1159.070 1444.760 1159.390 ;
        RECT 1444.560 1145.450 1444.700 1159.070 ;
        RECT 1444.040 1145.130 1444.300 1145.450 ;
        RECT 1444.500 1145.130 1444.760 1145.450 ;
        RECT 1444.100 1097.365 1444.240 1145.130 ;
        RECT 1444.030 1096.995 1444.310 1097.365 ;
        RECT 1444.950 1096.995 1445.230 1097.365 ;
        RECT 1444.960 1096.850 1445.220 1096.995 ;
        RECT 1446.800 1096.850 1447.060 1097.170 ;
        RECT 1446.860 1090.030 1447.000 1096.850 ;
        RECT 1446.800 1089.710 1447.060 1090.030 ;
        RECT 1446.800 1048.570 1447.060 1048.890 ;
        RECT 1446.860 1000.805 1447.000 1048.570 ;
        RECT 1445.410 1000.435 1445.690 1000.805 ;
        RECT 1446.790 1000.435 1447.070 1000.805 ;
        RECT 1445.480 953.205 1445.620 1000.435 ;
        RECT 1445.410 952.835 1445.690 953.205 ;
        RECT 1444.490 952.155 1444.770 952.525 ;
        RECT 1444.560 917.900 1444.700 952.155 ;
        RECT 1444.560 917.760 1445.160 917.900 ;
        RECT 1445.020 883.730 1445.160 917.760 ;
        RECT 1445.020 883.590 1445.620 883.730 ;
        RECT 1445.480 862.910 1445.620 883.590 ;
        RECT 1444.500 862.590 1444.760 862.910 ;
        RECT 1445.420 862.590 1445.680 862.910 ;
        RECT 1444.560 814.370 1444.700 862.590 ;
        RECT 1444.560 814.230 1445.160 814.370 ;
        RECT 1445.020 807.150 1445.160 814.230 ;
        RECT 1444.960 806.830 1445.220 807.150 ;
        RECT 1444.960 783.030 1445.220 783.350 ;
        RECT 1445.020 724.530 1445.160 783.030 ;
        RECT 1444.960 724.210 1445.220 724.530 ;
        RECT 1445.420 724.210 1445.680 724.530 ;
        RECT 1445.480 676.445 1445.620 724.210 ;
        RECT 1444.490 676.075 1444.770 676.445 ;
        RECT 1445.410 676.075 1445.690 676.445 ;
        RECT 1444.500 675.930 1444.760 676.075 ;
        RECT 1445.420 675.930 1445.680 676.075 ;
        RECT 1445.480 628.310 1445.620 675.930 ;
        RECT 1445.420 627.990 1445.680 628.310 ;
        RECT 1444.500 620.850 1444.760 621.170 ;
        RECT 1444.560 572.890 1444.700 620.850 ;
        RECT 1444.500 572.570 1444.760 572.890 ;
        RECT 1445.420 572.570 1445.680 572.890 ;
        RECT 1445.480 537.610 1445.620 572.570 ;
        RECT 1445.480 537.470 1446.080 537.610 ;
        RECT 1445.940 530.810 1446.080 537.470 ;
        RECT 1445.480 530.670 1446.080 530.810 ;
        RECT 1445.480 483.890 1445.620 530.670 ;
        RECT 1445.480 483.750 1446.080 483.890 ;
        RECT 1445.940 476.525 1446.080 483.750 ;
        RECT 1444.950 476.410 1445.230 476.525 ;
        RECT 1444.560 476.270 1445.230 476.410 ;
        RECT 1444.560 475.990 1444.700 476.270 ;
        RECT 1444.950 476.155 1445.230 476.270 ;
        RECT 1445.870 476.155 1446.150 476.525 ;
        RECT 1444.500 475.670 1444.760 475.990 ;
        RECT 1444.960 434.190 1445.220 434.510 ;
        RECT 1445.020 379.770 1445.160 434.190 ;
        RECT 1444.500 379.450 1444.760 379.770 ;
        RECT 1444.960 379.450 1445.220 379.770 ;
        RECT 1444.560 276.070 1444.700 379.450 ;
        RECT 1444.500 275.750 1444.760 276.070 ;
        RECT 1444.500 227.810 1444.760 228.130 ;
        RECT 1444.560 196.250 1444.700 227.810 ;
        RECT 1444.560 196.110 1445.160 196.250 ;
        RECT 1445.020 159.110 1445.160 196.110 ;
        RECT 1444.960 158.790 1445.220 159.110 ;
        RECT 1444.960 131.250 1445.220 131.570 ;
        RECT 1445.020 83.290 1445.160 131.250 ;
        RECT 1444.040 82.970 1444.300 83.290 ;
        RECT 1444.960 82.970 1445.220 83.290 ;
        RECT 1444.100 36.370 1444.240 82.970 ;
        RECT 1444.040 36.050 1444.300 36.370 ;
        RECT 1102.720 27.550 1102.980 27.870 ;
        RECT 1102.780 2.400 1102.920 27.550 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
      LAYER via2 ;
        RECT 1444.030 1097.040 1444.310 1097.320 ;
        RECT 1444.950 1097.040 1445.230 1097.320 ;
        RECT 1445.410 1000.480 1445.690 1000.760 ;
        RECT 1446.790 1000.480 1447.070 1000.760 ;
        RECT 1445.410 952.880 1445.690 953.160 ;
        RECT 1444.490 952.200 1444.770 952.480 ;
        RECT 1444.490 676.120 1444.770 676.400 ;
        RECT 1445.410 676.120 1445.690 676.400 ;
        RECT 1444.950 476.200 1445.230 476.480 ;
        RECT 1445.870 476.200 1446.150 476.480 ;
      LAYER met3 ;
        RECT 1444.005 1097.330 1444.335 1097.345 ;
        RECT 1444.925 1097.330 1445.255 1097.345 ;
        RECT 1444.005 1097.030 1445.255 1097.330 ;
        RECT 1444.005 1097.015 1444.335 1097.030 ;
        RECT 1444.925 1097.015 1445.255 1097.030 ;
        RECT 1445.385 1000.770 1445.715 1000.785 ;
        RECT 1446.765 1000.770 1447.095 1000.785 ;
        RECT 1445.385 1000.470 1447.095 1000.770 ;
        RECT 1445.385 1000.455 1445.715 1000.470 ;
        RECT 1446.765 1000.455 1447.095 1000.470 ;
        RECT 1445.385 953.170 1445.715 953.185 ;
        RECT 1443.790 952.870 1445.715 953.170 ;
        RECT 1443.790 952.490 1444.090 952.870 ;
        RECT 1445.385 952.855 1445.715 952.870 ;
        RECT 1444.465 952.490 1444.795 952.505 ;
        RECT 1443.790 952.190 1444.795 952.490 ;
        RECT 1444.465 952.175 1444.795 952.190 ;
        RECT 1444.465 676.410 1444.795 676.425 ;
        RECT 1445.385 676.410 1445.715 676.425 ;
        RECT 1444.465 676.110 1445.715 676.410 ;
        RECT 1444.465 676.095 1444.795 676.110 ;
        RECT 1445.385 676.095 1445.715 676.110 ;
        RECT 1444.925 476.490 1445.255 476.505 ;
        RECT 1445.845 476.490 1446.175 476.505 ;
        RECT 1444.925 476.190 1446.175 476.490 ;
        RECT 1444.925 476.175 1445.255 476.190 ;
        RECT 1445.845 476.175 1446.175 476.190 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1103.610 1680.860 1103.930 1680.920 ;
        RECT 1448.610 1680.860 1448.930 1680.920 ;
        RECT 1103.610 1680.720 1448.930 1680.860 ;
        RECT 1103.610 1680.660 1103.930 1680.720 ;
        RECT 1448.610 1680.660 1448.930 1680.720 ;
      LAYER via ;
        RECT 1103.640 1680.660 1103.900 1680.920 ;
        RECT 1448.640 1680.660 1448.900 1680.920 ;
      LAYER met2 ;
        RECT 1448.630 1700.000 1448.910 1704.000 ;
        RECT 1448.700 1680.950 1448.840 1700.000 ;
        RECT 1103.640 1680.630 1103.900 1680.950 ;
        RECT 1448.640 1680.630 1448.900 1680.950 ;
        RECT 1103.700 3.130 1103.840 1680.630 ;
        RECT 1103.240 2.990 1103.840 3.130 ;
        RECT 1103.240 2.960 1103.380 2.990 ;
        RECT 1102.780 2.820 1103.380 2.960 ;
        RECT 1102.780 2.400 1102.920 2.820 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 0.300 ;
=======
      LAYER li1 ;
        RECT 1450.985 923.525 1451.155 965.855 ;
      LAYER mcon ;
        RECT 1450.985 965.685 1451.155 965.855 ;
      LAYER met1 ;
        RECT 1450.910 965.840 1451.230 965.900 ;
        RECT 1450.715 965.700 1451.230 965.840 ;
        RECT 1450.910 965.640 1451.230 965.700 ;
        RECT 1450.910 923.680 1451.230 923.740 ;
        RECT 1450.715 923.540 1451.230 923.680 ;
        RECT 1450.910 923.480 1451.230 923.540 ;
        RECT 1124.310 48.860 1124.630 48.920 ;
        RECT 1450.910 48.860 1451.230 48.920 ;
        RECT 1124.310 48.720 1451.230 48.860 ;
        RECT 1124.310 48.660 1124.630 48.720 ;
        RECT 1450.910 48.660 1451.230 48.720 ;
      LAYER via ;
        RECT 1450.940 965.640 1451.200 965.900 ;
        RECT 1450.940 923.480 1451.200 923.740 ;
        RECT 1124.340 48.660 1124.600 48.920 ;
        RECT 1450.940 48.660 1451.200 48.920 ;
      LAYER met2 ;
        RECT 1452.310 1700.410 1452.590 1704.000 ;
        RECT 1451.000 1700.270 1452.590 1700.410 ;
        RECT 1451.000 965.930 1451.140 1700.270 ;
        RECT 1452.310 1700.000 1452.590 1700.270 ;
        RECT 1450.940 965.610 1451.200 965.930 ;
        RECT 1450.940 923.450 1451.200 923.770 ;
        RECT 1451.000 48.950 1451.140 923.450 ;
        RECT 1124.340 48.630 1124.600 48.950 ;
        RECT 1450.940 48.630 1451.200 48.950 ;
        RECT 1124.400 16.050 1124.540 48.630 ;
        RECT 1120.720 15.910 1124.540 16.050 ;
        RECT 1120.720 2.400 1120.860 15.910 ;
=======
      LAYER met1 ;
        RECT 1124.310 1576.820 1124.630 1576.880 ;
        RECT 1450.450 1576.820 1450.770 1576.880 ;
        RECT 1124.310 1576.680 1450.770 1576.820 ;
        RECT 1124.310 1576.620 1124.630 1576.680 ;
        RECT 1450.450 1576.620 1450.770 1576.680 ;
        RECT 1120.630 2.960 1120.950 3.020 ;
        RECT 1124.310 2.960 1124.630 3.020 ;
        RECT 1120.630 2.820 1124.630 2.960 ;
        RECT 1120.630 2.760 1120.950 2.820 ;
        RECT 1124.310 2.760 1124.630 2.820 ;
      LAYER via ;
        RECT 1124.340 1576.620 1124.600 1576.880 ;
        RECT 1450.480 1576.620 1450.740 1576.880 ;
        RECT 1120.660 2.760 1120.920 3.020 ;
        RECT 1124.340 2.760 1124.600 3.020 ;
      LAYER met2 ;
        RECT 1453.690 1700.410 1453.970 1704.000 ;
        RECT 1452.380 1700.270 1453.970 1700.410 ;
        RECT 1452.380 1677.290 1452.520 1700.270 ;
        RECT 1453.690 1700.000 1453.970 1700.270 ;
        RECT 1451.000 1677.150 1452.520 1677.290 ;
        RECT 1451.000 1607.250 1451.140 1677.150 ;
        RECT 1450.540 1607.110 1451.140 1607.250 ;
        RECT 1450.540 1576.910 1450.680 1607.110 ;
        RECT 1124.340 1576.590 1124.600 1576.910 ;
        RECT 1450.480 1576.590 1450.740 1576.910 ;
        RECT 1124.400 3.050 1124.540 1576.590 ;
        RECT 1120.660 2.730 1120.920 3.050 ;
        RECT 1124.340 2.730 1124.600 3.050 ;
        RECT 1120.720 2.400 1120.860 2.730 ;
>>>>>>> re-updated local openlane
        RECT 1120.510 -4.800 1121.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1145.010 1473.120 1145.330 1473.180 ;
        RECT 1457.350 1473.120 1457.670 1473.180 ;
        RECT 1145.010 1472.980 1457.670 1473.120 ;
        RECT 1145.010 1472.920 1145.330 1472.980 ;
        RECT 1457.350 1472.920 1457.670 1472.980 ;
        RECT 1138.570 13.840 1138.890 13.900 ;
        RECT 1145.010 13.840 1145.330 13.900 ;
        RECT 1138.570 13.700 1145.330 13.840 ;
        RECT 1138.570 13.640 1138.890 13.700 ;
        RECT 1145.010 13.640 1145.330 13.700 ;
      LAYER via ;
        RECT 1145.040 1472.920 1145.300 1473.180 ;
        RECT 1457.380 1472.920 1457.640 1473.180 ;
        RECT 1138.600 13.640 1138.860 13.900 ;
        RECT 1145.040 13.640 1145.300 13.900 ;
      LAYER met2 ;
        RECT 1458.290 1700.410 1458.570 1704.000 ;
        RECT 1457.440 1700.270 1458.570 1700.410 ;
        RECT 1457.440 1473.210 1457.580 1700.270 ;
        RECT 1458.290 1700.000 1458.570 1700.270 ;
        RECT 1145.040 1472.890 1145.300 1473.210 ;
        RECT 1457.380 1472.890 1457.640 1473.210 ;
        RECT 1145.100 13.930 1145.240 1472.890 ;
        RECT 1138.600 13.610 1138.860 13.930 ;
        RECT 1145.040 13.610 1145.300 13.930 ;
        RECT 1138.660 2.400 1138.800 13.610 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 0.300 ;
=======
      LAYER met1 ;
        RECT 1459.650 1689.360 1459.970 1689.420 ;
        RECT 1463.330 1689.360 1463.650 1689.420 ;
        RECT 1459.650 1689.220 1463.650 1689.360 ;
        RECT 1459.650 1689.160 1459.970 1689.220 ;
        RECT 1463.330 1689.160 1463.650 1689.220 ;
        RECT 1158.810 79.460 1159.130 79.520 ;
        RECT 1459.650 79.460 1459.970 79.520 ;
        RECT 1158.810 79.320 1459.970 79.460 ;
        RECT 1158.810 79.260 1159.130 79.320 ;
        RECT 1459.650 79.260 1459.970 79.320 ;
      LAYER via ;
        RECT 1459.680 1689.160 1459.940 1689.420 ;
        RECT 1463.360 1689.160 1463.620 1689.420 ;
        RECT 1158.840 79.260 1159.100 79.520 ;
        RECT 1459.680 79.260 1459.940 79.520 ;
      LAYER met2 ;
        RECT 1463.350 1700.000 1463.630 1704.000 ;
        RECT 1463.420 1689.450 1463.560 1700.000 ;
        RECT 1459.680 1689.130 1459.940 1689.450 ;
        RECT 1463.360 1689.130 1463.620 1689.450 ;
        RECT 1459.740 79.550 1459.880 1689.130 ;
        RECT 1158.840 79.230 1159.100 79.550 ;
        RECT 1459.680 79.230 1459.940 79.550 ;
        RECT 1158.900 3.130 1159.040 79.230 ;
        RECT 1156.600 2.990 1159.040 3.130 ;
        RECT 1156.600 2.400 1156.740 2.990 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 674.310 -4.800 674.870 0.300 ;
=======
        RECT 1331.790 1700.410 1332.070 1704.000 ;
        RECT 1331.790 1700.270 1332.460 1700.410 ;
        RECT 1331.790 1700.000 1332.070 1700.270 ;
        RECT 1332.320 34.525 1332.460 1700.270 ;
        RECT 674.450 34.155 674.730 34.525 ;
        RECT 1332.250 34.155 1332.530 34.525 ;
        RECT 674.520 2.400 674.660 34.155 ;
=======
      LAYER li1 ;
        RECT 1332.305 1604.205 1332.475 1642.115 ;
        RECT 1332.305 1490.645 1332.475 1538.755 ;
        RECT 1332.305 1213.205 1332.475 1290.215 ;
        RECT 1333.225 1151.325 1333.395 1193.655 ;
        RECT 1332.305 918.765 1332.475 1000.535 ;
        RECT 1333.685 862.325 1333.855 903.975 ;
        RECT 1333.685 758.965 1333.855 807.075 ;
        RECT 1332.305 662.405 1332.475 710.515 ;
        RECT 1332.305 524.365 1332.475 613.955 ;
      LAYER mcon ;
        RECT 1332.305 1641.945 1332.475 1642.115 ;
        RECT 1332.305 1538.585 1332.475 1538.755 ;
        RECT 1332.305 1290.045 1332.475 1290.215 ;
        RECT 1333.225 1193.485 1333.395 1193.655 ;
        RECT 1332.305 1000.365 1332.475 1000.535 ;
        RECT 1333.685 903.805 1333.855 903.975 ;
        RECT 1333.685 806.905 1333.855 807.075 ;
        RECT 1332.305 710.345 1332.475 710.515 ;
        RECT 1332.305 613.785 1332.475 613.955 ;
      LAYER met1 ;
        RECT 1331.770 1683.920 1332.090 1683.980 ;
        RECT 1332.230 1683.920 1332.550 1683.980 ;
        RECT 1331.770 1683.780 1332.550 1683.920 ;
        RECT 1331.770 1683.720 1332.090 1683.780 ;
        RECT 1332.230 1683.720 1332.550 1683.780 ;
        RECT 1332.230 1642.100 1332.550 1642.160 ;
        RECT 1332.035 1641.960 1332.550 1642.100 ;
        RECT 1332.230 1641.900 1332.550 1641.960 ;
        RECT 1332.245 1604.360 1332.535 1604.405 ;
        RECT 1332.690 1604.360 1333.010 1604.420 ;
        RECT 1332.245 1604.220 1333.010 1604.360 ;
        RECT 1332.245 1604.175 1332.535 1604.220 ;
        RECT 1332.690 1604.160 1333.010 1604.220 ;
        RECT 1332.245 1538.740 1332.535 1538.785 ;
        RECT 1332.690 1538.740 1333.010 1538.800 ;
        RECT 1332.245 1538.600 1333.010 1538.740 ;
        RECT 1332.245 1538.555 1332.535 1538.600 ;
        RECT 1332.690 1538.540 1333.010 1538.600 ;
        RECT 1332.230 1490.800 1332.550 1490.860 ;
        RECT 1332.035 1490.660 1332.550 1490.800 ;
        RECT 1332.230 1490.600 1332.550 1490.660 ;
        RECT 1332.230 1352.760 1332.550 1352.820 ;
        RECT 1332.690 1352.760 1333.010 1352.820 ;
        RECT 1332.230 1352.620 1333.010 1352.760 ;
        RECT 1332.230 1352.560 1332.550 1352.620 ;
        RECT 1332.690 1352.560 1333.010 1352.620 ;
        RECT 1332.230 1297.340 1332.550 1297.400 ;
        RECT 1333.150 1297.340 1333.470 1297.400 ;
        RECT 1332.230 1297.200 1333.470 1297.340 ;
        RECT 1332.230 1297.140 1332.550 1297.200 ;
        RECT 1333.150 1297.140 1333.470 1297.200 ;
        RECT 1332.230 1290.200 1332.550 1290.260 ;
        RECT 1332.035 1290.060 1332.550 1290.200 ;
        RECT 1332.230 1290.000 1332.550 1290.060 ;
        RECT 1332.230 1213.360 1332.550 1213.420 ;
        RECT 1332.035 1213.220 1332.550 1213.360 ;
        RECT 1332.230 1213.160 1332.550 1213.220 ;
        RECT 1333.150 1193.640 1333.470 1193.700 ;
        RECT 1332.955 1193.500 1333.470 1193.640 ;
        RECT 1333.150 1193.440 1333.470 1193.500 ;
        RECT 1333.150 1151.480 1333.470 1151.540 ;
        RECT 1332.955 1151.340 1333.470 1151.480 ;
        RECT 1333.150 1151.280 1333.470 1151.340 ;
        RECT 1332.690 1055.940 1333.010 1056.000 ;
        RECT 1333.150 1055.940 1333.470 1056.000 ;
        RECT 1332.690 1055.800 1333.470 1055.940 ;
        RECT 1332.690 1055.740 1333.010 1055.800 ;
        RECT 1333.150 1055.740 1333.470 1055.800 ;
        RECT 1332.230 1007.320 1332.550 1007.380 ;
        RECT 1333.150 1007.320 1333.470 1007.380 ;
        RECT 1332.230 1007.180 1333.470 1007.320 ;
        RECT 1332.230 1007.120 1332.550 1007.180 ;
        RECT 1333.150 1007.120 1333.470 1007.180 ;
        RECT 1332.245 1000.520 1332.535 1000.565 ;
        RECT 1333.150 1000.520 1333.470 1000.580 ;
        RECT 1332.245 1000.380 1333.470 1000.520 ;
        RECT 1332.245 1000.335 1332.535 1000.380 ;
        RECT 1333.150 1000.320 1333.470 1000.380 ;
        RECT 1332.230 918.920 1332.550 918.980 ;
        RECT 1332.035 918.780 1332.550 918.920 ;
        RECT 1332.230 918.720 1332.550 918.780 ;
        RECT 1332.230 910.760 1332.550 910.820 ;
        RECT 1333.610 910.760 1333.930 910.820 ;
        RECT 1332.230 910.620 1333.930 910.760 ;
        RECT 1332.230 910.560 1332.550 910.620 ;
        RECT 1333.610 910.560 1333.930 910.620 ;
        RECT 1333.610 903.960 1333.930 904.020 ;
        RECT 1333.415 903.820 1333.930 903.960 ;
        RECT 1333.610 903.760 1333.930 903.820 ;
        RECT 1333.610 862.480 1333.930 862.540 ;
        RECT 1333.415 862.340 1333.930 862.480 ;
        RECT 1333.610 862.280 1333.930 862.340 ;
        RECT 1332.230 823.040 1332.550 823.100 ;
        RECT 1333.610 823.040 1333.930 823.100 ;
        RECT 1332.230 822.900 1333.930 823.040 ;
        RECT 1332.230 822.840 1332.550 822.900 ;
        RECT 1333.610 822.840 1333.930 822.900 ;
        RECT 1332.230 814.200 1332.550 814.260 ;
        RECT 1333.610 814.200 1333.930 814.260 ;
        RECT 1332.230 814.060 1333.930 814.200 ;
        RECT 1332.230 814.000 1332.550 814.060 ;
        RECT 1333.610 814.000 1333.930 814.060 ;
        RECT 1333.610 807.060 1333.930 807.120 ;
        RECT 1333.415 806.920 1333.930 807.060 ;
        RECT 1333.610 806.860 1333.930 806.920 ;
        RECT 1333.610 759.120 1333.930 759.180 ;
        RECT 1333.415 758.980 1333.930 759.120 ;
        RECT 1333.610 758.920 1333.930 758.980 ;
        RECT 1332.230 710.500 1332.550 710.560 ;
        RECT 1332.035 710.360 1332.550 710.500 ;
        RECT 1332.230 710.300 1332.550 710.360 ;
        RECT 1332.245 662.560 1332.535 662.605 ;
        RECT 1332.690 662.560 1333.010 662.620 ;
        RECT 1332.245 662.420 1333.010 662.560 ;
        RECT 1332.245 662.375 1332.535 662.420 ;
        RECT 1332.690 662.360 1333.010 662.420 ;
        RECT 1332.245 613.940 1332.535 613.985 ;
        RECT 1332.690 613.940 1333.010 614.000 ;
        RECT 1332.245 613.800 1333.010 613.940 ;
        RECT 1332.245 613.755 1332.535 613.800 ;
        RECT 1332.690 613.740 1333.010 613.800 ;
        RECT 1332.230 524.520 1332.550 524.580 ;
        RECT 1332.035 524.380 1332.550 524.520 ;
        RECT 1332.230 524.320 1332.550 524.380 ;
        RECT 1331.310 476.240 1331.630 476.300 ;
        RECT 1332.690 476.240 1333.010 476.300 ;
        RECT 1331.310 476.100 1333.010 476.240 ;
        RECT 1331.310 476.040 1331.630 476.100 ;
        RECT 1332.690 476.040 1333.010 476.100 ;
        RECT 1331.310 379.340 1331.630 379.400 ;
        RECT 1332.690 379.340 1333.010 379.400 ;
        RECT 1331.310 379.200 1333.010 379.340 ;
        RECT 1331.310 379.140 1331.630 379.200 ;
        RECT 1332.690 379.140 1333.010 379.200 ;
        RECT 1332.230 331.060 1332.550 331.120 ;
        RECT 1332.690 331.060 1333.010 331.120 ;
        RECT 1332.230 330.920 1333.010 331.060 ;
        RECT 1332.230 330.860 1332.550 330.920 ;
        RECT 1332.690 330.860 1333.010 330.920 ;
        RECT 1332.690 255.580 1333.010 255.640 ;
        RECT 1332.320 255.440 1333.010 255.580 ;
        RECT 1332.320 255.300 1332.460 255.440 ;
        RECT 1332.690 255.380 1333.010 255.440 ;
        RECT 1332.230 255.040 1332.550 255.300 ;
        RECT 1331.310 193.360 1331.630 193.420 ;
        RECT 1332.690 193.360 1333.010 193.420 ;
        RECT 1331.310 193.220 1333.010 193.360 ;
        RECT 1331.310 193.160 1331.630 193.220 ;
        RECT 1332.690 193.160 1333.010 193.220 ;
        RECT 1332.690 159.020 1333.010 159.080 ;
        RECT 1332.320 158.880 1333.010 159.020 ;
        RECT 1332.320 158.740 1332.460 158.880 ;
        RECT 1332.690 158.820 1333.010 158.880 ;
        RECT 1332.230 158.480 1332.550 158.740 ;
        RECT 675.810 107.000 676.130 107.060 ;
        RECT 1332.230 107.000 1332.550 107.060 ;
        RECT 675.810 106.860 1332.550 107.000 ;
        RECT 675.810 106.800 676.130 106.860 ;
        RECT 1332.230 106.800 1332.550 106.860 ;
      LAYER via ;
        RECT 1331.800 1683.720 1332.060 1683.980 ;
        RECT 1332.260 1683.720 1332.520 1683.980 ;
        RECT 1332.260 1641.900 1332.520 1642.160 ;
        RECT 1332.720 1604.160 1332.980 1604.420 ;
        RECT 1332.720 1538.540 1332.980 1538.800 ;
        RECT 1332.260 1490.600 1332.520 1490.860 ;
        RECT 1332.260 1352.560 1332.520 1352.820 ;
        RECT 1332.720 1352.560 1332.980 1352.820 ;
        RECT 1332.260 1297.140 1332.520 1297.400 ;
        RECT 1333.180 1297.140 1333.440 1297.400 ;
        RECT 1332.260 1290.000 1332.520 1290.260 ;
        RECT 1332.260 1213.160 1332.520 1213.420 ;
        RECT 1333.180 1193.440 1333.440 1193.700 ;
        RECT 1333.180 1151.280 1333.440 1151.540 ;
        RECT 1332.720 1055.740 1332.980 1056.000 ;
        RECT 1333.180 1055.740 1333.440 1056.000 ;
        RECT 1332.260 1007.120 1332.520 1007.380 ;
        RECT 1333.180 1007.120 1333.440 1007.380 ;
        RECT 1333.180 1000.320 1333.440 1000.580 ;
        RECT 1332.260 918.720 1332.520 918.980 ;
        RECT 1332.260 910.560 1332.520 910.820 ;
        RECT 1333.640 910.560 1333.900 910.820 ;
        RECT 1333.640 903.760 1333.900 904.020 ;
        RECT 1333.640 862.280 1333.900 862.540 ;
        RECT 1332.260 822.840 1332.520 823.100 ;
        RECT 1333.640 822.840 1333.900 823.100 ;
        RECT 1332.260 814.000 1332.520 814.260 ;
        RECT 1333.640 814.000 1333.900 814.260 ;
        RECT 1333.640 806.860 1333.900 807.120 ;
        RECT 1333.640 758.920 1333.900 759.180 ;
        RECT 1332.260 710.300 1332.520 710.560 ;
        RECT 1332.720 662.360 1332.980 662.620 ;
        RECT 1332.720 613.740 1332.980 614.000 ;
        RECT 1332.260 524.320 1332.520 524.580 ;
        RECT 1331.340 476.040 1331.600 476.300 ;
        RECT 1332.720 476.040 1332.980 476.300 ;
        RECT 1331.340 379.140 1331.600 379.400 ;
        RECT 1332.720 379.140 1332.980 379.400 ;
        RECT 1332.260 330.860 1332.520 331.120 ;
        RECT 1332.720 330.860 1332.980 331.120 ;
        RECT 1332.720 255.380 1332.980 255.640 ;
        RECT 1332.260 255.040 1332.520 255.300 ;
        RECT 1331.340 193.160 1331.600 193.420 ;
        RECT 1332.720 193.160 1332.980 193.420 ;
        RECT 1332.720 158.820 1332.980 159.080 ;
        RECT 1332.260 158.480 1332.520 158.740 ;
        RECT 675.840 106.800 676.100 107.060 ;
        RECT 1332.260 106.800 1332.520 107.060 ;
      LAYER met2 ;
        RECT 1332.710 1700.410 1332.990 1704.000 ;
        RECT 1331.860 1700.270 1332.990 1700.410 ;
        RECT 1331.860 1684.010 1332.000 1700.270 ;
        RECT 1332.710 1700.000 1332.990 1700.270 ;
        RECT 1331.800 1683.690 1332.060 1684.010 ;
        RECT 1332.260 1683.690 1332.520 1684.010 ;
        RECT 1332.320 1642.190 1332.460 1683.690 ;
        RECT 1332.260 1641.870 1332.520 1642.190 ;
        RECT 1332.720 1604.130 1332.980 1604.450 ;
        RECT 1332.780 1538.830 1332.920 1604.130 ;
        RECT 1332.720 1538.510 1332.980 1538.830 ;
        RECT 1332.260 1490.570 1332.520 1490.890 ;
        RECT 1332.320 1352.850 1332.460 1490.570 ;
        RECT 1332.260 1352.530 1332.520 1352.850 ;
        RECT 1332.720 1352.530 1332.980 1352.850 ;
        RECT 1332.780 1318.250 1332.920 1352.530 ;
        RECT 1332.780 1318.110 1333.380 1318.250 ;
        RECT 1333.240 1297.430 1333.380 1318.110 ;
        RECT 1332.260 1297.110 1332.520 1297.430 ;
        RECT 1333.180 1297.110 1333.440 1297.430 ;
        RECT 1332.320 1290.290 1332.460 1297.110 ;
        RECT 1332.260 1289.970 1332.520 1290.290 ;
        RECT 1332.260 1213.130 1332.520 1213.450 ;
        RECT 1332.320 1200.610 1332.460 1213.130 ;
        RECT 1332.320 1200.470 1333.380 1200.610 ;
        RECT 1333.240 1193.730 1333.380 1200.470 ;
        RECT 1333.180 1193.410 1333.440 1193.730 ;
        RECT 1333.180 1151.250 1333.440 1151.570 ;
        RECT 1333.240 1124.450 1333.380 1151.250 ;
        RECT 1332.780 1124.310 1333.380 1124.450 ;
        RECT 1332.780 1104.050 1332.920 1124.310 ;
        RECT 1332.780 1103.910 1333.380 1104.050 ;
        RECT 1333.240 1056.030 1333.380 1103.910 ;
        RECT 1332.720 1055.710 1332.980 1056.030 ;
        RECT 1333.180 1055.710 1333.440 1056.030 ;
        RECT 1332.780 1031.290 1332.920 1055.710 ;
        RECT 1332.320 1031.150 1332.920 1031.290 ;
        RECT 1332.320 1007.410 1332.460 1031.150 ;
        RECT 1332.260 1007.090 1332.520 1007.410 ;
        RECT 1333.180 1007.090 1333.440 1007.410 ;
        RECT 1333.240 1000.610 1333.380 1007.090 ;
        RECT 1333.180 1000.290 1333.440 1000.610 ;
        RECT 1332.260 918.690 1332.520 919.010 ;
        RECT 1332.320 910.850 1332.460 918.690 ;
        RECT 1332.260 910.530 1332.520 910.850 ;
        RECT 1333.640 910.530 1333.900 910.850 ;
        RECT 1333.700 904.050 1333.840 910.530 ;
        RECT 1333.640 903.730 1333.900 904.050 ;
        RECT 1333.640 862.250 1333.900 862.570 ;
        RECT 1333.700 823.130 1333.840 862.250 ;
        RECT 1332.260 822.810 1332.520 823.130 ;
        RECT 1333.640 822.810 1333.900 823.130 ;
        RECT 1332.320 814.290 1332.460 822.810 ;
        RECT 1332.260 813.970 1332.520 814.290 ;
        RECT 1333.640 813.970 1333.900 814.290 ;
        RECT 1333.700 807.150 1333.840 813.970 ;
        RECT 1333.640 806.830 1333.900 807.150 ;
        RECT 1333.640 758.890 1333.900 759.210 ;
        RECT 1333.700 723.930 1333.840 758.890 ;
        RECT 1332.780 723.790 1333.840 723.930 ;
        RECT 1332.780 717.810 1332.920 723.790 ;
        RECT 1332.320 717.670 1332.920 717.810 ;
        RECT 1332.320 710.590 1332.460 717.670 ;
        RECT 1332.260 710.270 1332.520 710.590 ;
        RECT 1332.720 662.330 1332.980 662.650 ;
        RECT 1332.780 641.650 1332.920 662.330 ;
        RECT 1332.320 641.510 1332.920 641.650 ;
        RECT 1332.320 620.570 1332.460 641.510 ;
        RECT 1332.320 620.430 1332.920 620.570 ;
        RECT 1332.780 614.030 1332.920 620.430 ;
        RECT 1332.720 613.710 1332.980 614.030 ;
        RECT 1332.260 524.290 1332.520 524.610 ;
        RECT 1332.320 524.125 1332.460 524.290 ;
        RECT 1331.330 523.755 1331.610 524.125 ;
        RECT 1332.250 523.755 1332.530 524.125 ;
        RECT 1331.400 476.330 1331.540 523.755 ;
        RECT 1331.340 476.010 1331.600 476.330 ;
        RECT 1332.720 476.010 1332.980 476.330 ;
        RECT 1332.780 475.730 1332.920 476.010 ;
        RECT 1332.780 475.590 1333.380 475.730 ;
        RECT 1333.240 386.650 1333.380 475.590 ;
        RECT 1332.320 386.510 1333.380 386.650 ;
        RECT 1332.320 379.850 1332.460 386.510 ;
        RECT 1332.320 379.710 1332.920 379.850 ;
        RECT 1332.780 379.430 1332.920 379.710 ;
        RECT 1331.340 379.110 1331.600 379.430 ;
        RECT 1332.720 379.110 1332.980 379.430 ;
        RECT 1331.400 331.685 1331.540 379.110 ;
        RECT 1331.330 331.315 1331.610 331.685 ;
        RECT 1332.250 331.315 1332.530 331.685 ;
        RECT 1332.320 331.150 1332.460 331.315 ;
        RECT 1332.260 330.830 1332.520 331.150 ;
        RECT 1332.720 330.830 1332.980 331.150 ;
        RECT 1332.780 255.670 1332.920 330.830 ;
        RECT 1332.720 255.350 1332.980 255.670 ;
        RECT 1332.260 255.010 1332.520 255.330 ;
        RECT 1332.320 241.245 1332.460 255.010 ;
        RECT 1331.330 240.875 1331.610 241.245 ;
        RECT 1332.250 240.875 1332.530 241.245 ;
        RECT 1331.400 193.450 1331.540 240.875 ;
        RECT 1331.340 193.130 1331.600 193.450 ;
        RECT 1332.720 193.130 1332.980 193.450 ;
        RECT 1332.780 159.110 1332.920 193.130 ;
        RECT 1332.720 158.790 1332.980 159.110 ;
        RECT 1332.260 158.450 1332.520 158.770 ;
        RECT 1332.320 107.090 1332.460 158.450 ;
        RECT 675.840 106.770 676.100 107.090 ;
        RECT 1332.260 106.770 1332.520 107.090 ;
        RECT 675.900 3.130 676.040 106.770 ;
        RECT 674.520 2.990 676.040 3.130 ;
        RECT 674.520 2.400 674.660 2.990 ;
>>>>>>> re-updated local openlane
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 1331.330 523.800 1331.610 524.080 ;
        RECT 1332.250 523.800 1332.530 524.080 ;
        RECT 1331.330 331.360 1331.610 331.640 ;
        RECT 1332.250 331.360 1332.530 331.640 ;
        RECT 1331.330 240.920 1331.610 241.200 ;
        RECT 1332.250 240.920 1332.530 241.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 674.425 34.490 674.755 34.505 ;
        RECT 1332.225 34.490 1332.555 34.505 ;
        RECT 674.425 34.190 1332.555 34.490 ;
        RECT 674.425 34.175 674.755 34.190 ;
        RECT 1332.225 34.175 1332.555 34.190 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1331.305 524.090 1331.635 524.105 ;
        RECT 1332.225 524.090 1332.555 524.105 ;
        RECT 1331.305 523.790 1332.555 524.090 ;
        RECT 1331.305 523.775 1331.635 523.790 ;
        RECT 1332.225 523.775 1332.555 523.790 ;
        RECT 1331.305 331.650 1331.635 331.665 ;
        RECT 1332.225 331.650 1332.555 331.665 ;
        RECT 1331.305 331.350 1332.555 331.650 ;
        RECT 1331.305 331.335 1331.635 331.350 ;
        RECT 1332.225 331.335 1332.555 331.350 ;
        RECT 1331.305 241.210 1331.635 241.225 ;
        RECT 1332.225 241.210 1332.555 241.225 ;
        RECT 1331.305 240.910 1332.555 241.210 ;
        RECT 1331.305 240.895 1331.635 240.910 ;
        RECT 1332.225 240.895 1332.555 240.910 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1463.790 1664.200 1464.110 1664.260 ;
        RECT 1467.010 1664.200 1467.330 1664.260 ;
        RECT 1463.790 1664.060 1467.330 1664.200 ;
        RECT 1463.790 1664.000 1464.110 1664.060 ;
        RECT 1467.010 1664.000 1467.330 1664.060 ;
        RECT 1179.510 58.720 1179.830 58.780 ;
        RECT 1463.790 58.720 1464.110 58.780 ;
        RECT 1179.510 58.580 1464.110 58.720 ;
        RECT 1179.510 58.520 1179.830 58.580 ;
        RECT 1463.790 58.520 1464.110 58.580 ;
        RECT 1173.990 2.960 1174.310 3.020 ;
        RECT 1179.510 2.960 1179.830 3.020 ;
        RECT 1173.990 2.820 1179.830 2.960 ;
        RECT 1173.990 2.760 1174.310 2.820 ;
        RECT 1179.510 2.760 1179.830 2.820 ;
      LAYER via ;
        RECT 1463.820 1664.000 1464.080 1664.260 ;
        RECT 1467.040 1664.000 1467.300 1664.260 ;
        RECT 1179.540 58.520 1179.800 58.780 ;
        RECT 1463.820 58.520 1464.080 58.780 ;
        RECT 1174.020 2.760 1174.280 3.020 ;
        RECT 1179.540 2.760 1179.800 3.020 ;
      LAYER met2 ;
        RECT 1467.950 1700.410 1468.230 1704.000 ;
        RECT 1467.100 1700.270 1468.230 1700.410 ;
        RECT 1467.100 1664.290 1467.240 1700.270 ;
        RECT 1467.950 1700.000 1468.230 1700.270 ;
        RECT 1463.820 1663.970 1464.080 1664.290 ;
        RECT 1467.040 1663.970 1467.300 1664.290 ;
        RECT 1463.880 58.810 1464.020 1663.970 ;
        RECT 1179.540 58.490 1179.800 58.810 ;
        RECT 1463.820 58.490 1464.080 58.810 ;
        RECT 1179.600 3.050 1179.740 58.490 ;
        RECT 1174.020 2.730 1174.280 3.050 ;
        RECT 1179.540 2.730 1179.800 3.050 ;
        RECT 1174.080 2.400 1174.220 2.730 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1174.010 17.200 1174.290 17.480 ;
        RECT 1462.890 17.200 1463.170 17.480 ;
      LAYER met3 ;
        RECT 1173.985 17.490 1174.315 17.505 ;
        RECT 1462.865 17.490 1463.195 17.505 ;
        RECT 1173.985 17.190 1463.195 17.490 ;
        RECT 1173.985 17.175 1174.315 17.190 ;
        RECT 1462.865 17.175 1463.195 17.190 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1191.810 -4.800 1192.370 0.300 ;
=======
        RECT 1471.630 1700.410 1471.910 1704.000 ;
        RECT 1470.320 1700.270 1471.910 1700.410 ;
        RECT 1470.320 18.205 1470.460 1700.270 ;
        RECT 1471.630 1700.000 1471.910 1700.270 ;
        RECT 1191.950 17.835 1192.230 18.205 ;
        RECT 1470.250 17.835 1470.530 18.205 ;
        RECT 1192.020 2.400 1192.160 17.835 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
      LAYER via2 ;
        RECT 1191.950 17.880 1192.230 18.160 ;
        RECT 1470.250 17.880 1470.530 18.160 ;
      LAYER met3 ;
        RECT 1191.925 18.170 1192.255 18.185 ;
        RECT 1470.225 18.170 1470.555 18.185 ;
        RECT 1191.925 17.870 1470.555 18.170 ;
        RECT 1191.925 17.855 1192.255 17.870 ;
        RECT 1470.225 17.855 1470.555 17.870 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1471.610 1665.900 1471.930 1665.960 ;
        RECT 1472.990 1665.900 1473.310 1665.960 ;
        RECT 1471.610 1665.760 1473.310 1665.900 ;
        RECT 1471.610 1665.700 1471.930 1665.760 ;
        RECT 1472.990 1665.700 1473.310 1665.760 ;
        RECT 1193.310 93.060 1193.630 93.120 ;
        RECT 1471.610 93.060 1471.930 93.120 ;
        RECT 1193.310 92.920 1471.930 93.060 ;
        RECT 1193.310 92.860 1193.630 92.920 ;
        RECT 1471.610 92.860 1471.930 92.920 ;
        RECT 1191.930 2.960 1192.250 3.020 ;
        RECT 1193.310 2.960 1193.630 3.020 ;
        RECT 1191.930 2.820 1193.630 2.960 ;
        RECT 1191.930 2.760 1192.250 2.820 ;
        RECT 1193.310 2.760 1193.630 2.820 ;
      LAYER via ;
        RECT 1471.640 1665.700 1471.900 1665.960 ;
        RECT 1473.020 1665.700 1473.280 1665.960 ;
        RECT 1193.340 92.860 1193.600 93.120 ;
        RECT 1471.640 92.860 1471.900 93.120 ;
        RECT 1191.960 2.760 1192.220 3.020 ;
        RECT 1193.340 2.760 1193.600 3.020 ;
      LAYER met2 ;
        RECT 1473.010 1700.000 1473.290 1704.000 ;
        RECT 1473.080 1665.990 1473.220 1700.000 ;
        RECT 1471.640 1665.670 1471.900 1665.990 ;
        RECT 1473.020 1665.670 1473.280 1665.990 ;
        RECT 1471.700 93.150 1471.840 1665.670 ;
        RECT 1193.340 92.830 1193.600 93.150 ;
        RECT 1471.640 92.830 1471.900 93.150 ;
        RECT 1193.400 3.050 1193.540 92.830 ;
        RECT 1191.960 2.730 1192.220 3.050 ;
        RECT 1193.340 2.730 1193.600 3.050 ;
        RECT 1192.020 2.400 1192.160 2.730 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1471.150 1678.480 1471.470 1678.540 ;
        RECT 1475.290 1678.480 1475.610 1678.540 ;
        RECT 1471.150 1678.340 1475.610 1678.480 ;
        RECT 1471.150 1678.280 1471.470 1678.340 ;
        RECT 1475.290 1678.280 1475.610 1678.340 ;
        RECT 1209.870 17.580 1210.190 17.640 ;
        RECT 1471.150 17.580 1471.470 17.640 ;
        RECT 1209.870 17.440 1471.470 17.580 ;
        RECT 1209.870 17.380 1210.190 17.440 ;
        RECT 1471.150 17.380 1471.470 17.440 ;
      LAYER via ;
        RECT 1471.180 1678.280 1471.440 1678.540 ;
        RECT 1475.320 1678.280 1475.580 1678.540 ;
        RECT 1209.900 17.380 1210.160 17.640 ;
        RECT 1471.180 17.380 1471.440 17.640 ;
      LAYER met2 ;
        RECT 1476.230 1700.410 1476.510 1704.000 ;
        RECT 1475.380 1700.270 1476.510 1700.410 ;
        RECT 1475.380 1678.570 1475.520 1700.270 ;
        RECT 1476.230 1700.000 1476.510 1700.270 ;
        RECT 1471.180 1678.250 1471.440 1678.570 ;
        RECT 1475.320 1678.250 1475.580 1678.570 ;
        RECT 1471.240 17.670 1471.380 1678.250 ;
        RECT 1209.900 17.350 1210.160 17.670 ;
        RECT 1471.180 17.350 1471.440 17.670 ;
        RECT 1209.960 2.400 1210.100 17.350 ;
=======
      LAYER li1 ;
        RECT 1438.105 1686.145 1438.275 1689.375 ;
      LAYER mcon ;
        RECT 1438.105 1689.205 1438.275 1689.375 ;
      LAYER met1 ;
        RECT 1438.045 1689.360 1438.335 1689.405 ;
        RECT 1371.880 1689.220 1438.335 1689.360 ;
        RECT 1362.590 1689.020 1362.910 1689.080 ;
        RECT 1371.880 1689.020 1372.020 1689.220 ;
        RECT 1438.045 1689.175 1438.335 1689.220 ;
        RECT 1362.590 1688.880 1372.020 1689.020 ;
        RECT 1362.590 1688.820 1362.910 1688.880 ;
        RECT 1438.045 1686.300 1438.335 1686.345 ;
        RECT 1477.590 1686.300 1477.910 1686.360 ;
        RECT 1438.045 1686.160 1477.910 1686.300 ;
        RECT 1438.045 1686.115 1438.335 1686.160 ;
        RECT 1477.590 1686.100 1477.910 1686.160 ;
        RECT 1214.010 65.860 1214.330 65.920 ;
        RECT 1362.590 65.860 1362.910 65.920 ;
        RECT 1214.010 65.720 1362.910 65.860 ;
        RECT 1214.010 65.660 1214.330 65.720 ;
        RECT 1362.590 65.660 1362.910 65.720 ;
        RECT 1209.870 20.300 1210.190 20.360 ;
        RECT 1214.010 20.300 1214.330 20.360 ;
        RECT 1209.870 20.160 1214.330 20.300 ;
        RECT 1209.870 20.100 1210.190 20.160 ;
        RECT 1214.010 20.100 1214.330 20.160 ;
      LAYER via ;
        RECT 1362.620 1688.820 1362.880 1689.080 ;
        RECT 1477.620 1686.100 1477.880 1686.360 ;
        RECT 1214.040 65.660 1214.300 65.920 ;
        RECT 1362.620 65.660 1362.880 65.920 ;
        RECT 1209.900 20.100 1210.160 20.360 ;
        RECT 1214.040 20.100 1214.300 20.360 ;
      LAYER met2 ;
        RECT 1477.610 1700.000 1477.890 1704.000 ;
        RECT 1362.620 1688.790 1362.880 1689.110 ;
        RECT 1362.680 65.950 1362.820 1688.790 ;
        RECT 1477.680 1686.390 1477.820 1700.000 ;
        RECT 1477.620 1686.070 1477.880 1686.390 ;
        RECT 1214.040 65.630 1214.300 65.950 ;
        RECT 1362.620 65.630 1362.880 65.950 ;
        RECT 1214.100 20.390 1214.240 65.630 ;
        RECT 1209.900 20.070 1210.160 20.390 ;
        RECT 1214.040 20.070 1214.300 20.390 ;
        RECT 1209.960 2.400 1210.100 20.070 ;
>>>>>>> re-updated local openlane
        RECT 1209.750 -4.800 1210.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1477.130 1678.140 1477.450 1678.200 ;
        RECT 1479.890 1678.140 1480.210 1678.200 ;
        RECT 1477.130 1678.000 1480.210 1678.140 ;
        RECT 1477.130 1677.940 1477.450 1678.000 ;
        RECT 1479.890 1677.940 1480.210 1678.000 ;
        RECT 1227.810 18.260 1228.130 18.320 ;
        RECT 1477.130 18.260 1477.450 18.320 ;
        RECT 1227.810 18.120 1423.540 18.260 ;
        RECT 1227.810 18.060 1228.130 18.120 ;
        RECT 1423.400 17.920 1423.540 18.120 ;
        RECT 1464.800 18.120 1477.450 18.260 ;
        RECT 1464.800 17.920 1464.940 18.120 ;
        RECT 1477.130 18.060 1477.450 18.120 ;
        RECT 1423.400 17.780 1464.940 17.920 ;
      LAYER via ;
        RECT 1477.160 1677.940 1477.420 1678.200 ;
        RECT 1479.920 1677.940 1480.180 1678.200 ;
        RECT 1227.840 18.060 1228.100 18.320 ;
        RECT 1477.160 18.060 1477.420 18.320 ;
      LAYER met2 ;
        RECT 1481.290 1700.410 1481.570 1704.000 ;
        RECT 1479.980 1700.270 1481.570 1700.410 ;
        RECT 1479.980 1678.230 1480.120 1700.270 ;
        RECT 1481.290 1700.000 1481.570 1700.270 ;
        RECT 1477.160 1677.910 1477.420 1678.230 ;
        RECT 1479.920 1677.910 1480.180 1678.230 ;
        RECT 1477.220 18.350 1477.360 1677.910 ;
        RECT 1227.840 18.030 1228.100 18.350 ;
        RECT 1477.160 18.030 1477.420 18.350 ;
        RECT 1227.900 2.400 1228.040 18.030 ;
=======
      LAYER li1 ;
        RECT 1227.885 13.685 1228.055 17.595 ;
      LAYER mcon ;
        RECT 1227.885 17.425 1228.055 17.595 ;
      LAYER met1 ;
        RECT 1459.190 1690.380 1459.510 1690.440 ;
        RECT 1481.270 1690.380 1481.590 1690.440 ;
        RECT 1459.190 1690.240 1481.590 1690.380 ;
        RECT 1459.190 1690.180 1459.510 1690.240 ;
        RECT 1481.270 1690.180 1481.590 1690.240 ;
        RECT 1227.350 72.660 1227.670 72.720 ;
        RECT 1459.190 72.660 1459.510 72.720 ;
        RECT 1227.350 72.520 1459.510 72.660 ;
        RECT 1227.350 72.460 1227.670 72.520 ;
        RECT 1459.190 72.460 1459.510 72.520 ;
        RECT 1227.350 17.580 1227.670 17.640 ;
        RECT 1227.825 17.580 1228.115 17.625 ;
        RECT 1227.350 17.440 1228.115 17.580 ;
        RECT 1227.350 17.380 1227.670 17.440 ;
        RECT 1227.825 17.395 1228.115 17.440 ;
        RECT 1227.810 13.840 1228.130 13.900 ;
        RECT 1227.615 13.700 1228.130 13.840 ;
        RECT 1227.810 13.640 1228.130 13.700 ;
      LAYER via ;
        RECT 1459.220 1690.180 1459.480 1690.440 ;
        RECT 1481.300 1690.180 1481.560 1690.440 ;
        RECT 1227.380 72.460 1227.640 72.720 ;
        RECT 1459.220 72.460 1459.480 72.720 ;
        RECT 1227.380 17.380 1227.640 17.640 ;
        RECT 1227.840 13.640 1228.100 13.900 ;
      LAYER met2 ;
        RECT 1482.670 1700.410 1482.950 1704.000 ;
        RECT 1481.360 1700.270 1482.950 1700.410 ;
        RECT 1481.360 1690.470 1481.500 1700.270 ;
        RECT 1482.670 1700.000 1482.950 1700.270 ;
        RECT 1459.220 1690.150 1459.480 1690.470 ;
        RECT 1481.300 1690.150 1481.560 1690.470 ;
        RECT 1459.280 72.750 1459.420 1690.150 ;
        RECT 1227.380 72.430 1227.640 72.750 ;
        RECT 1459.220 72.430 1459.480 72.750 ;
        RECT 1227.440 17.670 1227.580 72.430 ;
        RECT 1227.380 17.350 1227.640 17.670 ;
        RECT 1227.840 13.610 1228.100 13.930 ;
        RECT 1227.900 2.400 1228.040 13.610 ;
>>>>>>> re-updated local openlane
        RECT 1227.690 -4.800 1228.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1484.490 1678.140 1484.810 1678.200 ;
        RECT 1486.330 1678.140 1486.650 1678.200 ;
        RECT 1484.490 1678.000 1486.650 1678.140 ;
        RECT 1484.490 1677.940 1484.810 1678.000 ;
        RECT 1486.330 1677.940 1486.650 1678.000 ;
        RECT 1245.750 37.980 1246.070 38.040 ;
        RECT 1484.490 37.980 1484.810 38.040 ;
        RECT 1245.750 37.840 1484.810 37.980 ;
        RECT 1245.750 37.780 1246.070 37.840 ;
        RECT 1484.490 37.780 1484.810 37.840 ;
      LAYER via ;
        RECT 1484.520 1677.940 1484.780 1678.200 ;
        RECT 1486.360 1677.940 1486.620 1678.200 ;
        RECT 1245.780 37.780 1246.040 38.040 ;
        RECT 1484.520 37.780 1484.780 38.040 ;
      LAYER met2 ;
        RECT 1487.270 1700.410 1487.550 1704.000 ;
        RECT 1486.420 1700.270 1487.550 1700.410 ;
        RECT 1486.420 1678.230 1486.560 1700.270 ;
        RECT 1487.270 1700.000 1487.550 1700.270 ;
        RECT 1484.520 1677.910 1484.780 1678.230 ;
        RECT 1486.360 1677.910 1486.620 1678.230 ;
        RECT 1484.580 38.070 1484.720 1677.910 ;
        RECT 1245.780 37.750 1246.040 38.070 ;
        RECT 1484.520 37.750 1484.780 38.070 ;
        RECT 1245.840 2.400 1245.980 37.750 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1263.230 38.320 1263.550 38.380 ;
        RECT 1491.850 38.320 1492.170 38.380 ;
        RECT 1263.230 38.180 1492.170 38.320 ;
        RECT 1263.230 38.120 1263.550 38.180 ;
        RECT 1491.850 38.120 1492.170 38.180 ;
      LAYER via ;
        RECT 1263.260 38.120 1263.520 38.380 ;
        RECT 1491.880 38.120 1492.140 38.380 ;
      LAYER met2 ;
        RECT 1492.330 1700.410 1492.610 1704.000 ;
        RECT 1491.940 1700.270 1492.610 1700.410 ;
        RECT 1491.940 38.410 1492.080 1700.270 ;
        RECT 1492.330 1700.000 1492.610 1700.270 ;
        RECT 1263.260 38.090 1263.520 38.410 ;
        RECT 1491.880 38.090 1492.140 38.410 ;
        RECT 1263.320 2.400 1263.460 38.090 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1491.390 1678.140 1491.710 1678.200 ;
        RECT 1495.990 1678.140 1496.310 1678.200 ;
        RECT 1491.390 1678.000 1496.310 1678.140 ;
        RECT 1491.390 1677.940 1491.710 1678.000 ;
        RECT 1495.990 1677.940 1496.310 1678.000 ;
        RECT 1281.170 38.660 1281.490 38.720 ;
        RECT 1491.390 38.660 1491.710 38.720 ;
        RECT 1281.170 38.520 1491.710 38.660 ;
        RECT 1281.170 38.460 1281.490 38.520 ;
        RECT 1491.390 38.460 1491.710 38.520 ;
      LAYER via ;
        RECT 1491.420 1677.940 1491.680 1678.200 ;
        RECT 1496.020 1677.940 1496.280 1678.200 ;
        RECT 1281.200 38.460 1281.460 38.720 ;
        RECT 1491.420 38.460 1491.680 38.720 ;
      LAYER met2 ;
        RECT 1496.930 1700.410 1497.210 1704.000 ;
        RECT 1496.080 1700.270 1497.210 1700.410 ;
        RECT 1496.080 1678.230 1496.220 1700.270 ;
        RECT 1496.930 1700.000 1497.210 1700.270 ;
        RECT 1491.420 1677.910 1491.680 1678.230 ;
        RECT 1496.020 1677.910 1496.280 1678.230 ;
        RECT 1491.480 38.750 1491.620 1677.910 ;
        RECT 1281.200 38.430 1281.460 38.750 ;
        RECT 1491.420 38.430 1491.680 38.750 ;
        RECT 1281.260 2.400 1281.400 38.430 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1487.710 18.600 1488.030 18.660 ;
        RECT 1498.290 18.600 1498.610 18.660 ;
        RECT 1487.710 18.460 1498.610 18.600 ;
        RECT 1487.710 18.400 1488.030 18.460 ;
        RECT 1498.290 18.400 1498.610 18.460 ;
        RECT 1299.110 17.920 1299.430 17.980 ;
        RECT 1485.410 17.920 1485.730 17.980 ;
        RECT 1299.110 17.780 1485.730 17.920 ;
        RECT 1299.110 17.720 1299.430 17.780 ;
        RECT 1485.410 17.720 1485.730 17.780 ;
      LAYER via ;
        RECT 1487.740 18.400 1488.000 18.660 ;
        RECT 1498.320 18.400 1498.580 18.660 ;
        RECT 1299.140 17.720 1299.400 17.980 ;
        RECT 1485.440 17.720 1485.700 17.980 ;
      LAYER met2 ;
        RECT 1501.990 1700.410 1502.270 1704.000 ;
        RECT 1500.680 1700.270 1502.270 1700.410 ;
        RECT 1500.680 1675.930 1500.820 1700.270 ;
        RECT 1501.990 1700.000 1502.270 1700.270 ;
        RECT 1498.380 1675.790 1500.820 1675.930 ;
        RECT 1498.380 18.690 1498.520 1675.790 ;
        RECT 1487.740 18.370 1488.000 18.690 ;
        RECT 1498.320 18.370 1498.580 18.690 ;
        RECT 1487.800 18.090 1487.940 18.370 ;
        RECT 1485.500 18.010 1487.940 18.090 ;
        RECT 1299.140 17.690 1299.400 18.010 ;
        RECT 1485.440 17.950 1487.940 18.010 ;
        RECT 1485.440 17.690 1485.700 17.950 ;
        RECT 1299.200 2.400 1299.340 17.690 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 0.300 ;
=======
      LAYER li1 ;
        RECT 1317.585 1684.105 1317.755 1687.335 ;
        RECT 1317.585 1580.065 1317.755 1594.175 ;
        RECT 1317.585 1207.425 1317.755 1255.875 ;
        RECT 1317.585 766.105 1317.755 814.215 ;
        RECT 1317.585 379.525 1317.755 427.635 ;
        RECT 1317.585 282.965 1317.755 331.075 ;
        RECT 1317.585 145.265 1317.755 234.515 ;
        RECT 1317.125 48.365 1317.295 137.615 ;
      LAYER mcon ;
        RECT 1317.585 1687.165 1317.755 1687.335 ;
        RECT 1317.585 1594.005 1317.755 1594.175 ;
        RECT 1317.585 1255.705 1317.755 1255.875 ;
        RECT 1317.585 814.045 1317.755 814.215 ;
        RECT 1317.585 427.465 1317.755 427.635 ;
        RECT 1317.585 330.905 1317.755 331.075 ;
        RECT 1317.585 234.345 1317.755 234.515 ;
        RECT 1317.125 137.445 1317.295 137.615 ;
      LAYER met1 ;
        RECT 1317.525 1687.320 1317.815 1687.365 ;
        RECT 1506.570 1687.320 1506.890 1687.380 ;
        RECT 1317.525 1687.180 1506.890 1687.320 ;
        RECT 1317.525 1687.135 1317.815 1687.180 ;
        RECT 1506.570 1687.120 1506.890 1687.180 ;
        RECT 1317.510 1684.260 1317.830 1684.320 ;
        RECT 1317.315 1684.120 1317.830 1684.260 ;
        RECT 1317.510 1684.060 1317.830 1684.120 ;
        RECT 1317.510 1642.240 1317.830 1642.500 ;
        RECT 1317.600 1641.760 1317.740 1642.240 ;
        RECT 1317.970 1641.760 1318.290 1641.820 ;
        RECT 1317.600 1641.620 1318.290 1641.760 ;
        RECT 1317.970 1641.560 1318.290 1641.620 ;
        RECT 1317.510 1594.160 1317.830 1594.220 ;
        RECT 1317.315 1594.020 1317.830 1594.160 ;
        RECT 1317.510 1593.960 1317.830 1594.020 ;
        RECT 1317.510 1580.220 1317.830 1580.280 ;
        RECT 1317.315 1580.080 1317.830 1580.220 ;
        RECT 1317.510 1580.020 1317.830 1580.080 ;
        RECT 1316.590 1531.940 1316.910 1532.000 ;
        RECT 1317.510 1531.940 1317.830 1532.000 ;
        RECT 1316.590 1531.800 1317.830 1531.940 ;
        RECT 1316.590 1531.740 1316.910 1531.800 ;
        RECT 1317.510 1531.740 1317.830 1531.800 ;
        RECT 1317.050 1483.660 1317.370 1483.720 ;
        RECT 1317.970 1483.660 1318.290 1483.720 ;
        RECT 1317.050 1483.520 1318.290 1483.660 ;
        RECT 1317.050 1483.460 1317.370 1483.520 ;
        RECT 1317.970 1483.460 1318.290 1483.520 ;
        RECT 1317.050 1442.180 1317.370 1442.240 ;
        RECT 1317.510 1442.180 1317.830 1442.240 ;
        RECT 1317.050 1442.040 1317.830 1442.180 ;
        RECT 1317.050 1441.980 1317.370 1442.040 ;
        RECT 1317.510 1441.980 1317.830 1442.040 ;
        RECT 1317.510 1255.860 1317.830 1255.920 ;
        RECT 1317.315 1255.720 1317.830 1255.860 ;
        RECT 1317.510 1255.660 1317.830 1255.720 ;
        RECT 1317.510 1207.580 1317.830 1207.640 ;
        RECT 1317.315 1207.440 1317.830 1207.580 ;
        RECT 1317.510 1207.380 1317.830 1207.440 ;
        RECT 1317.510 1152.500 1317.830 1152.560 ;
        RECT 1318.430 1152.500 1318.750 1152.560 ;
        RECT 1317.510 1152.360 1318.750 1152.500 ;
        RECT 1317.510 1152.300 1317.830 1152.360 ;
        RECT 1318.430 1152.300 1318.750 1152.360 ;
        RECT 1317.510 1007.320 1317.830 1007.380 ;
        RECT 1318.430 1007.320 1318.750 1007.380 ;
        RECT 1317.510 1007.180 1318.750 1007.320 ;
        RECT 1317.510 1007.120 1317.830 1007.180 ;
        RECT 1318.430 1007.120 1318.750 1007.180 ;
        RECT 1317.510 910.760 1317.830 910.820 ;
        RECT 1318.430 910.760 1318.750 910.820 ;
        RECT 1317.510 910.620 1318.750 910.760 ;
        RECT 1317.510 910.560 1317.830 910.620 ;
        RECT 1318.430 910.560 1318.750 910.620 ;
        RECT 1317.510 814.200 1317.830 814.260 ;
        RECT 1317.315 814.060 1317.830 814.200 ;
        RECT 1317.510 814.000 1317.830 814.060 ;
        RECT 1317.510 766.260 1317.830 766.320 ;
        RECT 1317.315 766.120 1317.830 766.260 ;
        RECT 1317.510 766.060 1317.830 766.120 ;
        RECT 1317.510 427.620 1317.830 427.680 ;
        RECT 1317.315 427.480 1317.830 427.620 ;
        RECT 1317.510 427.420 1317.830 427.480 ;
        RECT 1317.510 379.680 1317.830 379.740 ;
        RECT 1317.315 379.540 1317.830 379.680 ;
        RECT 1317.510 379.480 1317.830 379.540 ;
        RECT 1317.510 331.060 1317.830 331.120 ;
        RECT 1317.315 330.920 1317.830 331.060 ;
        RECT 1317.510 330.860 1317.830 330.920 ;
        RECT 1317.525 283.120 1317.815 283.165 ;
        RECT 1317.970 283.120 1318.290 283.180 ;
        RECT 1317.525 282.980 1318.290 283.120 ;
        RECT 1317.525 282.935 1317.815 282.980 ;
        RECT 1317.970 282.920 1318.290 282.980 ;
        RECT 1317.510 234.500 1317.830 234.560 ;
        RECT 1317.315 234.360 1317.830 234.500 ;
        RECT 1317.510 234.300 1317.830 234.360 ;
        RECT 1317.510 145.420 1317.830 145.480 ;
        RECT 1317.315 145.280 1317.830 145.420 ;
        RECT 1317.510 145.220 1317.830 145.280 ;
        RECT 1317.510 137.740 1317.830 138.000 ;
        RECT 1317.065 137.600 1317.355 137.645 ;
        RECT 1317.600 137.600 1317.740 137.740 ;
        RECT 1317.065 137.460 1317.740 137.600 ;
        RECT 1317.065 137.415 1317.355 137.460 ;
        RECT 1317.050 48.520 1317.370 48.580 ;
        RECT 1316.855 48.380 1317.370 48.520 ;
        RECT 1317.050 48.320 1317.370 48.380 ;
      LAYER via ;
        RECT 1506.600 1687.120 1506.860 1687.380 ;
        RECT 1317.540 1684.060 1317.800 1684.320 ;
        RECT 1317.540 1642.240 1317.800 1642.500 ;
        RECT 1318.000 1641.560 1318.260 1641.820 ;
        RECT 1317.540 1593.960 1317.800 1594.220 ;
        RECT 1317.540 1580.020 1317.800 1580.280 ;
        RECT 1316.620 1531.740 1316.880 1532.000 ;
        RECT 1317.540 1531.740 1317.800 1532.000 ;
        RECT 1317.080 1483.460 1317.340 1483.720 ;
        RECT 1318.000 1483.460 1318.260 1483.720 ;
        RECT 1317.080 1441.980 1317.340 1442.240 ;
        RECT 1317.540 1441.980 1317.800 1442.240 ;
        RECT 1317.540 1255.660 1317.800 1255.920 ;
        RECT 1317.540 1207.380 1317.800 1207.640 ;
        RECT 1317.540 1152.300 1317.800 1152.560 ;
        RECT 1318.460 1152.300 1318.720 1152.560 ;
        RECT 1317.540 1007.120 1317.800 1007.380 ;
        RECT 1318.460 1007.120 1318.720 1007.380 ;
        RECT 1317.540 910.560 1317.800 910.820 ;
        RECT 1318.460 910.560 1318.720 910.820 ;
        RECT 1317.540 814.000 1317.800 814.260 ;
        RECT 1317.540 766.060 1317.800 766.320 ;
        RECT 1317.540 427.420 1317.800 427.680 ;
        RECT 1317.540 379.480 1317.800 379.740 ;
        RECT 1317.540 330.860 1317.800 331.120 ;
        RECT 1318.000 282.920 1318.260 283.180 ;
        RECT 1317.540 234.300 1317.800 234.560 ;
        RECT 1317.540 145.220 1317.800 145.480 ;
        RECT 1317.540 137.740 1317.800 138.000 ;
        RECT 1317.080 48.320 1317.340 48.580 ;
      LAYER met2 ;
        RECT 1506.590 1700.000 1506.870 1704.000 ;
        RECT 1506.660 1687.410 1506.800 1700.000 ;
        RECT 1506.600 1687.090 1506.860 1687.410 ;
        RECT 1317.540 1684.030 1317.800 1684.350 ;
        RECT 1317.600 1642.530 1317.740 1684.030 ;
        RECT 1317.540 1642.210 1317.800 1642.530 ;
        RECT 1318.000 1641.530 1318.260 1641.850 ;
        RECT 1318.060 1628.330 1318.200 1641.530 ;
        RECT 1317.600 1628.190 1318.200 1628.330 ;
        RECT 1317.600 1594.250 1317.740 1628.190 ;
        RECT 1317.540 1593.930 1317.800 1594.250 ;
        RECT 1317.540 1579.990 1317.800 1580.310 ;
        RECT 1317.600 1532.030 1317.740 1579.990 ;
        RECT 1316.620 1531.770 1316.880 1532.030 ;
        RECT 1317.070 1531.770 1317.350 1531.885 ;
        RECT 1316.620 1531.710 1317.350 1531.770 ;
        RECT 1317.540 1531.710 1317.800 1532.030 ;
        RECT 1316.680 1531.630 1317.350 1531.710 ;
        RECT 1317.070 1531.515 1317.350 1531.630 ;
        RECT 1317.990 1531.515 1318.270 1531.885 ;
        RECT 1318.060 1483.750 1318.200 1531.515 ;
        RECT 1317.080 1483.430 1317.340 1483.750 ;
        RECT 1318.000 1483.430 1318.260 1483.750 ;
        RECT 1317.140 1442.270 1317.280 1483.430 ;
        RECT 1317.080 1441.950 1317.340 1442.270 ;
        RECT 1317.540 1441.950 1317.800 1442.270 ;
        RECT 1317.600 1255.950 1317.740 1441.950 ;
        RECT 1317.540 1255.630 1317.800 1255.950 ;
        RECT 1317.540 1207.350 1317.800 1207.670 ;
        RECT 1317.600 1200.725 1317.740 1207.350 ;
        RECT 1317.530 1200.355 1317.810 1200.725 ;
        RECT 1318.450 1200.355 1318.730 1200.725 ;
        RECT 1318.520 1152.590 1318.660 1200.355 ;
        RECT 1317.540 1152.270 1317.800 1152.590 ;
        RECT 1318.460 1152.270 1318.720 1152.590 ;
        RECT 1317.600 1104.165 1317.740 1152.270 ;
        RECT 1317.530 1103.795 1317.810 1104.165 ;
        RECT 1318.450 1103.795 1318.730 1104.165 ;
        RECT 1318.520 1055.885 1318.660 1103.795 ;
        RECT 1317.530 1055.515 1317.810 1055.885 ;
        RECT 1318.450 1055.515 1318.730 1055.885 ;
        RECT 1317.600 1007.410 1317.740 1055.515 ;
        RECT 1317.540 1007.090 1317.800 1007.410 ;
        RECT 1318.460 1007.090 1318.720 1007.410 ;
        RECT 1318.520 959.325 1318.660 1007.090 ;
        RECT 1317.530 958.955 1317.810 959.325 ;
        RECT 1318.450 958.955 1318.730 959.325 ;
        RECT 1317.600 910.850 1317.740 958.955 ;
        RECT 1317.540 910.530 1317.800 910.850 ;
        RECT 1318.460 910.530 1318.720 910.850 ;
        RECT 1318.520 862.765 1318.660 910.530 ;
        RECT 1317.530 862.395 1317.810 862.765 ;
        RECT 1318.450 862.395 1318.730 862.765 ;
        RECT 1317.600 814.290 1317.740 862.395 ;
        RECT 1317.540 813.970 1317.800 814.290 ;
        RECT 1317.540 766.030 1317.800 766.350 ;
        RECT 1317.600 427.710 1317.740 766.030 ;
        RECT 1317.540 427.390 1317.800 427.710 ;
        RECT 1317.540 379.450 1317.800 379.770 ;
        RECT 1317.600 331.150 1317.740 379.450 ;
        RECT 1317.540 330.830 1317.800 331.150 ;
        RECT 1318.000 282.890 1318.260 283.210 ;
        RECT 1318.060 241.810 1318.200 282.890 ;
        RECT 1317.600 241.670 1318.200 241.810 ;
        RECT 1317.600 234.590 1317.740 241.670 ;
        RECT 1317.540 234.270 1317.800 234.590 ;
        RECT 1317.540 145.190 1317.800 145.510 ;
        RECT 1317.600 138.030 1317.740 145.190 ;
        RECT 1317.540 137.710 1317.800 138.030 ;
        RECT 1317.080 48.290 1317.340 48.610 ;
        RECT 1317.140 2.400 1317.280 48.290 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
      LAYER via2 ;
        RECT 1317.070 1531.560 1317.350 1531.840 ;
        RECT 1317.990 1531.560 1318.270 1531.840 ;
        RECT 1317.530 1200.400 1317.810 1200.680 ;
        RECT 1318.450 1200.400 1318.730 1200.680 ;
        RECT 1317.530 1103.840 1317.810 1104.120 ;
        RECT 1318.450 1103.840 1318.730 1104.120 ;
        RECT 1317.530 1055.560 1317.810 1055.840 ;
        RECT 1318.450 1055.560 1318.730 1055.840 ;
        RECT 1317.530 959.000 1317.810 959.280 ;
        RECT 1318.450 959.000 1318.730 959.280 ;
        RECT 1317.530 862.440 1317.810 862.720 ;
        RECT 1318.450 862.440 1318.730 862.720 ;
      LAYER met3 ;
        RECT 1317.045 1531.850 1317.375 1531.865 ;
        RECT 1317.965 1531.850 1318.295 1531.865 ;
        RECT 1317.045 1531.550 1318.295 1531.850 ;
        RECT 1317.045 1531.535 1317.375 1531.550 ;
        RECT 1317.965 1531.535 1318.295 1531.550 ;
        RECT 1317.505 1200.690 1317.835 1200.705 ;
        RECT 1318.425 1200.690 1318.755 1200.705 ;
        RECT 1317.505 1200.390 1318.755 1200.690 ;
        RECT 1317.505 1200.375 1317.835 1200.390 ;
<<<<<<< HEAD
        RECT 1317.045 1007.570 1317.375 1007.585 ;
        RECT 1317.045 1007.270 1318.050 1007.570 ;
        RECT 1317.045 1007.255 1317.375 1007.270 ;
        RECT 1317.045 1006.890 1317.375 1006.905 ;
        RECT 1317.750 1006.890 1318.050 1007.270 ;
        RECT 1317.045 1006.590 1318.050 1006.890 ;
        RECT 1317.045 1006.575 1317.375 1006.590 ;
        RECT 1316.585 911.010 1316.915 911.025 ;
        RECT 1317.505 911.010 1317.835 911.025 ;
        RECT 1316.585 910.710 1317.835 911.010 ;
        RECT 1316.585 910.695 1316.915 910.710 ;
        RECT 1317.505 910.695 1317.835 910.710 ;
        RECT 1316.585 669.610 1316.915 669.625 ;
        RECT 1317.505 669.610 1317.835 669.625 ;
        RECT 1316.585 669.310 1317.835 669.610 ;
        RECT 1316.585 669.295 1316.915 669.310 ;
        RECT 1317.505 669.295 1317.835 669.310 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1318.425 1200.375 1318.755 1200.390 ;
        RECT 1317.505 1104.130 1317.835 1104.145 ;
        RECT 1318.425 1104.130 1318.755 1104.145 ;
        RECT 1317.505 1103.830 1318.755 1104.130 ;
        RECT 1317.505 1103.815 1317.835 1103.830 ;
        RECT 1318.425 1103.815 1318.755 1103.830 ;
        RECT 1317.505 1055.850 1317.835 1055.865 ;
        RECT 1318.425 1055.850 1318.755 1055.865 ;
        RECT 1317.505 1055.550 1318.755 1055.850 ;
        RECT 1317.505 1055.535 1317.835 1055.550 ;
        RECT 1318.425 1055.535 1318.755 1055.550 ;
        RECT 1317.505 959.290 1317.835 959.305 ;
        RECT 1318.425 959.290 1318.755 959.305 ;
        RECT 1317.505 958.990 1318.755 959.290 ;
        RECT 1317.505 958.975 1317.835 958.990 ;
        RECT 1318.425 958.975 1318.755 958.990 ;
        RECT 1317.505 862.730 1317.835 862.745 ;
        RECT 1318.425 862.730 1318.755 862.745 ;
        RECT 1317.505 862.430 1318.755 862.730 ;
        RECT 1317.505 862.415 1317.835 862.430 ;
        RECT 1318.425 862.415 1318.755 862.430 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1338.210 1688.000 1338.530 1688.060 ;
        RECT 1511.630 1688.000 1511.950 1688.060 ;
        RECT 1338.210 1687.860 1511.950 1688.000 ;
        RECT 1338.210 1687.800 1338.530 1687.860 ;
        RECT 1511.630 1687.800 1511.950 1687.860 ;
        RECT 1334.990 20.640 1335.310 20.700 ;
        RECT 1338.210 20.640 1338.530 20.700 ;
        RECT 1334.990 20.500 1338.530 20.640 ;
        RECT 1334.990 20.440 1335.310 20.500 ;
        RECT 1338.210 20.440 1338.530 20.500 ;
      LAYER via ;
        RECT 1338.240 1687.800 1338.500 1688.060 ;
        RECT 1511.660 1687.800 1511.920 1688.060 ;
        RECT 1335.020 20.440 1335.280 20.700 ;
        RECT 1338.240 20.440 1338.500 20.700 ;
      LAYER met2 ;
        RECT 1511.650 1700.000 1511.930 1704.000 ;
        RECT 1511.720 1688.090 1511.860 1700.000 ;
        RECT 1338.240 1687.770 1338.500 1688.090 ;
        RECT 1511.660 1687.770 1511.920 1688.090 ;
        RECT 1338.300 20.730 1338.440 1687.770 ;
        RECT 1335.020 20.410 1335.280 20.730 ;
        RECT 1338.240 20.410 1338.500 20.730 ;
        RECT 1335.080 2.400 1335.220 20.410 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1334.070 1642.440 1334.390 1642.500 ;
        RECT 1336.830 1642.440 1337.150 1642.500 ;
        RECT 1334.070 1642.300 1337.150 1642.440 ;
        RECT 1334.070 1642.240 1334.390 1642.300 ;
        RECT 1336.830 1642.240 1337.150 1642.300 ;
        RECT 696.510 1590.760 696.830 1590.820 ;
        RECT 1334.070 1590.760 1334.390 1590.820 ;
        RECT 696.510 1590.620 1334.390 1590.760 ;
        RECT 696.510 1590.560 696.830 1590.620 ;
        RECT 1334.070 1590.560 1334.390 1590.620 ;
        RECT 692.370 2.960 692.690 3.020 ;
        RECT 696.510 2.960 696.830 3.020 ;
        RECT 692.370 2.820 696.830 2.960 ;
        RECT 692.370 2.760 692.690 2.820 ;
        RECT 696.510 2.760 696.830 2.820 ;
      LAYER via ;
        RECT 1334.100 1642.240 1334.360 1642.500 ;
        RECT 1336.860 1642.240 1337.120 1642.500 ;
        RECT 696.540 1590.560 696.800 1590.820 ;
        RECT 1334.100 1590.560 1334.360 1590.820 ;
        RECT 692.400 2.760 692.660 3.020 ;
        RECT 696.540 2.760 696.800 3.020 ;
      LAYER met2 ;
        RECT 1337.310 1700.410 1337.590 1704.000 ;
        RECT 1336.920 1700.270 1337.590 1700.410 ;
        RECT 1336.920 1642.530 1337.060 1700.270 ;
        RECT 1337.310 1700.000 1337.590 1700.270 ;
        RECT 1334.100 1642.210 1334.360 1642.530 ;
        RECT 1336.860 1642.210 1337.120 1642.530 ;
        RECT 1334.160 1590.850 1334.300 1642.210 ;
        RECT 696.540 1590.530 696.800 1590.850 ;
        RECT 1334.100 1590.530 1334.360 1590.850 ;
        RECT 696.600 3.050 696.740 1590.530 ;
        RECT 692.400 2.730 692.660 3.050 ;
        RECT 696.540 2.730 696.800 3.050 ;
        RECT 692.460 2.400 692.600 2.730 ;
        RECT 692.250 -4.800 692.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 0.300 ;
=======
      LAYER li1 ;
        RECT 1484.565 17.425 1484.735 18.955 ;
      LAYER mcon ;
        RECT 1484.565 18.785 1484.735 18.955 ;
      LAYER met1 ;
        RECT 1512.090 1678.140 1512.410 1678.200 ;
        RECT 1515.310 1678.140 1515.630 1678.200 ;
        RECT 1512.090 1678.000 1515.630 1678.140 ;
        RECT 1512.090 1677.940 1512.410 1678.000 ;
        RECT 1515.310 1677.940 1515.630 1678.000 ;
        RECT 1352.470 18.940 1352.790 19.000 ;
        RECT 1484.505 18.940 1484.795 18.985 ;
        RECT 1352.470 18.800 1484.795 18.940 ;
        RECT 1352.470 18.740 1352.790 18.800 ;
        RECT 1484.505 18.755 1484.795 18.800 ;
        RECT 1512.090 17.920 1512.410 17.980 ;
        RECT 1485.960 17.780 1512.410 17.920 ;
        RECT 1484.505 17.580 1484.795 17.625 ;
        RECT 1485.960 17.580 1486.100 17.780 ;
        RECT 1512.090 17.720 1512.410 17.780 ;
        RECT 1484.505 17.440 1486.100 17.580 ;
        RECT 1484.505 17.395 1484.795 17.440 ;
      LAYER via ;
        RECT 1512.120 1677.940 1512.380 1678.200 ;
        RECT 1515.340 1677.940 1515.600 1678.200 ;
        RECT 1352.500 18.740 1352.760 19.000 ;
        RECT 1512.120 17.720 1512.380 17.980 ;
      LAYER met2 ;
        RECT 1516.250 1700.410 1516.530 1704.000 ;
        RECT 1515.400 1700.270 1516.530 1700.410 ;
        RECT 1515.400 1678.230 1515.540 1700.270 ;
        RECT 1516.250 1700.000 1516.530 1700.270 ;
        RECT 1512.120 1677.910 1512.380 1678.230 ;
        RECT 1515.340 1677.910 1515.600 1678.230 ;
        RECT 1352.500 18.710 1352.760 19.030 ;
        RECT 1352.560 2.400 1352.700 18.710 ;
        RECT 1512.180 18.010 1512.320 1677.910 ;
        RECT 1512.120 17.690 1512.380 18.010 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1393.960 20.500 1512.780 20.640 ;
        RECT 1370.410 20.300 1370.730 20.360 ;
        RECT 1393.960 20.300 1394.100 20.500 ;
        RECT 1370.410 20.160 1394.100 20.300 ;
        RECT 1512.640 20.300 1512.780 20.500 ;
        RECT 1519.450 20.300 1519.770 20.360 ;
        RECT 1512.640 20.160 1519.770 20.300 ;
        RECT 1370.410 20.100 1370.730 20.160 ;
        RECT 1519.450 20.100 1519.770 20.160 ;
      LAYER via ;
        RECT 1370.440 20.100 1370.700 20.360 ;
        RECT 1519.480 20.100 1519.740 20.360 ;
      LAYER met2 ;
        RECT 1519.930 1700.410 1520.210 1704.000 ;
        RECT 1519.540 1700.270 1520.210 1700.410 ;
        RECT 1519.540 20.390 1519.680 1700.270 ;
        RECT 1519.930 1700.000 1520.210 1700.270 ;
        RECT 1370.440 20.070 1370.700 20.390 ;
        RECT 1519.480 20.070 1519.740 20.390 ;
        RECT 1370.500 2.400 1370.640 20.070 ;
=======
      LAYER li1 ;
        RECT 1485.945 17.595 1486.115 19.295 ;
        RECT 1485.945 17.425 1486.575 17.595 ;
      LAYER mcon ;
        RECT 1485.945 19.125 1486.115 19.295 ;
        RECT 1486.405 17.425 1486.575 17.595 ;
      LAYER met1 ;
        RECT 1370.410 19.280 1370.730 19.340 ;
        RECT 1485.885 19.280 1486.175 19.325 ;
        RECT 1370.410 19.140 1486.175 19.280 ;
        RECT 1370.410 19.080 1370.730 19.140 ;
        RECT 1485.885 19.095 1486.175 19.140 ;
        RECT 1486.345 17.580 1486.635 17.625 ;
        RECT 1519.910 17.580 1520.230 17.640 ;
        RECT 1486.345 17.440 1520.230 17.580 ;
        RECT 1486.345 17.395 1486.635 17.440 ;
        RECT 1519.910 17.380 1520.230 17.440 ;
      LAYER via ;
        RECT 1370.440 19.080 1370.700 19.340 ;
        RECT 1519.940 17.380 1520.200 17.640 ;
      LAYER met2 ;
        RECT 1521.310 1700.410 1521.590 1704.000 ;
        RECT 1520.000 1700.270 1521.590 1700.410 ;
        RECT 1370.440 19.050 1370.700 19.370 ;
        RECT 1370.500 2.400 1370.640 19.050 ;
        RECT 1520.000 17.670 1520.140 1700.270 ;
        RECT 1521.310 1700.000 1521.590 1700.270 ;
        RECT 1519.940 17.350 1520.200 17.670 ;
>>>>>>> re-updated local openlane
        RECT 1370.290 -4.800 1370.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 0.300 ;
=======
      LAYER li1 ;
        RECT 1404.065 1241.765 1404.235 1256.215 ;
      LAYER mcon ;
        RECT 1404.065 1256.045 1404.235 1256.215 ;
      LAYER met1 ;
        RECT 1405.830 1689.700 1406.150 1689.760 ;
        RECT 1525.890 1689.700 1526.210 1689.760 ;
        RECT 1405.830 1689.560 1526.210 1689.700 ;
        RECT 1405.830 1689.500 1406.150 1689.560 ;
        RECT 1525.890 1689.500 1526.210 1689.560 ;
        RECT 1403.990 1628.640 1404.310 1628.900 ;
        RECT 1404.080 1628.220 1404.220 1628.640 ;
        RECT 1403.990 1627.960 1404.310 1628.220 ;
        RECT 1403.990 1256.200 1404.310 1256.260 ;
        RECT 1403.795 1256.060 1404.310 1256.200 ;
        RECT 1403.990 1256.000 1404.310 1256.060 ;
        RECT 1403.990 1241.920 1404.310 1241.980 ;
        RECT 1403.795 1241.780 1404.310 1241.920 ;
        RECT 1403.990 1241.720 1404.310 1241.780 ;
        RECT 1388.350 20.300 1388.670 20.360 ;
        RECT 1403.990 20.300 1404.310 20.360 ;
        RECT 1388.350 20.160 1404.310 20.300 ;
        RECT 1388.350 20.100 1388.670 20.160 ;
        RECT 1403.990 20.100 1404.310 20.160 ;
      LAYER via ;
        RECT 1405.860 1689.500 1406.120 1689.760 ;
        RECT 1525.920 1689.500 1526.180 1689.760 ;
        RECT 1404.020 1628.640 1404.280 1628.900 ;
        RECT 1404.020 1627.960 1404.280 1628.220 ;
        RECT 1404.020 1256.000 1404.280 1256.260 ;
        RECT 1404.020 1241.720 1404.280 1241.980 ;
        RECT 1388.380 20.100 1388.640 20.360 ;
        RECT 1404.020 20.100 1404.280 20.360 ;
      LAYER met2 ;
        RECT 1525.910 1700.000 1526.190 1704.000 ;
        RECT 1525.980 1689.790 1526.120 1700.000 ;
        RECT 1405.860 1689.470 1406.120 1689.790 ;
        RECT 1525.920 1689.470 1526.180 1689.790 ;
        RECT 1405.920 1673.210 1406.060 1689.470 ;
        RECT 1404.080 1673.070 1406.060 1673.210 ;
        RECT 1404.080 1628.930 1404.220 1673.070 ;
        RECT 1404.020 1628.610 1404.280 1628.930 ;
        RECT 1404.020 1627.930 1404.280 1628.250 ;
        RECT 1404.080 1256.290 1404.220 1627.930 ;
        RECT 1404.020 1255.970 1404.280 1256.290 ;
        RECT 1404.020 1241.690 1404.280 1242.010 ;
        RECT 1404.080 20.390 1404.220 1241.690 ;
        RECT 1388.380 20.070 1388.640 20.390 ;
        RECT 1404.020 20.070 1404.280 20.390 ;
        RECT 1388.440 2.400 1388.580 20.070 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 0.300 ;
=======
      LAYER li1 ;
        RECT 1479.505 1684.445 1479.675 1685.635 ;
      LAYER mcon ;
        RECT 1479.505 1685.465 1479.675 1685.635 ;
      LAYER met1 ;
        RECT 1407.210 1685.620 1407.530 1685.680 ;
        RECT 1479.445 1685.620 1479.735 1685.665 ;
        RECT 1407.210 1685.480 1479.735 1685.620 ;
        RECT 1407.210 1685.420 1407.530 1685.480 ;
        RECT 1479.445 1685.435 1479.735 1685.480 ;
        RECT 1479.445 1684.600 1479.735 1684.645 ;
        RECT 1529.570 1684.600 1529.890 1684.660 ;
        RECT 1479.445 1684.460 1529.890 1684.600 ;
        RECT 1479.445 1684.415 1479.735 1684.460 ;
        RECT 1529.570 1684.400 1529.890 1684.460 ;
        RECT 1406.290 2.960 1406.610 3.020 ;
        RECT 1407.210 2.960 1407.530 3.020 ;
        RECT 1406.290 2.820 1407.530 2.960 ;
        RECT 1406.290 2.760 1406.610 2.820 ;
        RECT 1407.210 2.760 1407.530 2.820 ;
      LAYER via ;
        RECT 1407.240 1685.420 1407.500 1685.680 ;
        RECT 1529.600 1684.400 1529.860 1684.660 ;
        RECT 1406.320 2.760 1406.580 3.020 ;
        RECT 1407.240 2.760 1407.500 3.020 ;
      LAYER met2 ;
        RECT 1529.590 1700.000 1529.870 1704.000 ;
        RECT 1407.240 1685.390 1407.500 1685.710 ;
        RECT 1407.300 3.050 1407.440 1685.390 ;
        RECT 1529.660 1684.690 1529.800 1700.000 ;
        RECT 1529.600 1684.370 1529.860 1684.690 ;
        RECT 1406.320 2.730 1406.580 3.050 ;
        RECT 1407.240 2.730 1407.500 3.050 ;
        RECT 1406.380 2.400 1406.520 2.730 ;
=======
      LAYER met1 ;
        RECT 1526.350 20.640 1526.670 20.700 ;
        RECT 1486.880 20.500 1526.670 20.640 ;
        RECT 1406.290 20.300 1406.610 20.360 ;
        RECT 1486.880 20.300 1487.020 20.500 ;
        RECT 1526.350 20.440 1526.670 20.500 ;
        RECT 1406.290 20.160 1487.020 20.300 ;
        RECT 1406.290 20.100 1406.610 20.160 ;
      LAYER via ;
        RECT 1406.320 20.100 1406.580 20.360 ;
        RECT 1526.380 20.440 1526.640 20.700 ;
      LAYER met2 ;
        RECT 1530.970 1700.410 1531.250 1704.000 ;
        RECT 1529.660 1700.270 1531.250 1700.410 ;
        RECT 1529.660 1678.650 1529.800 1700.270 ;
        RECT 1530.970 1700.000 1531.250 1700.270 ;
        RECT 1526.440 1678.510 1529.800 1678.650 ;
        RECT 1526.440 20.730 1526.580 1678.510 ;
        RECT 1526.380 20.410 1526.640 20.730 ;
        RECT 1406.320 20.070 1406.580 20.390 ;
        RECT 1406.380 2.400 1406.520 20.070 ;
>>>>>>> re-updated local openlane
        RECT 1406.170 -4.800 1406.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 0.300 ;
=======
=======
      LAYER li1 ;
        RECT 1452.825 16.065 1452.995 20.655 ;
        RECT 1486.405 20.485 1487.035 20.655 ;
        RECT 1486.865 19.125 1487.035 20.485 ;
      LAYER mcon ;
        RECT 1452.825 20.485 1452.995 20.655 ;
>>>>>>> re-updated local openlane
      LAYER met1 ;
        RECT 1452.765 20.640 1453.055 20.685 ;
        RECT 1486.345 20.640 1486.635 20.685 ;
        RECT 1452.765 20.500 1486.635 20.640 ;
        RECT 1452.765 20.455 1453.055 20.500 ;
        RECT 1486.345 20.455 1486.635 20.500 ;
        RECT 1486.805 19.280 1487.095 19.325 ;
        RECT 1532.790 19.280 1533.110 19.340 ;
        RECT 1486.805 19.140 1533.110 19.280 ;
        RECT 1486.805 19.095 1487.095 19.140 ;
        RECT 1532.790 19.080 1533.110 19.140 ;
        RECT 1423.770 16.220 1424.090 16.280 ;
        RECT 1452.765 16.220 1453.055 16.265 ;
        RECT 1423.770 16.080 1453.055 16.220 ;
        RECT 1423.770 16.020 1424.090 16.080 ;
        RECT 1452.765 16.035 1453.055 16.080 ;
      LAYER via ;
        RECT 1532.820 19.080 1533.080 19.340 ;
        RECT 1423.800 16.020 1424.060 16.280 ;
      LAYER met2 ;
        RECT 1535.570 1700.410 1535.850 1704.000 ;
        RECT 1534.720 1700.270 1535.850 1700.410 ;
        RECT 1534.720 1677.970 1534.860 1700.270 ;
        RECT 1535.570 1700.000 1535.850 1700.270 ;
        RECT 1532.880 1677.830 1534.860 1677.970 ;
        RECT 1532.880 19.370 1533.020 1677.830 ;
        RECT 1532.820 19.050 1533.080 19.370 ;
        RECT 1423.800 15.990 1424.060 16.310 ;
        RECT 1423.860 2.400 1424.000 15.990 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 0.300 ;
=======
      LAYER met1 ;
        RECT 1441.710 1690.040 1442.030 1690.100 ;
        RECT 1540.610 1690.040 1540.930 1690.100 ;
        RECT 1441.710 1689.900 1540.930 1690.040 ;
        RECT 1441.710 1689.840 1442.030 1689.900 ;
        RECT 1540.610 1689.840 1540.930 1689.900 ;
      LAYER via ;
        RECT 1441.740 1689.840 1442.000 1690.100 ;
        RECT 1540.640 1689.840 1540.900 1690.100 ;
      LAYER met2 ;
        RECT 1540.630 1700.000 1540.910 1704.000 ;
        RECT 1540.700 1690.130 1540.840 1700.000 ;
        RECT 1441.740 1689.810 1442.000 1690.130 ;
        RECT 1540.640 1689.810 1540.900 1690.130 ;
        RECT 1441.800 2.400 1441.940 1689.810 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1539.230 1678.480 1539.550 1678.540 ;
        RECT 1544.290 1678.480 1544.610 1678.540 ;
        RECT 1539.230 1678.340 1544.610 1678.480 ;
        RECT 1539.230 1678.280 1539.550 1678.340 ;
        RECT 1544.290 1678.280 1544.610 1678.340 ;
        RECT 1511.630 17.240 1511.950 17.300 ;
        RECT 1539.230 17.240 1539.550 17.300 ;
        RECT 1511.630 17.100 1539.550 17.240 ;
        RECT 1511.630 17.040 1511.950 17.100 ;
        RECT 1539.230 17.040 1539.550 17.100 ;
        RECT 1459.650 15.880 1459.970 15.940 ;
        RECT 1510.250 15.880 1510.570 15.940 ;
        RECT 1459.650 15.740 1510.570 15.880 ;
        RECT 1459.650 15.680 1459.970 15.740 ;
        RECT 1510.250 15.680 1510.570 15.740 ;
      LAYER via ;
        RECT 1539.260 1678.280 1539.520 1678.540 ;
        RECT 1544.320 1678.280 1544.580 1678.540 ;
        RECT 1511.660 17.040 1511.920 17.300 ;
        RECT 1539.260 17.040 1539.520 17.300 ;
        RECT 1459.680 15.680 1459.940 15.940 ;
        RECT 1510.280 15.680 1510.540 15.940 ;
      LAYER met2 ;
        RECT 1545.230 1700.410 1545.510 1704.000 ;
        RECT 1544.380 1700.270 1545.510 1700.410 ;
        RECT 1544.380 1678.570 1544.520 1700.270 ;
        RECT 1545.230 1700.000 1545.510 1700.270 ;
        RECT 1539.260 1678.250 1539.520 1678.570 ;
        RECT 1544.320 1678.250 1544.580 1678.570 ;
        RECT 1539.320 17.330 1539.460 1678.250 ;
        RECT 1511.660 17.010 1511.920 17.330 ;
        RECT 1539.260 17.010 1539.520 17.330 ;
        RECT 1511.720 16.165 1511.860 17.010 ;
        RECT 1459.680 15.650 1459.940 15.970 ;
        RECT 1510.270 15.795 1510.550 16.165 ;
        RECT 1511.650 15.795 1511.930 16.165 ;
        RECT 1510.280 15.650 1510.540 15.795 ;
        RECT 1459.740 2.400 1459.880 15.650 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 1510.270 15.840 1510.550 16.120 ;
        RECT 1511.650 15.840 1511.930 16.120 ;
      LAYER met3 ;
        RECT 1510.245 16.130 1510.575 16.145 ;
        RECT 1511.625 16.130 1511.955 16.145 ;
        RECT 1510.245 15.830 1511.955 16.130 ;
        RECT 1510.245 15.815 1510.575 15.830 ;
        RECT 1511.625 15.815 1511.955 15.830 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1546.130 1678.140 1546.450 1678.200 ;
        RECT 1548.890 1678.140 1549.210 1678.200 ;
        RECT 1546.130 1678.000 1549.210 1678.140 ;
        RECT 1546.130 1677.940 1546.450 1678.000 ;
        RECT 1548.890 1677.940 1549.210 1678.000 ;
        RECT 1546.130 15.540 1546.450 15.600 ;
        RECT 1524.600 15.400 1546.450 15.540 ;
        RECT 1477.590 15.200 1477.910 15.260 ;
        RECT 1524.600 15.200 1524.740 15.400 ;
        RECT 1546.130 15.340 1546.450 15.400 ;
        RECT 1477.590 15.060 1524.740 15.200 ;
        RECT 1477.590 15.000 1477.910 15.060 ;
      LAYER via ;
        RECT 1546.160 1677.940 1546.420 1678.200 ;
        RECT 1548.920 1677.940 1549.180 1678.200 ;
        RECT 1477.620 15.000 1477.880 15.260 ;
        RECT 1546.160 15.340 1546.420 15.600 ;
      LAYER met2 ;
        RECT 1550.290 1700.410 1550.570 1704.000 ;
        RECT 1548.980 1700.270 1550.570 1700.410 ;
        RECT 1548.980 1678.230 1549.120 1700.270 ;
        RECT 1550.290 1700.000 1550.570 1700.270 ;
        RECT 1546.160 1677.910 1546.420 1678.230 ;
        RECT 1548.920 1677.910 1549.180 1678.230 ;
        RECT 1546.220 15.630 1546.360 1677.910 ;
        RECT 1546.160 15.310 1546.420 15.630 ;
        RECT 1477.620 14.970 1477.880 15.290 ;
        RECT 1477.680 2.400 1477.820 14.970 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 0.300 ;
=======
      LAYER li1 ;
        RECT 1514.465 1655.545 1514.635 1687.675 ;
      LAYER mcon ;
        RECT 1514.465 1687.505 1514.635 1687.675 ;
      LAYER met1 ;
        RECT 1514.405 1687.660 1514.695 1687.705 ;
        RECT 1553.490 1687.660 1553.810 1687.720 ;
        RECT 1514.405 1687.520 1553.810 1687.660 ;
        RECT 1514.405 1687.475 1514.695 1687.520 ;
        RECT 1553.490 1687.460 1553.810 1687.520 ;
        RECT 1514.390 1655.700 1514.710 1655.760 ;
        RECT 1514.195 1655.560 1514.710 1655.700 ;
        RECT 1514.390 1655.500 1514.710 1655.560 ;
        RECT 1495.530 16.220 1495.850 16.280 ;
        RECT 1514.390 16.220 1514.710 16.280 ;
        RECT 1495.530 16.080 1514.710 16.220 ;
        RECT 1495.530 16.020 1495.850 16.080 ;
        RECT 1514.390 16.020 1514.710 16.080 ;
      LAYER via ;
        RECT 1553.520 1687.460 1553.780 1687.720 ;
        RECT 1514.420 1655.500 1514.680 1655.760 ;
        RECT 1495.560 16.020 1495.820 16.280 ;
        RECT 1514.420 16.020 1514.680 16.280 ;
      LAYER met2 ;
        RECT 1553.510 1700.000 1553.790 1704.000 ;
        RECT 1553.580 1687.750 1553.720 1700.000 ;
        RECT 1553.520 1687.430 1553.780 1687.750 ;
        RECT 1514.420 1655.470 1514.680 1655.790 ;
        RECT 1514.480 16.310 1514.620 1655.470 ;
        RECT 1495.560 15.990 1495.820 16.310 ;
        RECT 1514.420 15.990 1514.680 16.310 ;
        RECT 1495.620 2.400 1495.760 15.990 ;
=======
      LAYER met1 ;
        RECT 1555.330 1689.360 1555.650 1689.420 ;
        RECT 1539.320 1689.220 1555.650 1689.360 ;
        RECT 1522.210 1689.020 1522.530 1689.080 ;
        RECT 1539.320 1689.020 1539.460 1689.220 ;
        RECT 1555.330 1689.160 1555.650 1689.220 ;
        RECT 1522.210 1688.880 1539.460 1689.020 ;
        RECT 1522.210 1688.820 1522.530 1688.880 ;
        RECT 1495.530 14.860 1495.850 14.920 ;
        RECT 1521.750 14.860 1522.070 14.920 ;
        RECT 1495.530 14.720 1522.070 14.860 ;
        RECT 1495.530 14.660 1495.850 14.720 ;
        RECT 1521.750 14.660 1522.070 14.720 ;
      LAYER via ;
        RECT 1522.240 1688.820 1522.500 1689.080 ;
        RECT 1555.360 1689.160 1555.620 1689.420 ;
        RECT 1495.560 14.660 1495.820 14.920 ;
        RECT 1521.780 14.660 1522.040 14.920 ;
      LAYER met2 ;
        RECT 1555.350 1700.000 1555.630 1704.000 ;
        RECT 1555.420 1689.450 1555.560 1700.000 ;
        RECT 1555.360 1689.130 1555.620 1689.450 ;
        RECT 1522.240 1688.790 1522.500 1689.110 ;
        RECT 1522.300 1677.290 1522.440 1688.790 ;
        RECT 1521.840 1677.150 1522.440 1677.290 ;
        RECT 1521.840 14.950 1521.980 1677.150 ;
        RECT 1495.560 14.630 1495.820 14.950 ;
        RECT 1521.780 14.630 1522.040 14.950 ;
        RECT 1495.620 2.400 1495.760 14.630 ;
>>>>>>> re-updated local openlane
        RECT 1495.410 -4.800 1495.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1530.030 1687.660 1530.350 1687.720 ;
        RECT 1559.930 1687.660 1560.250 1687.720 ;
        RECT 1530.030 1687.520 1560.250 1687.660 ;
        RECT 1530.030 1687.460 1530.350 1687.520 ;
        RECT 1559.930 1687.460 1560.250 1687.520 ;
        RECT 1513.010 19.960 1513.330 20.020 ;
        RECT 1528.190 19.960 1528.510 20.020 ;
        RECT 1513.010 19.820 1528.510 19.960 ;
        RECT 1513.010 19.760 1513.330 19.820 ;
        RECT 1528.190 19.760 1528.510 19.820 ;
      LAYER via ;
        RECT 1530.060 1687.460 1530.320 1687.720 ;
        RECT 1559.960 1687.460 1560.220 1687.720 ;
        RECT 1513.040 19.760 1513.300 20.020 ;
        RECT 1528.220 19.760 1528.480 20.020 ;
      LAYER met2 ;
        RECT 1559.950 1700.000 1560.230 1704.000 ;
        RECT 1560.020 1687.750 1560.160 1700.000 ;
        RECT 1530.060 1687.430 1530.320 1687.750 ;
        RECT 1559.960 1687.430 1560.220 1687.750 ;
        RECT 1530.120 1671.850 1530.260 1687.430 ;
        RECT 1528.280 1671.710 1530.260 1671.850 ;
        RECT 1528.280 20.050 1528.420 1671.710 ;
        RECT 1513.040 19.730 1513.300 20.050 ;
        RECT 1528.220 19.730 1528.480 20.050 ;
        RECT 1513.100 2.400 1513.240 19.730 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1339.590 1693.440 1339.910 1693.500 ;
        RECT 1342.350 1693.440 1342.670 1693.500 ;
        RECT 1339.590 1693.300 1342.670 1693.440 ;
        RECT 1339.590 1693.240 1339.910 1693.300 ;
        RECT 1342.350 1693.240 1342.670 1693.300 ;
        RECT 709.850 1583.620 710.170 1583.680 ;
        RECT 1339.590 1583.620 1339.910 1583.680 ;
        RECT 709.850 1583.480 1339.910 1583.620 ;
        RECT 709.850 1583.420 710.170 1583.480 ;
        RECT 1339.590 1583.420 1339.910 1583.480 ;
      LAYER via ;
        RECT 1339.620 1693.240 1339.880 1693.500 ;
        RECT 1342.380 1693.240 1342.640 1693.500 ;
        RECT 709.880 1583.420 710.140 1583.680 ;
        RECT 1339.620 1583.420 1339.880 1583.680 ;
      LAYER met2 ;
        RECT 1342.370 1700.000 1342.650 1704.000 ;
        RECT 1342.440 1693.530 1342.580 1700.000 ;
        RECT 1339.620 1693.210 1339.880 1693.530 ;
        RECT 1342.380 1693.210 1342.640 1693.530 ;
        RECT 1339.680 1583.710 1339.820 1693.210 ;
        RECT 709.880 1583.390 710.140 1583.710 ;
        RECT 1339.620 1583.390 1339.880 1583.710 ;
        RECT 709.940 17.410 710.080 1583.390 ;
        RECT 709.940 17.270 710.540 17.410 ;
        RECT 710.400 2.400 710.540 17.270 ;
        RECT 710.190 -4.800 710.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1560.390 1667.600 1560.710 1667.660 ;
        RECT 1563.610 1667.600 1563.930 1667.660 ;
        RECT 1560.390 1667.460 1563.930 1667.600 ;
        RECT 1560.390 1667.400 1560.710 1667.460 ;
        RECT 1563.610 1667.400 1563.930 1667.460 ;
        RECT 1530.950 19.620 1531.270 19.680 ;
        RECT 1560.390 19.620 1560.710 19.680 ;
        RECT 1530.950 19.480 1560.710 19.620 ;
        RECT 1530.950 19.420 1531.270 19.480 ;
        RECT 1560.390 19.420 1560.710 19.480 ;
      LAYER via ;
        RECT 1560.420 1667.400 1560.680 1667.660 ;
        RECT 1563.640 1667.400 1563.900 1667.660 ;
        RECT 1530.980 19.420 1531.240 19.680 ;
        RECT 1560.420 19.420 1560.680 19.680 ;
      LAYER met2 ;
        RECT 1565.010 1700.410 1565.290 1704.000 ;
        RECT 1563.700 1700.270 1565.290 1700.410 ;
        RECT 1563.700 1667.690 1563.840 1700.270 ;
        RECT 1565.010 1700.000 1565.290 1700.270 ;
        RECT 1560.420 1667.370 1560.680 1667.690 ;
        RECT 1563.640 1667.370 1563.900 1667.690 ;
        RECT 1560.480 19.710 1560.620 1667.370 ;
        RECT 1530.980 19.390 1531.240 19.710 ;
        RECT 1560.420 19.390 1560.680 19.710 ;
        RECT 1531.040 2.400 1531.180 19.390 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1552.110 1689.020 1552.430 1689.080 ;
        RECT 1569.590 1689.020 1569.910 1689.080 ;
        RECT 1552.110 1688.880 1569.910 1689.020 ;
        RECT 1552.110 1688.820 1552.430 1688.880 ;
        RECT 1569.590 1688.820 1569.910 1688.880 ;
        RECT 1548.890 20.640 1549.210 20.700 ;
        RECT 1552.110 20.640 1552.430 20.700 ;
        RECT 1548.890 20.500 1552.430 20.640 ;
        RECT 1548.890 20.440 1549.210 20.500 ;
        RECT 1552.110 20.440 1552.430 20.500 ;
      LAYER via ;
        RECT 1552.140 1688.820 1552.400 1689.080 ;
        RECT 1569.620 1688.820 1569.880 1689.080 ;
        RECT 1548.920 20.440 1549.180 20.700 ;
        RECT 1552.140 20.440 1552.400 20.700 ;
      LAYER met2 ;
        RECT 1569.610 1700.000 1569.890 1704.000 ;
        RECT 1569.680 1689.110 1569.820 1700.000 ;
        RECT 1552.140 1688.790 1552.400 1689.110 ;
        RECT 1569.620 1688.790 1569.880 1689.110 ;
        RECT 1552.200 20.730 1552.340 1688.790 ;
        RECT 1548.920 20.410 1549.180 20.730 ;
        RECT 1552.140 20.410 1552.400 20.730 ;
        RECT 1548.980 2.400 1549.120 20.410 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1566.830 15.200 1567.150 15.260 ;
        RECT 1573.270 15.200 1573.590 15.260 ;
        RECT 1566.830 15.060 1573.590 15.200 ;
        RECT 1566.830 15.000 1567.150 15.060 ;
        RECT 1573.270 15.000 1573.590 15.060 ;
      LAYER via ;
        RECT 1566.860 15.000 1567.120 15.260 ;
        RECT 1573.300 15.000 1573.560 15.260 ;
      LAYER met2 ;
        RECT 1574.670 1700.410 1574.950 1704.000 ;
        RECT 1573.360 1700.270 1574.950 1700.410 ;
        RECT 1573.360 15.290 1573.500 1700.270 ;
        RECT 1574.670 1700.000 1574.950 1700.270 ;
        RECT 1566.860 14.970 1567.120 15.290 ;
        RECT 1573.300 14.970 1573.560 15.290 ;
        RECT 1566.920 2.400 1567.060 14.970 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 0.300 ;
=======
      LAYER met1 ;
        RECT 1579.250 1683.920 1579.570 1683.980 ;
        RECT 1582.010 1683.920 1582.330 1683.980 ;
        RECT 1579.250 1683.780 1582.330 1683.920 ;
        RECT 1579.250 1683.720 1579.570 1683.780 ;
        RECT 1582.010 1683.720 1582.330 1683.780 ;
        RECT 1582.010 2.960 1582.330 3.020 ;
        RECT 1584.770 2.960 1585.090 3.020 ;
        RECT 1582.010 2.820 1585.090 2.960 ;
        RECT 1582.010 2.760 1582.330 2.820 ;
        RECT 1584.770 2.760 1585.090 2.820 ;
      LAYER via ;
        RECT 1579.280 1683.720 1579.540 1683.980 ;
        RECT 1582.040 1683.720 1582.300 1683.980 ;
        RECT 1582.040 2.760 1582.300 3.020 ;
        RECT 1584.800 2.760 1585.060 3.020 ;
      LAYER met2 ;
        RECT 1579.270 1700.000 1579.550 1704.000 ;
        RECT 1579.340 1684.010 1579.480 1700.000 ;
        RECT 1579.280 1683.690 1579.540 1684.010 ;
        RECT 1582.040 1683.690 1582.300 1684.010 ;
        RECT 1582.100 3.050 1582.240 1683.690 ;
        RECT 1582.040 2.730 1582.300 3.050 ;
        RECT 1584.800 2.730 1585.060 3.050 ;
        RECT 1584.860 2.400 1585.000 2.730 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1584.310 1683.920 1584.630 1683.980 ;
        RECT 1586.610 1683.920 1586.930 1683.980 ;
        RECT 1584.310 1683.780 1586.930 1683.920 ;
        RECT 1584.310 1683.720 1584.630 1683.780 ;
        RECT 1586.610 1683.720 1586.930 1683.780 ;
        RECT 1586.610 20.300 1586.930 20.360 ;
        RECT 1602.250 20.300 1602.570 20.360 ;
        RECT 1586.610 20.160 1602.570 20.300 ;
        RECT 1586.610 20.100 1586.930 20.160 ;
        RECT 1602.250 20.100 1602.570 20.160 ;
      LAYER via ;
        RECT 1584.340 1683.720 1584.600 1683.980 ;
        RECT 1586.640 1683.720 1586.900 1683.980 ;
        RECT 1586.640 20.100 1586.900 20.360 ;
        RECT 1602.280 20.100 1602.540 20.360 ;
      LAYER met2 ;
        RECT 1584.330 1700.000 1584.610 1704.000 ;
        RECT 1584.400 1684.010 1584.540 1700.000 ;
        RECT 1584.340 1683.690 1584.600 1684.010 ;
        RECT 1586.640 1683.690 1586.900 1684.010 ;
        RECT 1586.700 20.390 1586.840 1683.690 ;
        RECT 1586.640 20.070 1586.900 20.390 ;
        RECT 1602.280 20.070 1602.540 20.390 ;
        RECT 1602.340 2.400 1602.480 20.070 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 0.300 ;
=======
      LAYER met1 ;
        RECT 1588.910 1683.920 1589.230 1683.980 ;
        RECT 1597.190 1683.920 1597.510 1683.980 ;
        RECT 1588.910 1683.780 1597.510 1683.920 ;
        RECT 1588.910 1683.720 1589.230 1683.780 ;
        RECT 1597.190 1683.720 1597.510 1683.780 ;
        RECT 1597.190 17.920 1597.510 17.980 ;
        RECT 1620.190 17.920 1620.510 17.980 ;
        RECT 1597.190 17.780 1620.510 17.920 ;
        RECT 1597.190 17.720 1597.510 17.780 ;
        RECT 1620.190 17.720 1620.510 17.780 ;
      LAYER via ;
        RECT 1588.940 1683.720 1589.200 1683.980 ;
        RECT 1597.220 1683.720 1597.480 1683.980 ;
        RECT 1597.220 17.720 1597.480 17.980 ;
        RECT 1620.220 17.720 1620.480 17.980 ;
      LAYER met2 ;
        RECT 1588.930 1700.000 1589.210 1704.000 ;
        RECT 1589.000 1684.010 1589.140 1700.000 ;
        RECT 1588.940 1683.690 1589.200 1684.010 ;
        RECT 1597.220 1683.690 1597.480 1684.010 ;
        RECT 1597.280 18.010 1597.420 1683.690 ;
        RECT 1597.220 17.690 1597.480 18.010 ;
        RECT 1620.220 17.690 1620.480 18.010 ;
        RECT 1620.280 2.400 1620.420 17.690 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1593.970 1684.940 1594.290 1685.000 ;
        RECT 1604.090 1684.940 1604.410 1685.000 ;
        RECT 1593.970 1684.800 1604.410 1684.940 ;
        RECT 1593.970 1684.740 1594.290 1684.800 ;
        RECT 1604.090 1684.740 1604.410 1684.800 ;
        RECT 1604.090 19.280 1604.410 19.340 ;
        RECT 1638.130 19.280 1638.450 19.340 ;
        RECT 1604.090 19.140 1638.450 19.280 ;
        RECT 1604.090 19.080 1604.410 19.140 ;
        RECT 1638.130 19.080 1638.450 19.140 ;
      LAYER via ;
        RECT 1594.000 1684.740 1594.260 1685.000 ;
        RECT 1604.120 1684.740 1604.380 1685.000 ;
        RECT 1604.120 19.080 1604.380 19.340 ;
        RECT 1638.160 19.080 1638.420 19.340 ;
      LAYER met2 ;
        RECT 1593.990 1700.000 1594.270 1704.000 ;
        RECT 1594.060 1685.030 1594.200 1700.000 ;
        RECT 1594.000 1684.710 1594.260 1685.030 ;
        RECT 1604.120 1684.710 1604.380 1685.030 ;
        RECT 1604.180 19.370 1604.320 1684.710 ;
        RECT 1604.120 19.050 1604.380 19.370 ;
        RECT 1638.160 19.050 1638.420 19.370 ;
        RECT 1638.220 2.400 1638.360 19.050 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 0.300 ;
=======
      LAYER li1 ;
        RECT 1632.225 17.765 1632.395 19.635 ;
      LAYER mcon ;
        RECT 1632.225 19.465 1632.395 19.635 ;
      LAYER met1 ;
        RECT 1598.570 1683.920 1598.890 1683.980 ;
        RECT 1600.410 1683.920 1600.730 1683.980 ;
        RECT 1598.570 1683.780 1600.730 1683.920 ;
        RECT 1598.570 1683.720 1598.890 1683.780 ;
        RECT 1600.410 1683.720 1600.730 1683.780 ;
        RECT 1600.410 19.620 1600.730 19.680 ;
        RECT 1632.165 19.620 1632.455 19.665 ;
        RECT 1600.410 19.480 1632.455 19.620 ;
        RECT 1600.410 19.420 1600.730 19.480 ;
        RECT 1632.165 19.435 1632.455 19.480 ;
        RECT 1632.165 17.920 1632.455 17.965 ;
        RECT 1656.070 17.920 1656.390 17.980 ;
        RECT 1632.165 17.780 1656.390 17.920 ;
        RECT 1632.165 17.735 1632.455 17.780 ;
        RECT 1656.070 17.720 1656.390 17.780 ;
      LAYER via ;
        RECT 1598.600 1683.720 1598.860 1683.980 ;
        RECT 1600.440 1683.720 1600.700 1683.980 ;
        RECT 1600.440 19.420 1600.700 19.680 ;
        RECT 1656.100 17.720 1656.360 17.980 ;
      LAYER met2 ;
        RECT 1598.590 1700.000 1598.870 1704.000 ;
        RECT 1598.660 1684.010 1598.800 1700.000 ;
        RECT 1598.600 1683.690 1598.860 1684.010 ;
        RECT 1600.440 1683.690 1600.700 1684.010 ;
        RECT 1600.500 19.710 1600.640 1683.690 ;
        RECT 1600.440 19.390 1600.700 19.710 ;
        RECT 1656.100 17.690 1656.360 18.010 ;
        RECT 1656.160 2.400 1656.300 17.690 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 0.300 ;
=======
      LAYER li1 ;
        RECT 1628.545 1686.485 1628.715 1688.015 ;
      LAYER mcon ;
        RECT 1628.545 1687.845 1628.715 1688.015 ;
      LAYER met1 ;
        RECT 1601.790 1688.000 1602.110 1688.060 ;
        RECT 1628.485 1688.000 1628.775 1688.045 ;
        RECT 1601.790 1687.860 1628.775 1688.000 ;
        RECT 1601.790 1687.800 1602.110 1687.860 ;
        RECT 1628.485 1687.815 1628.775 1687.860 ;
        RECT 1628.485 1686.640 1628.775 1686.685 ;
        RECT 1666.190 1686.640 1666.510 1686.700 ;
        RECT 1628.485 1686.500 1666.510 1686.640 ;
        RECT 1628.485 1686.455 1628.775 1686.500 ;
        RECT 1666.190 1686.440 1666.510 1686.500 ;
        RECT 1666.190 17.580 1666.510 17.640 ;
        RECT 1673.550 17.580 1673.870 17.640 ;
        RECT 1666.190 17.440 1673.870 17.580 ;
        RECT 1666.190 17.380 1666.510 17.440 ;
        RECT 1673.550 17.380 1673.870 17.440 ;
      LAYER via ;
        RECT 1601.820 1687.800 1602.080 1688.060 ;
        RECT 1666.220 1686.440 1666.480 1686.700 ;
        RECT 1666.220 17.380 1666.480 17.640 ;
        RECT 1673.580 17.380 1673.840 17.640 ;
=======
      LAYER met1 ;
        RECT 1603.630 1683.920 1603.950 1683.980 ;
        RECT 1606.850 1683.920 1607.170 1683.980 ;
        RECT 1603.630 1683.780 1607.170 1683.920 ;
        RECT 1603.630 1683.720 1603.950 1683.780 ;
        RECT 1606.850 1683.720 1607.170 1683.780 ;
        RECT 1606.850 17.240 1607.170 17.300 ;
        RECT 1673.550 17.240 1673.870 17.300 ;
        RECT 1606.850 17.100 1673.870 17.240 ;
        RECT 1606.850 17.040 1607.170 17.100 ;
        RECT 1673.550 17.040 1673.870 17.100 ;
      LAYER via ;
        RECT 1603.660 1683.720 1603.920 1683.980 ;
        RECT 1606.880 1683.720 1607.140 1683.980 ;
        RECT 1606.880 17.040 1607.140 17.300 ;
        RECT 1673.580 17.040 1673.840 17.300 ;
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1603.650 1700.000 1603.930 1704.000 ;
        RECT 1603.720 1684.010 1603.860 1700.000 ;
        RECT 1603.660 1683.690 1603.920 1684.010 ;
        RECT 1606.880 1683.690 1607.140 1684.010 ;
        RECT 1606.940 17.330 1607.080 1683.690 ;
        RECT 1606.880 17.010 1607.140 17.330 ;
        RECT 1673.580 17.010 1673.840 17.330 ;
        RECT 1673.640 2.400 1673.780 17.010 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1608.230 1683.920 1608.550 1683.980 ;
        RECT 1614.210 1683.920 1614.530 1683.980 ;
        RECT 1608.230 1683.780 1614.530 1683.920 ;
        RECT 1608.230 1683.720 1608.550 1683.780 ;
        RECT 1614.210 1683.720 1614.530 1683.780 ;
        RECT 1613.750 14.860 1614.070 14.920 ;
        RECT 1691.490 14.860 1691.810 14.920 ;
        RECT 1613.750 14.720 1691.810 14.860 ;
        RECT 1613.750 14.660 1614.070 14.720 ;
        RECT 1691.490 14.660 1691.810 14.720 ;
      LAYER via ;
        RECT 1608.260 1683.720 1608.520 1683.980 ;
        RECT 1614.240 1683.720 1614.500 1683.980 ;
        RECT 1613.780 14.660 1614.040 14.920 ;
        RECT 1691.520 14.660 1691.780 14.920 ;
      LAYER met2 ;
        RECT 1608.250 1700.000 1608.530 1704.000 ;
        RECT 1608.320 1684.010 1608.460 1700.000 ;
        RECT 1608.260 1683.690 1608.520 1684.010 ;
        RECT 1614.240 1683.690 1614.500 1684.010 ;
        RECT 1614.300 38.490 1614.440 1683.690 ;
        RECT 1613.840 38.350 1614.440 38.490 ;
        RECT 1613.840 14.950 1613.980 38.350 ;
        RECT 1613.780 14.630 1614.040 14.950 ;
        RECT 1691.520 14.630 1691.780 14.950 ;
        RECT 1691.580 2.400 1691.720 14.630 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1346.950 1656.380 1347.270 1656.440 ;
        RECT 1346.580 1656.240 1347.270 1656.380 ;
        RECT 1346.580 1656.100 1346.720 1656.240 ;
        RECT 1346.950 1656.180 1347.270 1656.240 ;
        RECT 1346.490 1655.840 1346.810 1656.100 ;
        RECT 1345.570 1598.920 1345.890 1598.980 ;
        RECT 1346.490 1598.920 1346.810 1598.980 ;
        RECT 1345.570 1598.780 1346.810 1598.920 ;
        RECT 1345.570 1598.720 1345.890 1598.780 ;
        RECT 1346.490 1598.720 1346.810 1598.780 ;
        RECT 1345.570 1545.880 1345.890 1545.940 ;
        RECT 1346.490 1545.880 1346.810 1545.940 ;
        RECT 1345.570 1545.740 1346.810 1545.880 ;
        RECT 1345.570 1545.680 1345.890 1545.740 ;
        RECT 1346.490 1545.680 1346.810 1545.740 ;
        RECT 1345.570 1419.400 1345.890 1419.460 ;
        RECT 1346.490 1419.400 1346.810 1419.460 ;
        RECT 1345.570 1419.260 1346.810 1419.400 ;
        RECT 1345.570 1419.200 1345.890 1419.260 ;
        RECT 1346.490 1419.200 1346.810 1419.260 ;
        RECT 1345.570 1352.760 1345.890 1352.820 ;
        RECT 1346.490 1352.760 1346.810 1352.820 ;
        RECT 1345.570 1352.620 1346.810 1352.760 ;
        RECT 1345.570 1352.560 1345.890 1352.620 ;
        RECT 1346.490 1352.560 1346.810 1352.620 ;
        RECT 731.010 1183.440 731.330 1183.500 ;
        RECT 1346.490 1183.440 1346.810 1183.500 ;
        RECT 731.010 1183.300 1346.810 1183.440 ;
        RECT 731.010 1183.240 731.330 1183.300 ;
        RECT 1346.490 1183.240 1346.810 1183.300 ;
        RECT 728.250 2.960 728.570 3.020 ;
        RECT 731.010 2.960 731.330 3.020 ;
        RECT 728.250 2.820 731.330 2.960 ;
        RECT 728.250 2.760 728.570 2.820 ;
        RECT 731.010 2.760 731.330 2.820 ;
      LAYER via ;
        RECT 1346.980 1656.180 1347.240 1656.440 ;
        RECT 1346.520 1655.840 1346.780 1656.100 ;
        RECT 1345.600 1598.720 1345.860 1598.980 ;
        RECT 1346.520 1598.720 1346.780 1598.980 ;
        RECT 1345.600 1545.680 1345.860 1545.940 ;
        RECT 1346.520 1545.680 1346.780 1545.940 ;
        RECT 1345.600 1419.200 1345.860 1419.460 ;
        RECT 1346.520 1419.200 1346.780 1419.460 ;
        RECT 1345.600 1352.560 1345.860 1352.820 ;
        RECT 1346.520 1352.560 1346.780 1352.820 ;
        RECT 731.040 1183.240 731.300 1183.500 ;
        RECT 1346.520 1183.240 1346.780 1183.500 ;
        RECT 728.280 2.760 728.540 3.020 ;
        RECT 731.040 2.760 731.300 3.020 ;
      LAYER met2 ;
        RECT 1346.970 1700.000 1347.250 1704.000 ;
        RECT 1347.040 1656.470 1347.180 1700.000 ;
        RECT 1346.980 1656.150 1347.240 1656.470 ;
        RECT 1346.520 1655.810 1346.780 1656.130 ;
        RECT 1346.580 1599.010 1346.720 1655.810 ;
        RECT 1345.600 1598.690 1345.860 1599.010 ;
        RECT 1346.520 1598.690 1346.780 1599.010 ;
        RECT 1345.660 1545.970 1345.800 1598.690 ;
        RECT 1345.600 1545.650 1345.860 1545.970 ;
        RECT 1346.520 1545.650 1346.780 1545.970 ;
        RECT 1346.580 1419.490 1346.720 1545.650 ;
        RECT 1345.600 1419.170 1345.860 1419.490 ;
        RECT 1346.520 1419.170 1346.780 1419.490 ;
        RECT 1345.660 1352.850 1345.800 1419.170 ;
        RECT 1345.600 1352.530 1345.860 1352.850 ;
        RECT 1346.520 1352.530 1346.780 1352.850 ;
        RECT 1346.580 1183.530 1346.720 1352.530 ;
        RECT 731.040 1183.210 731.300 1183.530 ;
        RECT 1346.520 1183.210 1346.780 1183.530 ;
        RECT 731.100 3.050 731.240 1183.210 ;
        RECT 728.280 2.730 728.540 3.050 ;
        RECT 731.040 2.730 731.300 3.050 ;
        RECT 728.340 2.400 728.480 2.730 ;
        RECT 728.130 -4.800 728.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 0.300 ;
=======
      LAYER met1 ;
        RECT 1611.450 1688.680 1611.770 1688.740 ;
        RECT 1614.210 1688.680 1614.530 1688.740 ;
        RECT 1611.450 1688.540 1614.530 1688.680 ;
        RECT 1611.450 1688.480 1611.770 1688.540 ;
        RECT 1614.210 1688.480 1614.530 1688.540 ;
        RECT 1614.210 18.600 1614.530 18.660 ;
        RECT 1709.430 18.600 1709.750 18.660 ;
        RECT 1614.210 18.460 1709.750 18.600 ;
        RECT 1614.210 18.400 1614.530 18.460 ;
        RECT 1709.430 18.400 1709.750 18.460 ;
      LAYER via ;
        RECT 1611.480 1688.480 1611.740 1688.740 ;
        RECT 1614.240 1688.480 1614.500 1688.740 ;
        RECT 1614.240 18.400 1614.500 18.660 ;
        RECT 1709.460 18.400 1709.720 18.660 ;
      LAYER met2 ;
        RECT 1611.470 1700.000 1611.750 1704.000 ;
        RECT 1611.540 1688.770 1611.680 1700.000 ;
        RECT 1611.480 1688.450 1611.740 1688.770 ;
        RECT 1614.240 1688.450 1614.500 1688.770 ;
        RECT 1614.300 18.690 1614.440 1688.450 ;
        RECT 1614.240 18.370 1614.500 18.690 ;
        RECT 1709.460 18.370 1709.720 18.690 ;
        RECT 1709.520 2.400 1709.660 18.370 ;
=======
      LAYER li1 ;
        RECT 1705.365 1642.285 1705.535 1686.995 ;
      LAYER mcon ;
        RECT 1705.365 1686.825 1705.535 1686.995 ;
      LAYER met1 ;
        RECT 1613.290 1686.980 1613.610 1687.040 ;
        RECT 1705.305 1686.980 1705.595 1687.025 ;
        RECT 1613.290 1686.840 1705.595 1686.980 ;
        RECT 1613.290 1686.780 1613.610 1686.840 ;
        RECT 1705.305 1686.795 1705.595 1686.840 ;
        RECT 1705.290 1642.440 1705.610 1642.500 ;
        RECT 1705.095 1642.300 1705.610 1642.440 ;
        RECT 1705.290 1642.240 1705.610 1642.300 ;
        RECT 1705.290 2.960 1705.610 3.020 ;
        RECT 1709.430 2.960 1709.750 3.020 ;
        RECT 1705.290 2.820 1709.750 2.960 ;
        RECT 1705.290 2.760 1705.610 2.820 ;
        RECT 1709.430 2.760 1709.750 2.820 ;
      LAYER via ;
        RECT 1613.320 1686.780 1613.580 1687.040 ;
        RECT 1705.320 1642.240 1705.580 1642.500 ;
        RECT 1705.320 2.760 1705.580 3.020 ;
        RECT 1709.460 2.760 1709.720 3.020 ;
      LAYER met2 ;
        RECT 1613.310 1700.000 1613.590 1704.000 ;
        RECT 1613.380 1687.070 1613.520 1700.000 ;
        RECT 1613.320 1686.750 1613.580 1687.070 ;
        RECT 1705.320 1642.210 1705.580 1642.530 ;
        RECT 1705.380 3.050 1705.520 1642.210 ;
        RECT 1705.320 2.730 1705.580 3.050 ;
        RECT 1709.460 2.730 1709.720 3.050 ;
        RECT 1709.520 2.400 1709.660 2.730 ;
>>>>>>> re-updated local openlane
        RECT 1709.310 -4.800 1709.870 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1619.270 1678.140 1619.590 1678.200 ;
        RECT 1621.110 1678.140 1621.430 1678.200 ;
        RECT 1619.270 1678.000 1621.430 1678.140 ;
        RECT 1619.270 1677.940 1619.590 1678.000 ;
        RECT 1621.110 1677.940 1621.430 1678.000 ;
        RECT 1727.370 15.880 1727.690 15.940 ;
        RECT 1651.560 15.740 1727.690 15.880 ;
        RECT 1621.110 15.540 1621.430 15.600 ;
        RECT 1651.560 15.540 1651.700 15.740 ;
        RECT 1727.370 15.680 1727.690 15.740 ;
        RECT 1621.110 15.400 1651.700 15.540 ;
        RECT 1621.110 15.340 1621.430 15.400 ;
      LAYER via ;
        RECT 1619.300 1677.940 1619.560 1678.200 ;
        RECT 1621.140 1677.940 1621.400 1678.200 ;
        RECT 1621.140 15.340 1621.400 15.600 ;
        RECT 1727.400 15.680 1727.660 15.940 ;
      LAYER met2 ;
        RECT 1617.910 1700.410 1618.190 1704.000 ;
        RECT 1617.910 1700.270 1619.500 1700.410 ;
        RECT 1617.910 1700.000 1618.190 1700.270 ;
        RECT 1619.360 1678.230 1619.500 1700.270 ;
        RECT 1619.300 1677.910 1619.560 1678.230 ;
        RECT 1621.140 1677.910 1621.400 1678.230 ;
        RECT 1621.200 15.630 1621.340 1677.910 ;
        RECT 1727.400 15.650 1727.660 15.970 ;
        RECT 1621.140 15.310 1621.400 15.630 ;
        RECT 1727.460 2.400 1727.600 15.650 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 0.300 ;
=======
      LAYER li1 ;
        RECT 1638.665 15.045 1638.835 16.235 ;
        RECT 1653.385 15.215 1653.555 16.575 ;
        RECT 1652.005 15.045 1653.555 15.215 ;
        RECT 1675.465 14.365 1675.635 16.575 ;
        RECT 1732.965 14.365 1734.515 14.535 ;
      LAYER mcon ;
        RECT 1653.385 16.405 1653.555 16.575 ;
        RECT 1638.665 16.065 1638.835 16.235 ;
        RECT 1675.465 16.405 1675.635 16.575 ;
        RECT 1734.345 14.365 1734.515 14.535 ;
      LAYER met1 ;
        RECT 1621.570 1684.940 1621.890 1685.000 ;
        RECT 1631.690 1684.940 1632.010 1685.000 ;
        RECT 1621.570 1684.800 1632.010 1684.940 ;
        RECT 1621.570 1684.740 1621.890 1684.800 ;
        RECT 1631.690 1684.740 1632.010 1684.800 ;
        RECT 1631.690 19.960 1632.010 20.020 ;
        RECT 1633.070 19.960 1633.390 20.020 ;
        RECT 1631.690 19.820 1633.390 19.960 ;
        RECT 1631.690 19.760 1632.010 19.820 ;
        RECT 1633.070 19.760 1633.390 19.820 ;
        RECT 1653.325 16.560 1653.615 16.605 ;
        RECT 1675.405 16.560 1675.695 16.605 ;
        RECT 1653.325 16.420 1675.695 16.560 ;
        RECT 1653.325 16.375 1653.615 16.420 ;
        RECT 1675.405 16.375 1675.695 16.420 ;
        RECT 1633.070 16.220 1633.390 16.280 ;
        RECT 1638.605 16.220 1638.895 16.265 ;
        RECT 1633.070 16.080 1638.895 16.220 ;
        RECT 1633.070 16.020 1633.390 16.080 ;
        RECT 1638.605 16.035 1638.895 16.080 ;
        RECT 1638.605 15.200 1638.895 15.245 ;
        RECT 1651.945 15.200 1652.235 15.245 ;
        RECT 1638.605 15.060 1652.235 15.200 ;
        RECT 1638.605 15.015 1638.895 15.060 ;
        RECT 1651.945 15.015 1652.235 15.060 ;
        RECT 1675.405 14.520 1675.695 14.565 ;
        RECT 1732.905 14.520 1733.195 14.565 ;
        RECT 1675.405 14.380 1733.195 14.520 ;
        RECT 1675.405 14.335 1675.695 14.380 ;
        RECT 1732.905 14.335 1733.195 14.380 ;
        RECT 1734.285 14.520 1734.575 14.565 ;
        RECT 1745.310 14.520 1745.630 14.580 ;
        RECT 1734.285 14.380 1745.630 14.520 ;
        RECT 1734.285 14.335 1734.575 14.380 ;
        RECT 1745.310 14.320 1745.630 14.380 ;
      LAYER via ;
        RECT 1621.600 1684.740 1621.860 1685.000 ;
        RECT 1631.720 1684.740 1631.980 1685.000 ;
        RECT 1631.720 19.760 1631.980 20.020 ;
        RECT 1633.100 19.760 1633.360 20.020 ;
        RECT 1633.100 16.020 1633.360 16.280 ;
        RECT 1745.340 14.320 1745.600 14.580 ;
      LAYER met2 ;
        RECT 1621.130 1700.000 1621.410 1704.000 ;
        RECT 1621.200 1686.130 1621.340 1700.000 ;
        RECT 1621.200 1685.990 1621.800 1686.130 ;
        RECT 1621.660 1685.030 1621.800 1685.990 ;
        RECT 1621.600 1684.710 1621.860 1685.030 ;
        RECT 1631.720 1684.710 1631.980 1685.030 ;
        RECT 1631.780 20.050 1631.920 1684.710 ;
        RECT 1631.720 19.730 1631.980 20.050 ;
        RECT 1633.100 19.730 1633.360 20.050 ;
        RECT 1633.160 16.310 1633.300 19.730 ;
        RECT 1633.100 15.990 1633.360 16.310 ;
        RECT 1745.340 14.290 1745.600 14.610 ;
        RECT 1745.400 2.400 1745.540 14.290 ;
=======
      LAYER met1 ;
        RECT 1622.950 1684.260 1623.270 1684.320 ;
        RECT 1628.010 1684.260 1628.330 1684.320 ;
        RECT 1622.950 1684.120 1628.330 1684.260 ;
        RECT 1622.950 1684.060 1623.270 1684.120 ;
        RECT 1628.010 1684.060 1628.330 1684.120 ;
        RECT 1628.010 16.220 1628.330 16.280 ;
        RECT 1745.310 16.220 1745.630 16.280 ;
        RECT 1628.010 16.080 1745.630 16.220 ;
        RECT 1628.010 16.020 1628.330 16.080 ;
        RECT 1745.310 16.020 1745.630 16.080 ;
      LAYER via ;
        RECT 1622.980 1684.060 1623.240 1684.320 ;
        RECT 1628.040 1684.060 1628.300 1684.320 ;
        RECT 1628.040 16.020 1628.300 16.280 ;
        RECT 1745.340 16.020 1745.600 16.280 ;
      LAYER met2 ;
        RECT 1622.970 1700.000 1623.250 1704.000 ;
        RECT 1623.040 1684.350 1623.180 1700.000 ;
        RECT 1622.980 1684.030 1623.240 1684.350 ;
        RECT 1628.040 1684.030 1628.300 1684.350 ;
        RECT 1628.100 16.310 1628.240 1684.030 ;
        RECT 1628.040 15.990 1628.300 16.310 ;
        RECT 1745.340 15.990 1745.600 16.310 ;
        RECT 1745.400 2.400 1745.540 15.990 ;
>>>>>>> re-updated local openlane
        RECT 1745.190 -4.800 1745.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 0.300 ;
=======
      LAYER met1 ;
        RECT 1625.710 1688.680 1626.030 1688.740 ;
        RECT 1628.010 1688.680 1628.330 1688.740 ;
        RECT 1625.710 1688.540 1628.330 1688.680 ;
        RECT 1625.710 1688.480 1626.030 1688.540 ;
        RECT 1628.010 1688.480 1628.330 1688.540 ;
        RECT 1628.010 15.540 1628.330 15.600 ;
        RECT 1628.010 15.400 1652.620 15.540 ;
        RECT 1628.010 15.340 1628.330 15.400 ;
        RECT 1652.480 15.200 1652.620 15.400 ;
        RECT 1762.790 15.200 1763.110 15.260 ;
        RECT 1652.480 15.060 1763.110 15.200 ;
        RECT 1762.790 15.000 1763.110 15.060 ;
      LAYER via ;
        RECT 1625.740 1688.480 1626.000 1688.740 ;
        RECT 1628.040 1688.480 1628.300 1688.740 ;
        RECT 1628.040 15.340 1628.300 15.600 ;
        RECT 1762.820 15.000 1763.080 15.260 ;
      LAYER met2 ;
        RECT 1625.730 1700.000 1626.010 1704.000 ;
        RECT 1625.800 1688.770 1625.940 1700.000 ;
        RECT 1625.740 1688.450 1626.000 1688.770 ;
        RECT 1628.040 1688.450 1628.300 1688.770 ;
        RECT 1628.100 15.630 1628.240 1688.450 ;
        RECT 1628.040 15.310 1628.300 15.630 ;
        RECT 1762.820 14.970 1763.080 15.290 ;
        RECT 1762.880 2.400 1763.020 14.970 ;
=======
      LAYER li1 ;
        RECT 1644.645 18.785 1644.815 20.655 ;
      LAYER mcon ;
        RECT 1644.645 20.485 1644.815 20.655 ;
      LAYER met1 ;
        RECT 1644.585 20.640 1644.875 20.685 ;
        RECT 1762.790 20.640 1763.110 20.700 ;
        RECT 1644.585 20.500 1763.110 20.640 ;
        RECT 1644.585 20.455 1644.875 20.500 ;
        RECT 1762.790 20.440 1763.110 20.500 ;
        RECT 1627.090 18.940 1627.410 19.000 ;
        RECT 1644.585 18.940 1644.875 18.985 ;
        RECT 1627.090 18.800 1644.875 18.940 ;
        RECT 1627.090 18.740 1627.410 18.800 ;
        RECT 1644.585 18.755 1644.875 18.800 ;
      LAYER via ;
        RECT 1762.820 20.440 1763.080 20.700 ;
        RECT 1627.120 18.740 1627.380 19.000 ;
      LAYER met2 ;
        RECT 1627.570 1700.410 1627.850 1704.000 ;
        RECT 1627.180 1700.270 1627.850 1700.410 ;
        RECT 1627.180 19.030 1627.320 1700.270 ;
        RECT 1627.570 1700.000 1627.850 1700.270 ;
        RECT 1762.820 20.410 1763.080 20.730 ;
        RECT 1627.120 18.710 1627.380 19.030 ;
        RECT 1762.880 2.400 1763.020 20.410 ;
>>>>>>> re-updated local openlane
        RECT 1762.670 -4.800 1763.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 0.300 ;
=======
      LAYER li1 ;
        RECT 1644.645 17.425 1644.815 19.975 ;
        RECT 1656.605 16.745 1656.775 17.595 ;
      LAYER mcon ;
        RECT 1644.645 19.805 1644.815 19.975 ;
        RECT 1656.605 17.425 1656.775 17.595 ;
      LAYER met1 ;
        RECT 1630.770 1688.340 1631.090 1688.400 ;
        RECT 1634.910 1688.340 1635.230 1688.400 ;
        RECT 1630.770 1688.200 1635.230 1688.340 ;
        RECT 1630.770 1688.140 1631.090 1688.200 ;
        RECT 1634.910 1688.140 1635.230 1688.200 ;
=======
      LAYER met1 ;
        RECT 1632.610 1683.920 1632.930 1683.980 ;
        RECT 1634.910 1683.920 1635.230 1683.980 ;
        RECT 1632.610 1683.780 1635.230 1683.920 ;
        RECT 1632.610 1683.720 1632.930 1683.780 ;
        RECT 1634.910 1683.720 1635.230 1683.780 ;
>>>>>>> re-updated local openlane
        RECT 1634.910 19.960 1635.230 20.020 ;
        RECT 1780.730 19.960 1781.050 20.020 ;
        RECT 1634.910 19.820 1781.050 19.960 ;
        RECT 1634.910 19.760 1635.230 19.820 ;
        RECT 1780.730 19.760 1781.050 19.820 ;
      LAYER via ;
        RECT 1632.640 1683.720 1632.900 1683.980 ;
        RECT 1634.940 1683.720 1635.200 1683.980 ;
        RECT 1634.940 19.760 1635.200 20.020 ;
        RECT 1780.760 19.760 1781.020 20.020 ;
      LAYER met2 ;
        RECT 1632.630 1700.000 1632.910 1704.000 ;
        RECT 1632.700 1684.010 1632.840 1700.000 ;
        RECT 1632.640 1683.690 1632.900 1684.010 ;
        RECT 1634.940 1683.690 1635.200 1684.010 ;
        RECT 1635.000 20.050 1635.140 1683.690 ;
        RECT 1634.940 19.730 1635.200 20.050 ;
        RECT 1780.760 19.730 1781.020 20.050 ;
        RECT 1780.820 2.400 1780.960 19.730 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1637.210 1684.260 1637.530 1684.320 ;
        RECT 1640.890 1684.260 1641.210 1684.320 ;
        RECT 1637.210 1684.120 1641.210 1684.260 ;
        RECT 1637.210 1684.060 1637.530 1684.120 ;
        RECT 1640.890 1684.060 1641.210 1684.120 ;
        RECT 1640.890 22.340 1641.210 22.400 ;
        RECT 1798.670 22.340 1798.990 22.400 ;
        RECT 1640.890 22.200 1798.990 22.340 ;
        RECT 1640.890 22.140 1641.210 22.200 ;
        RECT 1798.670 22.140 1798.990 22.200 ;
      LAYER via ;
        RECT 1637.240 1684.060 1637.500 1684.320 ;
        RECT 1640.920 1684.060 1641.180 1684.320 ;
        RECT 1640.920 22.140 1641.180 22.400 ;
        RECT 1798.700 22.140 1798.960 22.400 ;
      LAYER met2 ;
        RECT 1637.230 1700.000 1637.510 1704.000 ;
        RECT 1637.300 1684.350 1637.440 1700.000 ;
        RECT 1637.240 1684.030 1637.500 1684.350 ;
        RECT 1640.920 1684.030 1641.180 1684.350 ;
        RECT 1640.980 22.430 1641.120 1684.030 ;
        RECT 1640.920 22.110 1641.180 22.430 ;
        RECT 1798.700 22.110 1798.960 22.430 ;
        RECT 1798.760 2.400 1798.900 22.110 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1642.270 1684.260 1642.590 1684.320 ;
        RECT 1647.330 1684.260 1647.650 1684.320 ;
        RECT 1642.270 1684.120 1647.650 1684.260 ;
        RECT 1642.270 1684.060 1642.590 1684.120 ;
        RECT 1647.330 1684.060 1647.650 1684.120 ;
        RECT 1647.330 22.680 1647.650 22.740 ;
        RECT 1816.610 22.680 1816.930 22.740 ;
        RECT 1647.330 22.540 1816.930 22.680 ;
        RECT 1647.330 22.480 1647.650 22.540 ;
        RECT 1816.610 22.480 1816.930 22.540 ;
      LAYER via ;
        RECT 1642.300 1684.060 1642.560 1684.320 ;
        RECT 1647.360 1684.060 1647.620 1684.320 ;
        RECT 1647.360 22.480 1647.620 22.740 ;
        RECT 1816.640 22.480 1816.900 22.740 ;
      LAYER met2 ;
        RECT 1642.290 1700.000 1642.570 1704.000 ;
        RECT 1642.360 1684.350 1642.500 1700.000 ;
        RECT 1642.300 1684.030 1642.560 1684.350 ;
        RECT 1647.360 1684.030 1647.620 1684.350 ;
        RECT 1647.420 22.770 1647.560 1684.030 ;
        RECT 1647.360 22.450 1647.620 22.770 ;
        RECT 1816.640 22.450 1816.900 22.770 ;
        RECT 1816.700 2.400 1816.840 22.450 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 0.300 ;
=======
      LAYER li1 ;
        RECT 1801.505 22.185 1801.675 23.375 ;
      LAYER mcon ;
        RECT 1801.505 23.205 1801.675 23.375 ;
      LAYER met1 ;
        RECT 1645.030 1688.340 1645.350 1688.400 ;
        RECT 1648.250 1688.340 1648.570 1688.400 ;
        RECT 1645.030 1688.200 1648.570 1688.340 ;
        RECT 1645.030 1688.140 1645.350 1688.200 ;
        RECT 1648.250 1688.140 1648.570 1688.200 ;
        RECT 1648.250 23.360 1648.570 23.420 ;
        RECT 1801.445 23.360 1801.735 23.405 ;
        RECT 1648.250 23.220 1801.735 23.360 ;
        RECT 1648.250 23.160 1648.570 23.220 ;
        RECT 1801.445 23.175 1801.735 23.220 ;
        RECT 1801.445 22.340 1801.735 22.385 ;
        RECT 1834.550 22.340 1834.870 22.400 ;
        RECT 1801.445 22.200 1834.870 22.340 ;
        RECT 1801.445 22.155 1801.735 22.200 ;
        RECT 1834.550 22.140 1834.870 22.200 ;
      LAYER via ;
        RECT 1645.060 1688.140 1645.320 1688.400 ;
        RECT 1648.280 1688.140 1648.540 1688.400 ;
        RECT 1648.280 23.160 1648.540 23.420 ;
        RECT 1834.580 22.140 1834.840 22.400 ;
      LAYER met2 ;
        RECT 1645.050 1700.000 1645.330 1704.000 ;
        RECT 1645.120 1688.430 1645.260 1700.000 ;
        RECT 1645.060 1688.110 1645.320 1688.430 ;
        RECT 1648.280 1688.110 1648.540 1688.430 ;
        RECT 1648.340 23.450 1648.480 1688.110 ;
        RECT 1648.280 23.130 1648.540 23.450 ;
        RECT 1834.580 22.110 1834.840 22.430 ;
        RECT 1834.640 2.400 1834.780 22.110 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1646.870 23.700 1647.190 23.760 ;
        RECT 1834.550 23.700 1834.870 23.760 ;
        RECT 1646.870 23.560 1834.870 23.700 ;
        RECT 1646.870 23.500 1647.190 23.560 ;
        RECT 1834.550 23.500 1834.870 23.560 ;
      LAYER via ;
        RECT 1646.900 23.500 1647.160 23.760 ;
        RECT 1834.580 23.500 1834.840 23.760 ;
      LAYER met2 ;
        RECT 1646.890 1700.000 1647.170 1704.000 ;
        RECT 1646.960 23.790 1647.100 1700.000 ;
        RECT 1646.900 23.470 1647.160 23.790 ;
        RECT 1834.580 23.470 1834.840 23.790 ;
        RECT 1834.640 2.400 1834.780 23.470 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 0.300 ;
=======
      LAYER met1 ;
        RECT 1654.690 27.100 1655.010 27.160 ;
        RECT 1852.030 27.100 1852.350 27.160 ;
        RECT 1654.690 26.960 1852.350 27.100 ;
        RECT 1654.690 26.900 1655.010 26.960 ;
        RECT 1852.030 26.900 1852.350 26.960 ;
      LAYER via ;
        RECT 1654.720 26.900 1654.980 27.160 ;
        RECT 1852.060 26.900 1852.320 27.160 ;
      LAYER met2 ;
        RECT 1651.950 1700.410 1652.230 1704.000 ;
        RECT 1651.950 1700.270 1653.080 1700.410 ;
        RECT 1651.950 1700.000 1652.230 1700.270 ;
        RECT 1652.940 1677.970 1653.080 1700.270 ;
        RECT 1652.940 1677.830 1654.920 1677.970 ;
        RECT 1654.780 27.190 1654.920 1677.830 ;
        RECT 1654.720 26.870 1654.980 27.190 ;
        RECT 1852.060 26.870 1852.320 27.190 ;
        RECT 1852.120 2.400 1852.260 26.870 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1656.530 1684.260 1656.850 1684.320 ;
        RECT 1661.590 1684.260 1661.910 1684.320 ;
        RECT 1656.530 1684.120 1661.910 1684.260 ;
        RECT 1656.530 1684.060 1656.850 1684.120 ;
        RECT 1661.590 1684.060 1661.910 1684.120 ;
        RECT 1661.590 26.420 1661.910 26.480 ;
        RECT 1869.970 26.420 1870.290 26.480 ;
        RECT 1661.590 26.280 1870.290 26.420 ;
        RECT 1661.590 26.220 1661.910 26.280 ;
        RECT 1869.970 26.220 1870.290 26.280 ;
      LAYER via ;
        RECT 1656.560 1684.060 1656.820 1684.320 ;
        RECT 1661.620 1684.060 1661.880 1684.320 ;
        RECT 1661.620 26.220 1661.880 26.480 ;
        RECT 1870.000 26.220 1870.260 26.480 ;
      LAYER met2 ;
        RECT 1656.550 1700.000 1656.830 1704.000 ;
        RECT 1656.620 1684.350 1656.760 1700.000 ;
        RECT 1656.560 1684.030 1656.820 1684.350 ;
        RECT 1661.620 1684.030 1661.880 1684.350 ;
        RECT 1661.680 26.510 1661.820 1684.030 ;
        RECT 1661.620 26.190 1661.880 26.510 ;
        RECT 1870.000 26.190 1870.260 26.510 ;
        RECT 1870.060 2.400 1870.200 26.190 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 0.300 ;
=======
      LAYER met1 ;
        RECT 1348.330 1608.100 1348.650 1608.160 ;
        RECT 1349.250 1608.100 1349.570 1608.160 ;
        RECT 1348.330 1607.960 1349.570 1608.100 ;
        RECT 1348.330 1607.900 1348.650 1607.960 ;
        RECT 1349.250 1607.900 1349.570 1607.960 ;
        RECT 751.710 1562.880 752.030 1562.940 ;
        RECT 1348.330 1562.880 1348.650 1562.940 ;
        RECT 751.710 1562.740 1348.650 1562.880 ;
        RECT 751.710 1562.680 752.030 1562.740 ;
        RECT 1348.330 1562.680 1348.650 1562.740 ;
        RECT 746.190 2.960 746.510 3.020 ;
        RECT 751.710 2.960 752.030 3.020 ;
        RECT 746.190 2.820 752.030 2.960 ;
        RECT 746.190 2.760 746.510 2.820 ;
        RECT 751.710 2.760 752.030 2.820 ;
      LAYER via ;
        RECT 1348.360 1607.900 1348.620 1608.160 ;
        RECT 1349.280 1607.900 1349.540 1608.160 ;
        RECT 751.740 1562.680 752.000 1562.940 ;
        RECT 1348.360 1562.680 1348.620 1562.940 ;
        RECT 746.220 2.760 746.480 3.020 ;
        RECT 751.740 2.760 752.000 3.020 ;
      LAYER met2 ;
        RECT 1352.030 1700.410 1352.310 1704.000 ;
        RECT 1351.180 1700.270 1352.310 1700.410 ;
        RECT 1351.180 1663.690 1351.320 1700.270 ;
        RECT 1352.030 1700.000 1352.310 1700.270 ;
        RECT 1349.340 1663.550 1351.320 1663.690 ;
        RECT 1349.340 1608.190 1349.480 1663.550 ;
        RECT 1348.360 1607.870 1348.620 1608.190 ;
        RECT 1349.280 1607.870 1349.540 1608.190 ;
        RECT 1348.420 1562.970 1348.560 1607.870 ;
        RECT 751.740 1562.650 752.000 1562.970 ;
        RECT 1348.360 1562.650 1348.620 1562.970 ;
        RECT 751.800 3.050 751.940 1562.650 ;
        RECT 746.220 2.730 746.480 3.050 ;
        RECT 751.740 2.730 752.000 3.050 ;
        RECT 746.280 2.400 746.420 2.730 ;
        RECT 746.070 -4.800 746.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1661.130 25.740 1661.450 25.800 ;
        RECT 1887.910 25.740 1888.230 25.800 ;
        RECT 1661.130 25.600 1888.230 25.740 ;
        RECT 1661.130 25.540 1661.450 25.600 ;
        RECT 1887.910 25.540 1888.230 25.600 ;
      LAYER via ;
        RECT 1661.160 25.540 1661.420 25.800 ;
        RECT 1887.940 25.540 1888.200 25.800 ;
      LAYER met2 ;
        RECT 1661.610 1700.410 1661.890 1704.000 ;
        RECT 1661.220 1700.270 1661.890 1700.410 ;
        RECT 1661.220 25.830 1661.360 1700.270 ;
        RECT 1661.610 1700.000 1661.890 1700.270 ;
        RECT 1661.160 25.510 1661.420 25.830 ;
        RECT 1887.940 25.510 1888.200 25.830 ;
        RECT 1888.000 2.400 1888.140 25.510 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1667.570 25.060 1667.890 25.120 ;
        RECT 1905.850 25.060 1906.170 25.120 ;
        RECT 1667.570 24.920 1906.170 25.060 ;
        RECT 1667.570 24.860 1667.890 24.920 ;
        RECT 1905.850 24.860 1906.170 24.920 ;
      LAYER via ;
        RECT 1667.600 24.860 1667.860 25.120 ;
        RECT 1905.880 24.860 1906.140 25.120 ;
      LAYER met2 ;
        RECT 1666.210 1700.410 1666.490 1704.000 ;
        RECT 1666.210 1700.270 1667.800 1700.410 ;
        RECT 1666.210 1700.000 1666.490 1700.270 ;
        RECT 1667.660 25.150 1667.800 1700.270 ;
        RECT 1667.600 24.830 1667.860 25.150 ;
        RECT 1905.880 24.830 1906.140 25.150 ;
        RECT 1905.940 2.400 1906.080 24.830 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1671.250 1684.260 1671.570 1684.320 ;
        RECT 1675.390 1684.260 1675.710 1684.320 ;
        RECT 1671.250 1684.120 1675.710 1684.260 ;
        RECT 1671.250 1684.060 1671.570 1684.120 ;
        RECT 1675.390 1684.060 1675.710 1684.120 ;
        RECT 1675.390 24.720 1675.710 24.780 ;
        RECT 1923.330 24.720 1923.650 24.780 ;
        RECT 1675.390 24.580 1923.650 24.720 ;
        RECT 1675.390 24.520 1675.710 24.580 ;
        RECT 1923.330 24.520 1923.650 24.580 ;
      LAYER via ;
        RECT 1671.280 1684.060 1671.540 1684.320 ;
        RECT 1675.420 1684.060 1675.680 1684.320 ;
        RECT 1675.420 24.520 1675.680 24.780 ;
        RECT 1923.360 24.520 1923.620 24.780 ;
      LAYER met2 ;
        RECT 1671.270 1700.000 1671.550 1704.000 ;
        RECT 1671.340 1684.350 1671.480 1700.000 ;
        RECT 1671.280 1684.030 1671.540 1684.350 ;
        RECT 1675.420 1684.030 1675.680 1684.350 ;
        RECT 1675.480 24.810 1675.620 1684.030 ;
        RECT 1675.420 24.490 1675.680 24.810 ;
        RECT 1923.360 24.490 1923.620 24.810 ;
        RECT 1923.420 2.400 1923.560 24.490 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 0.300 ;
=======
      LAYER met1 ;
        RECT 1674.930 34.920 1675.250 34.980 ;
        RECT 1941.270 34.920 1941.590 34.980 ;
        RECT 1674.930 34.780 1941.590 34.920 ;
        RECT 1674.930 34.720 1675.250 34.780 ;
        RECT 1941.270 34.720 1941.590 34.780 ;
      LAYER via ;
        RECT 1674.960 34.720 1675.220 34.980 ;
        RECT 1941.300 34.720 1941.560 34.980 ;
      LAYER met2 ;
        RECT 1675.870 1700.410 1676.150 1704.000 ;
        RECT 1675.020 1700.270 1676.150 1700.410 ;
        RECT 1675.020 35.010 1675.160 1700.270 ;
        RECT 1675.870 1700.000 1676.150 1700.270 ;
        RECT 1674.960 34.690 1675.220 35.010 ;
        RECT 1941.300 34.690 1941.560 35.010 ;
        RECT 1941.360 2.400 1941.500 34.690 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1680.910 1684.260 1681.230 1684.320 ;
        RECT 1682.290 1684.260 1682.610 1684.320 ;
        RECT 1680.910 1684.120 1682.610 1684.260 ;
        RECT 1680.910 1684.060 1681.230 1684.120 ;
        RECT 1682.290 1684.060 1682.610 1684.120 ;
        RECT 1682.290 35.260 1682.610 35.320 ;
        RECT 1959.210 35.260 1959.530 35.320 ;
        RECT 1682.290 35.120 1959.530 35.260 ;
        RECT 1682.290 35.060 1682.610 35.120 ;
        RECT 1959.210 35.060 1959.530 35.120 ;
      LAYER via ;
        RECT 1680.940 1684.060 1681.200 1684.320 ;
        RECT 1682.320 1684.060 1682.580 1684.320 ;
        RECT 1682.320 35.060 1682.580 35.320 ;
        RECT 1959.240 35.060 1959.500 35.320 ;
      LAYER met2 ;
        RECT 1680.930 1700.000 1681.210 1704.000 ;
        RECT 1681.000 1684.350 1681.140 1700.000 ;
        RECT 1680.940 1684.030 1681.200 1684.350 ;
        RECT 1682.320 1684.030 1682.580 1684.350 ;
        RECT 1682.380 35.350 1682.520 1684.030 ;
        RECT 1682.320 35.030 1682.580 35.350 ;
        RECT 1959.240 35.030 1959.500 35.350 ;
        RECT 1959.300 2.400 1959.440 35.030 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1685.970 1683.920 1686.290 1683.980 ;
        RECT 1689.190 1683.920 1689.510 1683.980 ;
        RECT 1685.970 1683.780 1689.510 1683.920 ;
        RECT 1685.970 1683.720 1686.290 1683.780 ;
        RECT 1689.190 1683.720 1689.510 1683.780 ;
        RECT 1689.190 35.600 1689.510 35.660 ;
        RECT 1977.150 35.600 1977.470 35.660 ;
        RECT 1689.190 35.460 1977.470 35.600 ;
        RECT 1689.190 35.400 1689.510 35.460 ;
        RECT 1977.150 35.400 1977.470 35.460 ;
      LAYER via ;
        RECT 1686.000 1683.720 1686.260 1683.980 ;
        RECT 1689.220 1683.720 1689.480 1683.980 ;
        RECT 1689.220 35.400 1689.480 35.660 ;
        RECT 1977.180 35.400 1977.440 35.660 ;
      LAYER met2 ;
        RECT 1685.990 1700.000 1686.270 1704.000 ;
        RECT 1686.060 1684.010 1686.200 1700.000 ;
        RECT 1686.000 1683.690 1686.260 1684.010 ;
        RECT 1689.220 1683.690 1689.480 1684.010 ;
        RECT 1689.280 35.690 1689.420 1683.690 ;
        RECT 1689.220 35.370 1689.480 35.690 ;
        RECT 1977.180 35.370 1977.440 35.690 ;
        RECT 1977.240 2.400 1977.380 35.370 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1690.570 1683.920 1690.890 1683.980 ;
        RECT 1696.550 1683.920 1696.870 1683.980 ;
        RECT 1690.570 1683.780 1696.870 1683.920 ;
        RECT 1690.570 1683.720 1690.890 1683.780 ;
        RECT 1696.550 1683.720 1696.870 1683.780 ;
        RECT 1696.550 35.940 1696.870 36.000 ;
        RECT 1995.090 35.940 1995.410 36.000 ;
        RECT 1696.550 35.800 1995.410 35.940 ;
        RECT 1696.550 35.740 1696.870 35.800 ;
        RECT 1995.090 35.740 1995.410 35.800 ;
      LAYER via ;
        RECT 1690.600 1683.720 1690.860 1683.980 ;
        RECT 1696.580 1683.720 1696.840 1683.980 ;
        RECT 1696.580 35.740 1696.840 36.000 ;
        RECT 1995.120 35.740 1995.380 36.000 ;
      LAYER met2 ;
        RECT 1690.590 1700.000 1690.870 1704.000 ;
        RECT 1690.660 1684.010 1690.800 1700.000 ;
        RECT 1690.600 1683.690 1690.860 1684.010 ;
        RECT 1696.580 1683.690 1696.840 1684.010 ;
        RECT 1696.640 36.030 1696.780 1683.690 ;
        RECT 1696.580 35.710 1696.840 36.030 ;
        RECT 1995.120 35.710 1995.380 36.030 ;
        RECT 1995.180 2.400 1995.320 35.710 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1696.090 43.760 1696.410 43.820 ;
        RECT 2012.570 43.760 2012.890 43.820 ;
        RECT 1696.090 43.620 2012.890 43.760 ;
        RECT 1696.090 43.560 1696.410 43.620 ;
        RECT 2012.570 43.560 2012.890 43.620 ;
      LAYER via ;
        RECT 1696.120 43.560 1696.380 43.820 ;
        RECT 2012.600 43.560 2012.860 43.820 ;
      LAYER met2 ;
        RECT 1695.650 1700.410 1695.930 1704.000 ;
        RECT 1695.650 1700.270 1696.320 1700.410 ;
        RECT 1695.650 1700.000 1695.930 1700.270 ;
        RECT 1696.180 43.850 1696.320 1700.270 ;
        RECT 1696.120 43.530 1696.380 43.850 ;
        RECT 2012.600 43.530 2012.860 43.850 ;
        RECT 2012.660 2.400 2012.800 43.530 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 0.300 ;
=======
      LAYER met1 ;
        RECT 1700.230 1684.260 1700.550 1684.320 ;
        RECT 1703.450 1684.260 1703.770 1684.320 ;
        RECT 1700.230 1684.120 1703.770 1684.260 ;
        RECT 1700.230 1684.060 1700.550 1684.120 ;
        RECT 1703.450 1684.060 1703.770 1684.120 ;
        RECT 1703.450 44.100 1703.770 44.160 ;
        RECT 2030.510 44.100 2030.830 44.160 ;
        RECT 1703.450 43.960 2030.830 44.100 ;
        RECT 1703.450 43.900 1703.770 43.960 ;
        RECT 2030.510 43.900 2030.830 43.960 ;
      LAYER via ;
        RECT 1700.260 1684.060 1700.520 1684.320 ;
        RECT 1703.480 1684.060 1703.740 1684.320 ;
        RECT 1703.480 43.900 1703.740 44.160 ;
        RECT 2030.540 43.900 2030.800 44.160 ;
      LAYER met2 ;
        RECT 1700.250 1700.000 1700.530 1704.000 ;
        RECT 1700.320 1684.350 1700.460 1700.000 ;
        RECT 1700.260 1684.030 1700.520 1684.350 ;
        RECT 1703.480 1684.030 1703.740 1684.350 ;
        RECT 1703.540 44.190 1703.680 1684.030 ;
        RECT 1703.480 43.870 1703.740 44.190 ;
        RECT 2030.540 43.870 2030.800 44.190 ;
        RECT 2030.600 2.400 2030.740 43.870 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 0.300 ;
=======
      LAYER met1 ;
        RECT 1705.290 1683.920 1705.610 1683.980 ;
        RECT 1710.350 1683.920 1710.670 1683.980 ;
        RECT 1705.290 1683.780 1710.670 1683.920 ;
        RECT 1705.290 1683.720 1705.610 1683.780 ;
        RECT 1710.350 1683.720 1710.670 1683.780 ;
        RECT 1710.350 44.440 1710.670 44.500 ;
        RECT 2048.450 44.440 2048.770 44.500 ;
        RECT 1710.350 44.300 2048.770 44.440 ;
        RECT 1710.350 44.240 1710.670 44.300 ;
        RECT 2048.450 44.240 2048.770 44.300 ;
      LAYER via ;
        RECT 1705.320 1683.720 1705.580 1683.980 ;
        RECT 1710.380 1683.720 1710.640 1683.980 ;
        RECT 1710.380 44.240 1710.640 44.500 ;
        RECT 2048.480 44.240 2048.740 44.500 ;
      LAYER met2 ;
        RECT 1705.310 1700.000 1705.590 1704.000 ;
        RECT 1705.380 1684.010 1705.520 1700.000 ;
        RECT 1705.320 1683.690 1705.580 1684.010 ;
        RECT 1710.380 1683.690 1710.640 1684.010 ;
        RECT 1710.440 44.530 1710.580 1683.690 ;
        RECT 1710.380 44.210 1710.640 44.530 ;
        RECT 2048.480 44.210 2048.740 44.530 ;
        RECT 2048.540 2.400 2048.680 44.210 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1348.790 1683.920 1349.110 1683.980 ;
        RECT 1356.610 1683.920 1356.930 1683.980 ;
        RECT 1348.790 1683.780 1356.930 1683.920 ;
        RECT 1348.790 1683.720 1349.110 1683.780 ;
        RECT 1356.610 1683.720 1356.930 1683.780 ;
        RECT 765.510 99.860 765.830 99.920 ;
        RECT 1348.790 99.860 1349.110 99.920 ;
        RECT 765.510 99.720 1349.110 99.860 ;
        RECT 765.510 99.660 765.830 99.720 ;
        RECT 1348.790 99.660 1349.110 99.720 ;
      LAYER via ;
        RECT 1348.820 1683.720 1349.080 1683.980 ;
        RECT 1356.640 1683.720 1356.900 1683.980 ;
        RECT 765.540 99.660 765.800 99.920 ;
        RECT 1348.820 99.660 1349.080 99.920 ;
      LAYER met2 ;
        RECT 1356.630 1700.000 1356.910 1704.000 ;
        RECT 1356.700 1684.010 1356.840 1700.000 ;
        RECT 1348.820 1683.690 1349.080 1684.010 ;
        RECT 1356.640 1683.690 1356.900 1684.010 ;
        RECT 1348.880 99.950 1349.020 1683.690 ;
        RECT 765.540 99.630 765.800 99.950 ;
        RECT 1348.820 99.630 1349.080 99.950 ;
        RECT 765.600 3.130 765.740 99.630 ;
        RECT 763.760 2.990 765.740 3.130 ;
        RECT 763.760 2.400 763.900 2.990 ;
        RECT 763.550 -4.800 764.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 0.300 ;
=======
      LAYER met1 ;
        RECT 1710.810 48.180 1711.130 48.240 ;
        RECT 2066.390 48.180 2066.710 48.240 ;
        RECT 1710.810 48.040 2066.710 48.180 ;
        RECT 1710.810 47.980 1711.130 48.040 ;
        RECT 2066.390 47.980 2066.710 48.040 ;
      LAYER via ;
        RECT 1710.840 47.980 1711.100 48.240 ;
        RECT 2066.420 47.980 2066.680 48.240 ;
      LAYER met2 ;
        RECT 1709.910 1700.410 1710.190 1704.000 ;
        RECT 1709.910 1700.270 1711.040 1700.410 ;
        RECT 1709.910 1700.000 1710.190 1700.270 ;
        RECT 1710.900 48.270 1711.040 1700.270 ;
        RECT 1710.840 47.950 1711.100 48.270 ;
        RECT 2066.420 47.950 2066.680 48.270 ;
        RECT 2066.480 2.400 2066.620 47.950 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1717.250 47.840 1717.570 47.900 ;
        RECT 2084.330 47.840 2084.650 47.900 ;
        RECT 1717.250 47.700 2084.650 47.840 ;
        RECT 1717.250 47.640 1717.570 47.700 ;
        RECT 2084.330 47.640 2084.650 47.700 ;
      LAYER via ;
        RECT 1717.280 47.640 1717.540 47.900 ;
        RECT 2084.360 47.640 2084.620 47.900 ;
      LAYER met2 ;
        RECT 1714.970 1700.410 1715.250 1704.000 ;
        RECT 1714.970 1700.270 1716.100 1700.410 ;
        RECT 1714.970 1700.000 1715.250 1700.270 ;
        RECT 1715.960 1684.770 1716.100 1700.270 ;
        RECT 1715.960 1684.630 1717.480 1684.770 ;
        RECT 1717.340 47.930 1717.480 1684.630 ;
        RECT 1717.280 47.610 1717.540 47.930 ;
        RECT 2084.360 47.610 2084.620 47.930 ;
        RECT 2084.420 2.400 2084.560 47.610 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1719.550 1684.260 1719.870 1684.320 ;
        RECT 1723.230 1684.260 1723.550 1684.320 ;
        RECT 1719.550 1684.120 1723.550 1684.260 ;
        RECT 1719.550 1684.060 1719.870 1684.120 ;
        RECT 1723.230 1684.060 1723.550 1684.120 ;
        RECT 1723.230 47.500 1723.550 47.560 ;
        RECT 2101.810 47.500 2102.130 47.560 ;
        RECT 1723.230 47.360 2102.130 47.500 ;
        RECT 1723.230 47.300 1723.550 47.360 ;
        RECT 2101.810 47.300 2102.130 47.360 ;
      LAYER via ;
        RECT 1719.580 1684.060 1719.840 1684.320 ;
        RECT 1723.260 1684.060 1723.520 1684.320 ;
        RECT 1723.260 47.300 1723.520 47.560 ;
        RECT 2101.840 47.300 2102.100 47.560 ;
      LAYER met2 ;
        RECT 1719.570 1700.000 1719.850 1704.000 ;
        RECT 1719.640 1684.350 1719.780 1700.000 ;
        RECT 1719.580 1684.030 1719.840 1684.350 ;
        RECT 1723.260 1684.030 1723.520 1684.350 ;
        RECT 1723.320 47.590 1723.460 1684.030 ;
        RECT 1723.260 47.270 1723.520 47.590 ;
        RECT 2101.840 47.270 2102.100 47.590 ;
        RECT 2101.900 2.400 2102.040 47.270 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1723.690 47.160 1724.010 47.220 ;
        RECT 2119.750 47.160 2120.070 47.220 ;
        RECT 1723.690 47.020 2120.070 47.160 ;
        RECT 1723.690 46.960 1724.010 47.020 ;
        RECT 2119.750 46.960 2120.070 47.020 ;
      LAYER via ;
        RECT 1723.720 46.960 1723.980 47.220 ;
        RECT 2119.780 46.960 2120.040 47.220 ;
      LAYER met2 ;
        RECT 1724.630 1700.410 1724.910 1704.000 ;
        RECT 1723.780 1700.270 1724.910 1700.410 ;
        RECT 1723.780 47.250 1723.920 1700.270 ;
        RECT 1724.630 1700.000 1724.910 1700.270 ;
        RECT 1723.720 46.930 1723.980 47.250 ;
        RECT 2119.780 46.930 2120.040 47.250 ;
        RECT 2119.840 2.400 2119.980 46.930 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 0.300 ;
=======
      LAYER met1 ;
        RECT 1730.590 46.820 1730.910 46.880 ;
        RECT 2137.690 46.820 2138.010 46.880 ;
        RECT 1730.590 46.680 2138.010 46.820 ;
        RECT 1730.590 46.620 1730.910 46.680 ;
        RECT 2137.690 46.620 2138.010 46.680 ;
      LAYER via ;
        RECT 1730.620 46.620 1730.880 46.880 ;
        RECT 2137.720 46.620 2137.980 46.880 ;
      LAYER met2 ;
        RECT 1729.230 1700.410 1729.510 1704.000 ;
        RECT 1729.230 1700.270 1730.820 1700.410 ;
        RECT 1729.230 1700.000 1729.510 1700.270 ;
        RECT 1730.680 46.910 1730.820 1700.270 ;
        RECT 1730.620 46.590 1730.880 46.910 ;
        RECT 2137.720 46.590 2137.980 46.910 ;
        RECT 2137.780 2.400 2137.920 46.590 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 0.300 ;
=======
      LAYER met1 ;
        RECT 1734.270 1683.920 1734.590 1683.980 ;
        RECT 1737.490 1683.920 1737.810 1683.980 ;
        RECT 1734.270 1683.780 1737.810 1683.920 ;
        RECT 1734.270 1683.720 1734.590 1683.780 ;
        RECT 1737.490 1683.720 1737.810 1683.780 ;
        RECT 1737.490 46.480 1737.810 46.540 ;
        RECT 2155.630 46.480 2155.950 46.540 ;
        RECT 1737.490 46.340 2155.950 46.480 ;
        RECT 1737.490 46.280 1737.810 46.340 ;
        RECT 2155.630 46.280 2155.950 46.340 ;
      LAYER via ;
        RECT 1734.300 1683.720 1734.560 1683.980 ;
        RECT 1737.520 1683.720 1737.780 1683.980 ;
        RECT 1737.520 46.280 1737.780 46.540 ;
        RECT 2155.660 46.280 2155.920 46.540 ;
      LAYER met2 ;
        RECT 1734.290 1700.000 1734.570 1704.000 ;
        RECT 1734.360 1684.010 1734.500 1700.000 ;
        RECT 1734.300 1683.690 1734.560 1684.010 ;
        RECT 1737.520 1683.690 1737.780 1684.010 ;
        RECT 1737.580 46.570 1737.720 1683.690 ;
        RECT 1737.520 46.250 1737.780 46.570 ;
        RECT 2155.660 46.250 2155.920 46.570 ;
        RECT 2155.720 2.400 2155.860 46.250 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1738.870 1684.260 1739.190 1684.320 ;
        RECT 1744.390 1684.260 1744.710 1684.320 ;
        RECT 1738.870 1684.120 1744.710 1684.260 ;
        RECT 1738.870 1684.060 1739.190 1684.120 ;
        RECT 1744.390 1684.060 1744.710 1684.120 ;
        RECT 1744.390 46.140 1744.710 46.200 ;
        RECT 2173.110 46.140 2173.430 46.200 ;
        RECT 1744.390 46.000 2173.430 46.140 ;
        RECT 1744.390 45.940 1744.710 46.000 ;
        RECT 2173.110 45.940 2173.430 46.000 ;
      LAYER via ;
        RECT 1738.900 1684.060 1739.160 1684.320 ;
        RECT 1744.420 1684.060 1744.680 1684.320 ;
        RECT 1744.420 45.940 1744.680 46.200 ;
        RECT 2173.140 45.940 2173.400 46.200 ;
      LAYER met2 ;
        RECT 1738.890 1700.000 1739.170 1704.000 ;
        RECT 1738.960 1684.350 1739.100 1700.000 ;
        RECT 1738.900 1684.030 1739.160 1684.350 ;
        RECT 1744.420 1684.030 1744.680 1684.350 ;
        RECT 1744.480 46.230 1744.620 1684.030 ;
        RECT 1744.420 45.910 1744.680 46.230 ;
        RECT 2173.140 45.910 2173.400 46.230 ;
        RECT 2173.200 2.400 2173.340 45.910 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1743.930 45.800 1744.250 45.860 ;
        RECT 2191.050 45.800 2191.370 45.860 ;
        RECT 1743.930 45.660 2191.370 45.800 ;
        RECT 1743.930 45.600 1744.250 45.660 ;
        RECT 2191.050 45.600 2191.370 45.660 ;
      LAYER via ;
        RECT 1743.960 45.600 1744.220 45.860 ;
        RECT 2191.080 45.600 2191.340 45.860 ;
      LAYER met2 ;
        RECT 1743.950 1700.000 1744.230 1704.000 ;
        RECT 1744.020 45.890 1744.160 1700.000 ;
        RECT 1743.960 45.570 1744.220 45.890 ;
        RECT 2191.080 45.570 2191.340 45.890 ;
        RECT 2191.140 2.400 2191.280 45.570 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1748.530 1685.280 1748.850 1685.340 ;
        RECT 1750.830 1685.280 1751.150 1685.340 ;
        RECT 1748.530 1685.140 1751.150 1685.280 ;
        RECT 1748.530 1685.080 1748.850 1685.140 ;
        RECT 1750.830 1685.080 1751.150 1685.140 ;
        RECT 1750.830 45.460 1751.150 45.520 ;
        RECT 2208.990 45.460 2209.310 45.520 ;
        RECT 1750.830 45.320 2209.310 45.460 ;
        RECT 1750.830 45.260 1751.150 45.320 ;
        RECT 2208.990 45.260 2209.310 45.320 ;
      LAYER via ;
        RECT 1748.560 1685.080 1748.820 1685.340 ;
        RECT 1750.860 1685.080 1751.120 1685.340 ;
        RECT 1750.860 45.260 1751.120 45.520 ;
        RECT 2209.020 45.260 2209.280 45.520 ;
      LAYER met2 ;
        RECT 1748.550 1700.000 1748.830 1704.000 ;
        RECT 1748.620 1685.370 1748.760 1700.000 ;
        RECT 1748.560 1685.050 1748.820 1685.370 ;
        RECT 1750.860 1685.050 1751.120 1685.370 ;
        RECT 1750.920 45.550 1751.060 1685.050 ;
        RECT 1750.860 45.230 1751.120 45.550 ;
        RECT 2209.020 45.230 2209.280 45.550 ;
        RECT 2209.080 2.400 2209.220 45.230 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 0.300 ;
=======
      LAYER met1 ;
        RECT 1753.590 1684.600 1753.910 1684.660 ;
        RECT 1758.190 1684.600 1758.510 1684.660 ;
        RECT 1753.590 1684.460 1758.510 1684.600 ;
        RECT 1753.590 1684.400 1753.910 1684.460 ;
        RECT 1758.190 1684.400 1758.510 1684.460 ;
        RECT 1758.190 45.120 1758.510 45.180 ;
        RECT 2226.930 45.120 2227.250 45.180 ;
        RECT 1758.190 44.980 2227.250 45.120 ;
        RECT 1758.190 44.920 1758.510 44.980 ;
        RECT 2226.930 44.920 2227.250 44.980 ;
      LAYER via ;
        RECT 1753.620 1684.400 1753.880 1684.660 ;
        RECT 1758.220 1684.400 1758.480 1684.660 ;
        RECT 1758.220 44.920 1758.480 45.180 ;
        RECT 2226.960 44.920 2227.220 45.180 ;
      LAYER met2 ;
        RECT 1753.610 1700.000 1753.890 1704.000 ;
        RECT 1753.680 1684.690 1753.820 1700.000 ;
        RECT 1753.620 1684.370 1753.880 1684.690 ;
        RECT 1758.220 1684.370 1758.480 1684.690 ;
        RECT 1758.280 45.210 1758.420 1684.370 ;
        RECT 1758.220 44.890 1758.480 45.210 ;
        RECT 2226.960 44.890 2227.220 45.210 ;
        RECT 2227.020 2.400 2227.160 44.890 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1359.370 1695.480 1359.690 1695.540 ;
        RECT 1361.670 1695.480 1361.990 1695.540 ;
        RECT 1359.370 1695.340 1361.990 1695.480 ;
        RECT 1359.370 1695.280 1359.690 1695.340 ;
        RECT 1361.670 1695.280 1361.990 1695.340 ;
        RECT 781.610 41.040 781.930 41.100 ;
        RECT 1359.370 41.040 1359.690 41.100 ;
        RECT 781.610 40.900 1359.690 41.040 ;
        RECT 781.610 40.840 781.930 40.900 ;
        RECT 1359.370 40.840 1359.690 40.900 ;
      LAYER via ;
        RECT 1359.400 1695.280 1359.660 1695.540 ;
        RECT 1361.700 1695.280 1361.960 1695.540 ;
        RECT 781.640 40.840 781.900 41.100 ;
        RECT 1359.400 40.840 1359.660 41.100 ;
      LAYER met2 ;
        RECT 1361.690 1700.000 1361.970 1704.000 ;
        RECT 1361.760 1695.570 1361.900 1700.000 ;
        RECT 1359.400 1695.250 1359.660 1695.570 ;
        RECT 1361.700 1695.250 1361.960 1695.570 ;
        RECT 1359.460 41.130 1359.600 1695.250 ;
        RECT 781.640 40.810 781.900 41.130 ;
        RECT 1359.400 40.810 1359.660 41.130 ;
        RECT 781.700 2.400 781.840 40.810 ;
        RECT 781.490 -4.800 782.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1758.650 44.780 1758.970 44.840 ;
        RECT 2244.870 44.780 2245.190 44.840 ;
        RECT 1758.650 44.640 2245.190 44.780 ;
        RECT 1758.650 44.580 1758.970 44.640 ;
        RECT 2244.870 44.580 2245.190 44.640 ;
      LAYER via ;
        RECT 1758.680 44.580 1758.940 44.840 ;
        RECT 2244.900 44.580 2245.160 44.840 ;
      LAYER met2 ;
        RECT 1758.210 1700.410 1758.490 1704.000 ;
        RECT 1758.210 1700.270 1758.880 1700.410 ;
        RECT 1758.210 1700.000 1758.490 1700.270 ;
        RECT 1758.740 44.870 1758.880 1700.270 ;
        RECT 1758.680 44.550 1758.940 44.870 ;
        RECT 2244.900 44.550 2245.160 44.870 ;
        RECT 2244.960 2.400 2245.100 44.550 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 0.300 ;
=======
      LAYER met1 ;
        RECT 1763.250 1684.260 1763.570 1684.320 ;
        RECT 1765.090 1684.260 1765.410 1684.320 ;
        RECT 1763.250 1684.120 1765.410 1684.260 ;
        RECT 1763.250 1684.060 1763.570 1684.120 ;
        RECT 1765.090 1684.060 1765.410 1684.120 ;
        RECT 1765.090 1562.880 1765.410 1562.940 ;
        RECT 2256.370 1562.880 2256.690 1562.940 ;
        RECT 1765.090 1562.740 2256.690 1562.880 ;
        RECT 1765.090 1562.680 1765.410 1562.740 ;
        RECT 2256.370 1562.680 2256.690 1562.740 ;
        RECT 2256.370 5.680 2256.690 5.740 ;
        RECT 2262.350 5.680 2262.670 5.740 ;
        RECT 2256.370 5.540 2262.670 5.680 ;
        RECT 2256.370 5.480 2256.690 5.540 ;
        RECT 2262.350 5.480 2262.670 5.540 ;
      LAYER via ;
        RECT 1763.280 1684.060 1763.540 1684.320 ;
        RECT 1765.120 1684.060 1765.380 1684.320 ;
        RECT 1765.120 1562.680 1765.380 1562.940 ;
        RECT 2256.400 1562.680 2256.660 1562.940 ;
        RECT 2256.400 5.480 2256.660 5.740 ;
        RECT 2262.380 5.480 2262.640 5.740 ;
      LAYER met2 ;
        RECT 1763.270 1700.000 1763.550 1704.000 ;
        RECT 1763.340 1684.350 1763.480 1700.000 ;
        RECT 1763.280 1684.030 1763.540 1684.350 ;
        RECT 1765.120 1684.030 1765.380 1684.350 ;
        RECT 1765.180 1562.970 1765.320 1684.030 ;
        RECT 1765.120 1562.650 1765.380 1562.970 ;
        RECT 2256.400 1562.650 2256.660 1562.970 ;
        RECT 2256.460 5.770 2256.600 1562.650 ;
        RECT 2256.400 5.450 2256.660 5.770 ;
        RECT 2262.380 5.450 2262.640 5.770 ;
        RECT 2262.440 2.400 2262.580 5.450 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1765.090 45.120 1765.410 45.180 ;
        RECT 2280.290 45.120 2280.610 45.180 ;
        RECT 1765.090 44.980 2280.610 45.120 ;
        RECT 1765.090 44.920 1765.410 44.980 ;
        RECT 2280.290 44.920 2280.610 44.980 ;
      LAYER via ;
        RECT 1765.120 44.920 1765.380 45.180 ;
        RECT 2280.320 44.920 2280.580 45.180 ;
      LAYER met2 ;
        RECT 1765.570 1700.410 1765.850 1704.000 ;
        RECT 1765.180 1700.270 1765.850 1700.410 ;
        RECT 1765.180 45.210 1765.320 1700.270 ;
        RECT 1765.570 1700.000 1765.850 1700.270 ;
        RECT 1765.120 44.890 1765.380 45.210 ;
        RECT 2280.320 44.890 2280.580 45.210 ;
        RECT 2280.380 2.400 2280.520 44.890 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 2277.145 1587.205 2277.315 1594.175 ;
        RECT 2277.145 766.105 2277.315 814.215 ;
        RECT 2277.145 669.545 2277.315 717.655 ;
        RECT 2277.145 572.645 2277.315 620.755 ;
        RECT 2277.145 476.085 2277.315 524.195 ;
        RECT 2277.145 379.525 2277.315 427.635 ;
        RECT 2277.145 331.245 2277.315 339.235 ;
        RECT 2277.145 186.405 2277.315 234.175 ;
      LAYER mcon ;
        RECT 2277.145 1594.005 2277.315 1594.175 ;
        RECT 2277.145 814.045 2277.315 814.215 ;
        RECT 2277.145 717.485 2277.315 717.655 ;
        RECT 2277.145 620.585 2277.315 620.755 ;
        RECT 2277.145 524.025 2277.315 524.195 ;
        RECT 2277.145 427.465 2277.315 427.635 ;
        RECT 2277.145 339.065 2277.315 339.235 ;
        RECT 2277.145 234.005 2277.315 234.175 ;
      LAYER met1 ;
        RECT 1767.850 1680.520 1768.170 1680.580 ;
        RECT 2277.070 1680.520 2277.390 1680.580 ;
        RECT 1767.850 1680.380 2277.390 1680.520 ;
        RECT 1767.850 1680.320 1768.170 1680.380 ;
        RECT 2277.070 1680.320 2277.390 1680.380 ;
        RECT 2277.070 1594.160 2277.390 1594.220 ;
        RECT 2276.875 1594.020 2277.390 1594.160 ;
        RECT 2277.070 1593.960 2277.390 1594.020 ;
        RECT 2277.070 1587.360 2277.390 1587.420 ;
        RECT 2276.875 1587.220 2277.390 1587.360 ;
        RECT 2277.070 1587.160 2277.390 1587.220 ;
        RECT 2277.070 1208.060 2277.390 1208.320 ;
        RECT 2277.160 1207.640 2277.300 1208.060 ;
        RECT 2277.070 1207.380 2277.390 1207.640 ;
        RECT 2276.150 1152.500 2276.470 1152.560 ;
        RECT 2276.610 1152.500 2276.930 1152.560 ;
        RECT 2276.150 1152.360 2276.930 1152.500 ;
        RECT 2276.150 1152.300 2276.470 1152.360 ;
        RECT 2276.610 1152.300 2276.930 1152.360 ;
        RECT 2276.150 911.100 2276.470 911.160 ;
        RECT 2277.070 911.100 2277.390 911.160 ;
        RECT 2276.150 910.960 2277.390 911.100 ;
        RECT 2276.150 910.900 2276.470 910.960 ;
        RECT 2277.070 910.900 2277.390 910.960 ;
        RECT 2276.150 869.280 2276.470 869.340 ;
        RECT 2277.070 869.280 2277.390 869.340 ;
        RECT 2276.150 869.140 2277.390 869.280 ;
        RECT 2276.150 869.080 2276.470 869.140 ;
        RECT 2277.070 869.080 2277.390 869.140 ;
        RECT 2277.070 814.200 2277.390 814.260 ;
        RECT 2276.875 814.060 2277.390 814.200 ;
        RECT 2277.070 814.000 2277.390 814.060 ;
        RECT 2277.070 766.260 2277.390 766.320 ;
        RECT 2276.875 766.120 2277.390 766.260 ;
        RECT 2277.070 766.060 2277.390 766.120 ;
        RECT 2277.070 717.640 2277.390 717.700 ;
        RECT 2276.875 717.500 2277.390 717.640 ;
        RECT 2277.070 717.440 2277.390 717.500 ;
        RECT 2277.070 669.700 2277.390 669.760 ;
        RECT 2276.875 669.560 2277.390 669.700 ;
        RECT 2277.070 669.500 2277.390 669.560 ;
        RECT 2277.070 620.740 2277.390 620.800 ;
        RECT 2276.875 620.600 2277.390 620.740 ;
        RECT 2277.070 620.540 2277.390 620.600 ;
        RECT 2277.070 572.800 2277.390 572.860 ;
        RECT 2276.875 572.660 2277.390 572.800 ;
        RECT 2277.070 572.600 2277.390 572.660 ;
        RECT 2277.070 524.180 2277.390 524.240 ;
        RECT 2276.875 524.040 2277.390 524.180 ;
        RECT 2277.070 523.980 2277.390 524.040 ;
        RECT 2277.070 476.240 2277.390 476.300 ;
        RECT 2276.875 476.100 2277.390 476.240 ;
        RECT 2277.070 476.040 2277.390 476.100 ;
        RECT 2277.070 427.620 2277.390 427.680 ;
        RECT 2276.875 427.480 2277.390 427.620 ;
        RECT 2277.070 427.420 2277.390 427.480 ;
        RECT 2277.070 379.680 2277.390 379.740 ;
        RECT 2276.875 379.540 2277.390 379.680 ;
        RECT 2277.070 379.480 2277.390 379.540 ;
        RECT 2277.070 339.220 2277.390 339.280 ;
        RECT 2276.875 339.080 2277.390 339.220 ;
        RECT 2277.070 339.020 2277.390 339.080 ;
        RECT 2277.070 331.400 2277.390 331.460 ;
        RECT 2276.875 331.260 2277.390 331.400 ;
        RECT 2277.070 331.200 2277.390 331.260 ;
        RECT 2275.690 283.120 2276.010 283.180 ;
        RECT 2277.070 283.120 2277.390 283.180 ;
        RECT 2275.690 282.980 2277.390 283.120 ;
        RECT 2275.690 282.920 2276.010 282.980 ;
        RECT 2277.070 282.920 2277.390 282.980 ;
        RECT 2277.070 234.160 2277.390 234.220 ;
        RECT 2276.875 234.020 2277.390 234.160 ;
        RECT 2277.070 233.960 2277.390 234.020 ;
        RECT 2277.070 186.560 2277.390 186.620 ;
        RECT 2276.875 186.420 2277.390 186.560 ;
        RECT 2277.070 186.360 2277.390 186.420 ;
        RECT 2276.610 138.620 2276.930 138.680 ;
        RECT 2277.070 138.620 2277.390 138.680 ;
        RECT 2276.610 138.480 2277.390 138.620 ;
        RECT 2276.610 138.420 2276.930 138.480 ;
        RECT 2277.070 138.420 2277.390 138.480 ;
        RECT 2276.610 137.940 2276.930 138.000 ;
        RECT 2280.290 137.940 2280.610 138.000 ;
        RECT 2276.610 137.800 2280.610 137.940 ;
        RECT 2276.610 137.740 2276.930 137.800 ;
        RECT 2280.290 137.740 2280.610 137.800 ;
      LAYER via ;
        RECT 1767.880 1680.320 1768.140 1680.580 ;
        RECT 2277.100 1680.320 2277.360 1680.580 ;
        RECT 2277.100 1593.960 2277.360 1594.220 ;
        RECT 2277.100 1587.160 2277.360 1587.420 ;
        RECT 2277.100 1208.060 2277.360 1208.320 ;
        RECT 2277.100 1207.380 2277.360 1207.640 ;
        RECT 2276.180 1152.300 2276.440 1152.560 ;
        RECT 2276.640 1152.300 2276.900 1152.560 ;
        RECT 2276.180 910.900 2276.440 911.160 ;
        RECT 2277.100 910.900 2277.360 911.160 ;
        RECT 2276.180 869.080 2276.440 869.340 ;
        RECT 2277.100 869.080 2277.360 869.340 ;
        RECT 2277.100 814.000 2277.360 814.260 ;
        RECT 2277.100 766.060 2277.360 766.320 ;
        RECT 2277.100 717.440 2277.360 717.700 ;
        RECT 2277.100 669.500 2277.360 669.760 ;
        RECT 2277.100 620.540 2277.360 620.800 ;
        RECT 2277.100 572.600 2277.360 572.860 ;
        RECT 2277.100 523.980 2277.360 524.240 ;
        RECT 2277.100 476.040 2277.360 476.300 ;
        RECT 2277.100 427.420 2277.360 427.680 ;
        RECT 2277.100 379.480 2277.360 379.740 ;
        RECT 2277.100 339.020 2277.360 339.280 ;
        RECT 2277.100 331.200 2277.360 331.460 ;
        RECT 2275.720 282.920 2275.980 283.180 ;
        RECT 2277.100 282.920 2277.360 283.180 ;
        RECT 2277.100 233.960 2277.360 234.220 ;
        RECT 2277.100 186.360 2277.360 186.620 ;
        RECT 2276.640 138.420 2276.900 138.680 ;
        RECT 2277.100 138.420 2277.360 138.680 ;
        RECT 2276.640 137.740 2276.900 138.000 ;
        RECT 2280.320 137.740 2280.580 138.000 ;
      LAYER met2 ;
        RECT 1767.870 1700.000 1768.150 1704.000 ;
        RECT 1767.940 1680.610 1768.080 1700.000 ;
        RECT 1767.880 1680.290 1768.140 1680.610 ;
        RECT 2277.100 1680.290 2277.360 1680.610 ;
        RECT 2277.160 1594.250 2277.300 1680.290 ;
        RECT 2277.100 1593.930 2277.360 1594.250 ;
        RECT 2277.100 1587.130 2277.360 1587.450 ;
        RECT 2277.160 1208.350 2277.300 1587.130 ;
        RECT 2277.100 1208.030 2277.360 1208.350 ;
        RECT 2277.100 1207.350 2277.360 1207.670 ;
        RECT 2277.160 1200.610 2277.300 1207.350 ;
        RECT 2276.700 1200.470 2277.300 1200.610 ;
        RECT 2276.700 1152.590 2276.840 1200.470 ;
        RECT 2276.180 1152.270 2276.440 1152.590 ;
        RECT 2276.640 1152.270 2276.900 1152.590 ;
        RECT 2276.240 1055.885 2276.380 1152.270 ;
        RECT 2276.170 1055.515 2276.450 1055.885 ;
        RECT 2277.090 1055.515 2277.370 1055.885 ;
        RECT 2277.160 911.190 2277.300 1055.515 ;
        RECT 2276.180 910.870 2276.440 911.190 ;
        RECT 2277.100 910.870 2277.360 911.190 ;
        RECT 2276.240 869.370 2276.380 910.870 ;
        RECT 2276.180 869.050 2276.440 869.370 ;
        RECT 2277.100 869.050 2277.360 869.370 ;
        RECT 2277.160 862.650 2277.300 869.050 ;
        RECT 2277.160 862.510 2277.760 862.650 ;
        RECT 2277.620 821.170 2277.760 862.510 ;
        RECT 2277.160 821.030 2277.760 821.170 ;
        RECT 2277.160 814.290 2277.300 821.030 ;
        RECT 2277.100 813.970 2277.360 814.290 ;
        RECT 2277.100 766.030 2277.360 766.350 ;
        RECT 2277.160 717.730 2277.300 766.030 ;
        RECT 2277.100 717.410 2277.360 717.730 ;
        RECT 2277.100 669.470 2277.360 669.790 ;
        RECT 2277.160 620.830 2277.300 669.470 ;
        RECT 2277.100 620.510 2277.360 620.830 ;
        RECT 2277.100 572.570 2277.360 572.890 ;
        RECT 2277.160 524.270 2277.300 572.570 ;
        RECT 2277.100 523.950 2277.360 524.270 ;
        RECT 2277.100 476.010 2277.360 476.330 ;
        RECT 2277.160 427.710 2277.300 476.010 ;
        RECT 2277.100 427.390 2277.360 427.710 ;
        RECT 2277.100 379.450 2277.360 379.770 ;
        RECT 2277.160 339.310 2277.300 379.450 ;
        RECT 2277.100 338.990 2277.360 339.310 ;
        RECT 2277.100 331.170 2277.360 331.490 ;
        RECT 2277.160 331.005 2277.300 331.170 ;
        RECT 2275.710 330.635 2275.990 331.005 ;
        RECT 2277.090 330.635 2277.370 331.005 ;
        RECT 2275.780 283.210 2275.920 330.635 ;
        RECT 2275.720 282.890 2275.980 283.210 ;
        RECT 2277.100 282.890 2277.360 283.210 ;
        RECT 2277.160 234.250 2277.300 282.890 ;
        RECT 2277.100 233.930 2277.360 234.250 ;
        RECT 2277.100 186.330 2277.360 186.650 ;
        RECT 2277.160 138.710 2277.300 186.330 ;
        RECT 2276.640 138.390 2276.900 138.710 ;
        RECT 2277.100 138.390 2277.360 138.710 ;
        RECT 2276.700 138.030 2276.840 138.390 ;
        RECT 2276.640 137.710 2276.900 138.030 ;
        RECT 2280.320 137.710 2280.580 138.030 ;
        RECT 2280.380 2.400 2280.520 137.710 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
      LAYER via2 ;
        RECT 2276.170 1055.560 2276.450 1055.840 ;
        RECT 2277.090 1055.560 2277.370 1055.840 ;
        RECT 2275.710 330.680 2275.990 330.960 ;
        RECT 2277.090 330.680 2277.370 330.960 ;
      LAYER met3 ;
        RECT 2276.145 1055.850 2276.475 1055.865 ;
        RECT 2277.065 1055.850 2277.395 1055.865 ;
        RECT 2276.145 1055.550 2277.395 1055.850 ;
        RECT 2276.145 1055.535 2276.475 1055.550 ;
        RECT 2277.065 1055.535 2277.395 1055.550 ;
        RECT 2275.685 330.970 2276.015 330.985 ;
        RECT 2277.065 330.970 2277.395 330.985 ;
        RECT 2275.685 330.670 2277.395 330.970 ;
        RECT 2275.685 330.655 2276.015 330.670 ;
        RECT 2277.065 330.655 2277.395 330.670 ;
>>>>>>> re-updated local openlane
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1772.910 1659.780 1773.230 1659.840 ;
        RECT 2298.230 1659.780 2298.550 1659.840 ;
        RECT 1772.910 1659.640 2298.550 1659.780 ;
        RECT 1772.910 1659.580 1773.230 1659.640 ;
        RECT 2298.230 1659.580 2298.550 1659.640 ;
      LAYER via ;
        RECT 1772.940 1659.580 1773.200 1659.840 ;
        RECT 2298.260 1659.580 2298.520 1659.840 ;
      LAYER met2 ;
        RECT 1772.930 1700.000 1773.210 1704.000 ;
        RECT 1773.000 1659.870 1773.140 1700.000 ;
        RECT 1772.940 1659.550 1773.200 1659.870 ;
        RECT 2298.260 1659.550 2298.520 1659.870 ;
        RECT 2298.320 2.400 2298.460 1659.550 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1778.890 1548.940 1779.210 1549.000 ;
        RECT 2311.570 1548.940 2311.890 1549.000 ;
        RECT 1778.890 1548.800 2311.890 1548.940 ;
        RECT 1778.890 1548.740 1779.210 1548.800 ;
        RECT 2311.570 1548.740 2311.890 1548.800 ;
        RECT 2311.570 62.120 2311.890 62.180 ;
        RECT 2316.170 62.120 2316.490 62.180 ;
        RECT 2311.570 61.980 2316.490 62.120 ;
        RECT 2311.570 61.920 2311.890 61.980 ;
        RECT 2316.170 61.920 2316.490 61.980 ;
      LAYER via ;
        RECT 1778.920 1548.740 1779.180 1549.000 ;
        RECT 2311.600 1548.740 2311.860 1549.000 ;
        RECT 2311.600 61.920 2311.860 62.180 ;
        RECT 2316.200 61.920 2316.460 62.180 ;
      LAYER met2 ;
        RECT 1777.530 1700.410 1777.810 1704.000 ;
        RECT 1777.530 1700.270 1779.120 1700.410 ;
        RECT 1777.530 1700.000 1777.810 1700.270 ;
        RECT 1778.980 1549.030 1779.120 1700.270 ;
        RECT 1778.920 1548.710 1779.180 1549.030 ;
        RECT 2311.600 1548.710 2311.860 1549.030 ;
        RECT 2311.660 62.210 2311.800 1548.710 ;
        RECT 2311.600 61.890 2311.860 62.210 ;
        RECT 2316.200 61.890 2316.460 62.210 ;
        RECT 2316.260 2.400 2316.400 61.890 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1782.570 1683.920 1782.890 1683.980 ;
        RECT 1785.790 1683.920 1786.110 1683.980 ;
        RECT 1782.570 1683.780 1786.110 1683.920 ;
        RECT 1782.570 1683.720 1782.890 1683.780 ;
        RECT 1785.790 1683.720 1786.110 1683.780 ;
        RECT 1785.790 1617.960 1786.110 1618.020 ;
        RECT 2332.270 1617.960 2332.590 1618.020 ;
        RECT 1785.790 1617.820 2332.590 1617.960 ;
        RECT 1785.790 1617.760 1786.110 1617.820 ;
        RECT 2332.270 1617.760 2332.590 1617.820 ;
        RECT 2331.810 48.520 2332.130 48.580 ;
        RECT 2334.110 48.520 2334.430 48.580 ;
        RECT 2331.810 48.380 2334.430 48.520 ;
        RECT 2331.810 48.320 2332.130 48.380 ;
        RECT 2334.110 48.320 2334.430 48.380 ;
      LAYER via ;
        RECT 1782.600 1683.720 1782.860 1683.980 ;
        RECT 1785.820 1683.720 1786.080 1683.980 ;
        RECT 1785.820 1617.760 1786.080 1618.020 ;
        RECT 2332.300 1617.760 2332.560 1618.020 ;
        RECT 2331.840 48.320 2332.100 48.580 ;
        RECT 2334.140 48.320 2334.400 48.580 ;
      LAYER met2 ;
        RECT 1782.590 1700.000 1782.870 1704.000 ;
        RECT 1782.660 1684.010 1782.800 1700.000 ;
        RECT 1782.600 1683.690 1782.860 1684.010 ;
        RECT 1785.820 1683.690 1786.080 1684.010 ;
        RECT 1785.880 1618.050 1786.020 1683.690 ;
        RECT 1785.820 1617.730 1786.080 1618.050 ;
        RECT 2332.300 1617.730 2332.560 1618.050 ;
        RECT 2332.360 72.490 2332.500 1617.730 ;
        RECT 2331.900 72.350 2332.500 72.490 ;
        RECT 2331.900 48.610 2332.040 72.350 ;
        RECT 2331.840 48.290 2332.100 48.610 ;
        RECT 2334.140 48.290 2334.400 48.610 ;
        RECT 2334.200 2.400 2334.340 48.290 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1787.170 1684.600 1787.490 1684.660 ;
        RECT 1792.690 1684.600 1793.010 1684.660 ;
        RECT 1787.170 1684.460 1793.010 1684.600 ;
        RECT 1787.170 1684.400 1787.490 1684.460 ;
        RECT 1792.690 1684.400 1793.010 1684.460 ;
        RECT 1792.690 1542.140 1793.010 1542.200 ;
        RECT 2346.070 1542.140 2346.390 1542.200 ;
        RECT 1792.690 1542.000 2346.390 1542.140 ;
        RECT 1792.690 1541.940 1793.010 1542.000 ;
        RECT 2346.070 1541.940 2346.390 1542.000 ;
        RECT 2346.070 62.120 2346.390 62.180 ;
        RECT 2351.590 62.120 2351.910 62.180 ;
        RECT 2346.070 61.980 2351.910 62.120 ;
        RECT 2346.070 61.920 2346.390 61.980 ;
        RECT 2351.590 61.920 2351.910 61.980 ;
      LAYER via ;
        RECT 1787.200 1684.400 1787.460 1684.660 ;
        RECT 1792.720 1684.400 1792.980 1684.660 ;
        RECT 1792.720 1541.940 1792.980 1542.200 ;
        RECT 2346.100 1541.940 2346.360 1542.200 ;
        RECT 2346.100 61.920 2346.360 62.180 ;
        RECT 2351.620 61.920 2351.880 62.180 ;
      LAYER met2 ;
        RECT 1787.190 1700.000 1787.470 1704.000 ;
        RECT 1787.260 1684.690 1787.400 1700.000 ;
        RECT 1787.200 1684.370 1787.460 1684.690 ;
        RECT 1792.720 1684.370 1792.980 1684.690 ;
        RECT 1792.780 1542.230 1792.920 1684.370 ;
        RECT 1792.720 1541.910 1792.980 1542.230 ;
        RECT 2346.100 1541.910 2346.360 1542.230 ;
        RECT 2346.160 62.210 2346.300 1541.910 ;
        RECT 2346.100 61.890 2346.360 62.210 ;
        RECT 2351.620 61.890 2351.880 62.210 ;
        RECT 2351.680 2.400 2351.820 61.890 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 0.300 ;
=======
      LAYER met1 ;
        RECT 1792.230 1624.760 1792.550 1624.820 ;
        RECT 2366.770 1624.760 2367.090 1624.820 ;
        RECT 1792.230 1624.620 2367.090 1624.760 ;
        RECT 1792.230 1624.560 1792.550 1624.620 ;
        RECT 2366.770 1624.560 2367.090 1624.620 ;
        RECT 2366.770 62.120 2367.090 62.180 ;
        RECT 2369.530 62.120 2369.850 62.180 ;
        RECT 2366.770 61.980 2369.850 62.120 ;
        RECT 2366.770 61.920 2367.090 61.980 ;
        RECT 2369.530 61.920 2369.850 61.980 ;
      LAYER via ;
        RECT 1792.260 1624.560 1792.520 1624.820 ;
        RECT 2366.800 1624.560 2367.060 1624.820 ;
        RECT 2366.800 61.920 2367.060 62.180 ;
        RECT 2369.560 61.920 2369.820 62.180 ;
      LAYER met2 ;
        RECT 1792.250 1700.000 1792.530 1704.000 ;
        RECT 1792.320 1624.850 1792.460 1700.000 ;
        RECT 1792.260 1624.530 1792.520 1624.850 ;
        RECT 2366.800 1624.530 2367.060 1624.850 ;
        RECT 2366.860 62.210 2367.000 1624.530 ;
        RECT 2366.800 61.890 2367.060 62.210 ;
        RECT 2369.560 61.890 2369.820 62.210 ;
        RECT 2369.620 2.400 2369.760 61.890 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1794.530 1687.660 1794.850 1687.720 ;
        RECT 1799.590 1687.660 1799.910 1687.720 ;
        RECT 1794.530 1687.520 1799.910 1687.660 ;
        RECT 1794.530 1687.460 1794.850 1687.520 ;
        RECT 1799.590 1687.460 1799.910 1687.520 ;
        RECT 1799.590 53.960 1799.910 54.020 ;
        RECT 2387.930 53.960 2388.250 54.020 ;
        RECT 1799.590 53.820 2388.250 53.960 ;
        RECT 1799.590 53.760 1799.910 53.820 ;
        RECT 2387.930 53.760 2388.250 53.820 ;
      LAYER via ;
        RECT 1794.560 1687.460 1794.820 1687.720 ;
        RECT 1799.620 1687.460 1799.880 1687.720 ;
        RECT 1799.620 53.760 1799.880 54.020 ;
        RECT 2387.960 53.760 2388.220 54.020 ;
      LAYER met2 ;
        RECT 1794.550 1700.000 1794.830 1704.000 ;
        RECT 1794.620 1687.750 1794.760 1700.000 ;
        RECT 1794.560 1687.430 1794.820 1687.750 ;
        RECT 1799.620 1687.430 1799.880 1687.750 ;
        RECT 1799.680 54.050 1799.820 1687.430 ;
        RECT 1799.620 53.730 1799.880 54.050 ;
        RECT 2387.960 53.730 2388.220 54.050 ;
        RECT 2388.020 17.410 2388.160 53.730 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
=======
      LAYER li1 ;
        RECT 2387.545 2.805 2387.715 14.195 ;
      LAYER mcon ;
        RECT 2387.545 14.025 2387.715 14.195 ;
      LAYER met1 ;
        RECT 1796.830 1684.260 1797.150 1684.320 ;
        RECT 1799.130 1684.260 1799.450 1684.320 ;
        RECT 1796.830 1684.120 1799.450 1684.260 ;
        RECT 1796.830 1684.060 1797.150 1684.120 ;
        RECT 1799.130 1684.060 1799.450 1684.120 ;
        RECT 1799.130 1535.340 1799.450 1535.400 ;
        RECT 2387.930 1535.340 2388.250 1535.400 ;
        RECT 1799.130 1535.200 2388.250 1535.340 ;
        RECT 1799.130 1535.140 1799.450 1535.200 ;
        RECT 2387.930 1535.140 2388.250 1535.200 ;
        RECT 2387.485 14.180 2387.775 14.225 ;
        RECT 2387.930 14.180 2388.250 14.240 ;
        RECT 2387.485 14.040 2388.250 14.180 ;
        RECT 2387.485 13.995 2387.775 14.040 ;
        RECT 2387.930 13.980 2388.250 14.040 ;
        RECT 2387.470 2.960 2387.790 3.020 ;
        RECT 2387.275 2.820 2387.790 2.960 ;
        RECT 2387.470 2.760 2387.790 2.820 ;
      LAYER via ;
        RECT 1796.860 1684.060 1797.120 1684.320 ;
        RECT 1799.160 1684.060 1799.420 1684.320 ;
        RECT 1799.160 1535.140 1799.420 1535.400 ;
        RECT 2387.960 1535.140 2388.220 1535.400 ;
        RECT 2387.960 13.980 2388.220 14.240 ;
        RECT 2387.500 2.760 2387.760 3.020 ;
      LAYER met2 ;
        RECT 1796.850 1700.000 1797.130 1704.000 ;
        RECT 1796.920 1684.350 1797.060 1700.000 ;
        RECT 1796.860 1684.030 1797.120 1684.350 ;
        RECT 1799.160 1684.030 1799.420 1684.350 ;
        RECT 1799.220 1535.430 1799.360 1684.030 ;
        RECT 1799.160 1535.110 1799.420 1535.430 ;
        RECT 2387.960 1535.110 2388.220 1535.430 ;
        RECT 2388.020 14.270 2388.160 1535.110 ;
        RECT 2387.960 13.950 2388.220 14.270 ;
        RECT 2387.500 2.730 2387.760 3.050 ;
        RECT 2387.560 2.400 2387.700 2.730 ;
>>>>>>> re-updated local openlane
        RECT 2387.350 -4.800 2387.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1802.350 1652.980 1802.670 1653.040 ;
        RECT 2401.270 1652.980 2401.590 1653.040 ;
        RECT 1802.350 1652.840 2401.590 1652.980 ;
        RECT 1802.350 1652.780 1802.670 1652.840 ;
        RECT 2401.270 1652.780 2401.590 1652.840 ;
        RECT 2401.270 62.120 2401.590 62.180 ;
        RECT 2405.410 62.120 2405.730 62.180 ;
        RECT 2401.270 61.980 2405.730 62.120 ;
        RECT 2401.270 61.920 2401.590 61.980 ;
        RECT 2405.410 61.920 2405.730 61.980 ;
      LAYER via ;
        RECT 1802.380 1652.780 1802.640 1653.040 ;
        RECT 2401.300 1652.780 2401.560 1653.040 ;
        RECT 2401.300 61.920 2401.560 62.180 ;
        RECT 2405.440 61.920 2405.700 62.180 ;
      LAYER met2 ;
        RECT 1801.910 1700.410 1802.190 1704.000 ;
        RECT 1801.910 1700.270 1802.580 1700.410 ;
        RECT 1801.910 1700.000 1802.190 1700.270 ;
        RECT 1802.440 1653.070 1802.580 1700.270 ;
        RECT 1802.380 1652.750 1802.640 1653.070 ;
        RECT 2401.300 1652.750 2401.560 1653.070 ;
        RECT 2401.360 62.210 2401.500 1652.750 ;
        RECT 2401.300 61.890 2401.560 62.210 ;
        RECT 2405.440 61.890 2405.700 62.210 ;
        RECT 2405.500 2.400 2405.640 61.890 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 0.300 ;
=======
      LAYER met1 ;
        RECT 799.550 41.380 799.870 41.440 ;
        RECT 1366.730 41.380 1367.050 41.440 ;
        RECT 799.550 41.240 1367.050 41.380 ;
        RECT 799.550 41.180 799.870 41.240 ;
        RECT 1366.730 41.180 1367.050 41.240 ;
      LAYER via ;
        RECT 799.580 41.180 799.840 41.440 ;
        RECT 1366.760 41.180 1367.020 41.440 ;
      LAYER met2 ;
        RECT 1366.290 1700.410 1366.570 1704.000 ;
        RECT 1366.290 1700.270 1366.960 1700.410 ;
        RECT 1366.290 1700.000 1366.570 1700.270 ;
        RECT 1366.820 41.470 1366.960 1700.270 ;
        RECT 799.580 41.150 799.840 41.470 ;
        RECT 1366.760 41.150 1367.020 41.470 ;
        RECT 799.640 2.400 799.780 41.150 ;
        RECT 799.430 -4.800 799.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1318.890 1678.140 1319.210 1678.200 ;
        RECT 1323.490 1678.140 1323.810 1678.200 ;
        RECT 1318.890 1678.000 1323.810 1678.140 ;
        RECT 1318.890 1677.940 1319.210 1678.000 ;
        RECT 1323.490 1677.940 1323.810 1678.000 ;
        RECT 644.990 40.700 645.310 40.760 ;
        RECT 1318.890 40.700 1319.210 40.760 ;
        RECT 644.990 40.560 1319.210 40.700 ;
        RECT 644.990 40.500 645.310 40.560 ;
        RECT 1318.890 40.500 1319.210 40.560 ;
      LAYER via ;
        RECT 1318.920 1677.940 1319.180 1678.200 ;
        RECT 1323.520 1677.940 1323.780 1678.200 ;
        RECT 645.020 40.500 645.280 40.760 ;
        RECT 1318.920 40.500 1319.180 40.760 ;
      LAYER met2 ;
        RECT 1324.430 1700.410 1324.710 1704.000 ;
        RECT 1323.580 1700.270 1324.710 1700.410 ;
        RECT 1323.580 1678.230 1323.720 1700.270 ;
        RECT 1324.430 1700.000 1324.710 1700.270 ;
        RECT 1318.920 1677.910 1319.180 1678.230 ;
        RECT 1323.520 1677.910 1323.780 1678.230 ;
        RECT 1318.980 40.790 1319.120 1677.910 ;
        RECT 645.020 40.470 645.280 40.790 ;
        RECT 1318.920 40.470 1319.180 40.790 ;
        RECT 645.080 2.400 645.220 40.470 ;
        RECT 644.870 -4.800 645.430 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 645.010 41.000 645.290 41.280 ;
        RECT 1320.290 41.000 1320.570 41.280 ;
      LAYER met3 ;
        RECT 644.985 41.290 645.315 41.305 ;
        RECT 1320.265 41.290 1320.595 41.305 ;
        RECT 644.985 40.990 1320.595 41.290 ;
        RECT 644.985 40.975 645.315 40.990 ;
        RECT 1320.265 40.975 1320.595 40.990 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1808.330 1684.260 1808.650 1684.320 ;
        RECT 1813.850 1684.260 1814.170 1684.320 ;
        RECT 1808.330 1684.120 1814.170 1684.260 ;
        RECT 1808.330 1684.060 1808.650 1684.120 ;
        RECT 1813.850 1684.060 1814.170 1684.120 ;
        RECT 1813.850 231.100 1814.170 231.160 ;
        RECT 2429.330 231.100 2429.650 231.160 ;
        RECT 1813.850 230.960 2429.650 231.100 ;
        RECT 1813.850 230.900 1814.170 230.960 ;
        RECT 2429.330 230.900 2429.650 230.960 ;
      LAYER via ;
        RECT 1808.360 1684.060 1808.620 1684.320 ;
        RECT 1813.880 1684.060 1814.140 1684.320 ;
        RECT 1813.880 230.900 1814.140 231.160 ;
        RECT 2429.360 230.900 2429.620 231.160 ;
      LAYER met2 ;
        RECT 1808.350 1700.000 1808.630 1704.000 ;
        RECT 1808.420 1684.350 1808.560 1700.000 ;
        RECT 1808.360 1684.030 1808.620 1684.350 ;
        RECT 1813.880 1684.030 1814.140 1684.350 ;
        RECT 1813.940 231.190 1814.080 1684.030 ;
        RECT 1813.880 230.870 1814.140 231.190 ;
        RECT 2429.360 230.870 2429.620 231.190 ;
        RECT 2429.420 35.090 2429.560 230.870 ;
        RECT 2428.960 34.950 2429.560 35.090 ;
        RECT 2428.960 2.400 2429.100 34.950 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 0.300 ;
=======
      LAYER met1 ;
        RECT 1813.390 1528.200 1813.710 1528.260 ;
        RECT 2442.670 1528.200 2442.990 1528.260 ;
        RECT 1813.390 1528.060 2442.990 1528.200 ;
        RECT 1813.390 1528.000 1813.710 1528.060 ;
        RECT 2442.670 1528.000 2442.990 1528.060 ;
        RECT 2442.670 62.120 2442.990 62.180 ;
        RECT 2446.810 62.120 2447.130 62.180 ;
        RECT 2442.670 61.980 2447.130 62.120 ;
        RECT 2442.670 61.920 2442.990 61.980 ;
        RECT 2446.810 61.920 2447.130 61.980 ;
      LAYER via ;
        RECT 1813.420 1528.000 1813.680 1528.260 ;
        RECT 2442.700 1528.000 2442.960 1528.260 ;
        RECT 2442.700 61.920 2442.960 62.180 ;
        RECT 2446.840 61.920 2447.100 62.180 ;
      LAYER met2 ;
        RECT 1812.950 1700.410 1813.230 1704.000 ;
        RECT 1812.950 1700.270 1813.620 1700.410 ;
        RECT 1812.950 1700.000 1813.230 1700.270 ;
        RECT 1813.480 1528.290 1813.620 1700.270 ;
        RECT 1813.420 1527.970 1813.680 1528.290 ;
        RECT 2442.700 1527.970 2442.960 1528.290 ;
        RECT 2442.760 62.210 2442.900 1527.970 ;
        RECT 2442.700 61.890 2442.960 62.210 ;
        RECT 2446.840 61.890 2447.100 62.210 ;
        RECT 2446.900 2.400 2447.040 61.890 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1815.230 1683.920 1815.550 1683.980 ;
        RECT 1819.370 1683.920 1819.690 1683.980 ;
        RECT 1815.230 1683.780 1819.690 1683.920 ;
        RECT 1815.230 1683.720 1815.550 1683.780 ;
        RECT 1819.370 1683.720 1819.690 1683.780 ;
        RECT 1819.830 52.600 1820.150 52.660 ;
        RECT 2463.370 52.600 2463.690 52.660 ;
        RECT 1819.830 52.460 2463.690 52.600 ;
        RECT 1819.830 52.400 1820.150 52.460 ;
        RECT 2463.370 52.400 2463.690 52.460 ;
        RECT 2463.370 2.960 2463.690 3.020 ;
=======
      LAYER li1 ;
        RECT 2463.905 1594.005 2464.075 1604.375 ;
        RECT 2463.445 1497.445 2463.615 1545.555 ;
        RECT 2463.445 1400.885 2463.615 1448.995 ;
        RECT 2463.445 1304.325 2463.615 1352.435 ;
        RECT 2463.445 1207.425 2463.615 1255.875 ;
        RECT 2463.445 628.065 2463.615 675.835 ;
        RECT 2463.445 531.505 2463.615 579.615 ;
        RECT 2463.445 434.945 2463.615 483.055 ;
        RECT 2463.445 338.045 2463.615 386.155 ;
        RECT 2463.445 145.605 2463.615 193.035 ;
        RECT 2463.445 48.365 2463.615 137.955 ;
      LAYER mcon ;
        RECT 2463.905 1604.205 2464.075 1604.375 ;
        RECT 2463.445 1545.385 2463.615 1545.555 ;
        RECT 2463.445 1448.825 2463.615 1448.995 ;
        RECT 2463.445 1352.265 2463.615 1352.435 ;
        RECT 2463.445 1255.705 2463.615 1255.875 ;
        RECT 2463.445 675.665 2463.615 675.835 ;
        RECT 2463.445 579.445 2463.615 579.615 ;
        RECT 2463.445 482.885 2463.615 483.055 ;
        RECT 2463.445 385.985 2463.615 386.155 ;
        RECT 2463.445 192.865 2463.615 193.035 ;
        RECT 2463.445 137.785 2463.615 137.955 ;
      LAYER met1 ;
        RECT 1819.830 1604.360 1820.150 1604.420 ;
        RECT 2463.845 1604.360 2464.135 1604.405 ;
        RECT 1819.830 1604.220 2464.135 1604.360 ;
        RECT 1819.830 1604.160 1820.150 1604.220 ;
        RECT 2463.845 1604.175 2464.135 1604.220 ;
        RECT 2463.370 1594.160 2463.690 1594.220 ;
        RECT 2463.845 1594.160 2464.135 1594.205 ;
        RECT 2463.370 1594.020 2464.135 1594.160 ;
        RECT 2463.370 1593.960 2463.690 1594.020 ;
        RECT 2463.845 1593.975 2464.135 1594.020 ;
        RECT 2463.370 1545.540 2463.690 1545.600 ;
        RECT 2463.370 1545.400 2463.885 1545.540 ;
        RECT 2463.370 1545.340 2463.690 1545.400 ;
        RECT 2463.370 1497.600 2463.690 1497.660 ;
        RECT 2463.370 1497.460 2463.885 1497.600 ;
        RECT 2463.370 1497.400 2463.690 1497.460 ;
        RECT 2463.370 1448.980 2463.690 1449.040 ;
        RECT 2463.370 1448.840 2463.885 1448.980 ;
        RECT 2463.370 1448.780 2463.690 1448.840 ;
        RECT 2463.370 1401.040 2463.690 1401.100 ;
        RECT 2463.370 1400.900 2463.885 1401.040 ;
        RECT 2463.370 1400.840 2463.690 1400.900 ;
        RECT 2463.370 1352.420 2463.690 1352.480 ;
        RECT 2463.370 1352.280 2463.885 1352.420 ;
        RECT 2463.370 1352.220 2463.690 1352.280 ;
        RECT 2463.370 1304.480 2463.690 1304.540 ;
        RECT 2463.370 1304.340 2463.885 1304.480 ;
        RECT 2463.370 1304.280 2463.690 1304.340 ;
        RECT 2463.370 1255.860 2463.690 1255.920 ;
        RECT 2463.370 1255.720 2463.885 1255.860 ;
        RECT 2463.370 1255.660 2463.690 1255.720 ;
        RECT 2463.370 1207.580 2463.690 1207.640 ;
        RECT 2463.370 1207.440 2463.885 1207.580 ;
        RECT 2463.370 1207.380 2463.690 1207.440 ;
        RECT 2463.370 1111.020 2463.690 1111.080 ;
        RECT 2464.290 1111.020 2464.610 1111.080 ;
        RECT 2463.370 1110.880 2464.610 1111.020 ;
        RECT 2463.370 1110.820 2463.690 1110.880 ;
        RECT 2464.290 1110.820 2464.610 1110.880 ;
        RECT 2463.370 1014.460 2463.690 1014.520 ;
        RECT 2464.290 1014.460 2464.610 1014.520 ;
        RECT 2463.370 1014.320 2464.610 1014.460 ;
        RECT 2463.370 1014.260 2463.690 1014.320 ;
        RECT 2464.290 1014.260 2464.610 1014.320 ;
        RECT 2463.370 917.900 2463.690 917.960 ;
        RECT 2464.290 917.900 2464.610 917.960 ;
        RECT 2463.370 917.760 2464.610 917.900 ;
        RECT 2463.370 917.700 2463.690 917.760 ;
        RECT 2464.290 917.700 2464.610 917.760 ;
        RECT 2463.370 772.720 2463.690 772.780 ;
        RECT 2464.290 772.720 2464.610 772.780 ;
        RECT 2463.370 772.580 2464.610 772.720 ;
        RECT 2463.370 772.520 2463.690 772.580 ;
        RECT 2464.290 772.520 2464.610 772.580 ;
        RECT 2463.370 675.820 2463.690 675.880 ;
        RECT 2463.370 675.680 2463.885 675.820 ;
        RECT 2463.370 675.620 2463.690 675.680 ;
        RECT 2463.370 628.220 2463.690 628.280 ;
        RECT 2463.370 628.080 2463.885 628.220 ;
        RECT 2463.370 628.020 2463.690 628.080 ;
        RECT 2463.370 579.600 2463.690 579.660 ;
        RECT 2463.370 579.460 2463.885 579.600 ;
        RECT 2463.370 579.400 2463.690 579.460 ;
        RECT 2463.370 531.660 2463.690 531.720 ;
        RECT 2463.370 531.520 2463.885 531.660 ;
        RECT 2463.370 531.460 2463.690 531.520 ;
        RECT 2463.370 483.040 2463.690 483.100 ;
        RECT 2463.370 482.900 2463.885 483.040 ;
        RECT 2463.370 482.840 2463.690 482.900 ;
        RECT 2463.370 435.100 2463.690 435.160 ;
        RECT 2463.370 434.960 2463.885 435.100 ;
        RECT 2463.370 434.900 2463.690 434.960 ;
        RECT 2463.370 386.140 2463.690 386.200 ;
        RECT 2463.370 386.000 2463.885 386.140 ;
        RECT 2463.370 385.940 2463.690 386.000 ;
        RECT 2463.370 338.200 2463.690 338.260 ;
        RECT 2463.370 338.060 2463.885 338.200 ;
        RECT 2463.370 338.000 2463.690 338.060 ;
        RECT 2463.370 193.020 2463.690 193.080 ;
        RECT 2463.370 192.880 2463.885 193.020 ;
        RECT 2463.370 192.820 2463.690 192.880 ;
        RECT 2463.370 145.760 2463.690 145.820 ;
        RECT 2463.370 145.620 2463.885 145.760 ;
        RECT 2463.370 145.560 2463.690 145.620 ;
        RECT 2463.370 137.940 2463.690 138.000 ;
        RECT 2463.175 137.800 2463.690 137.940 ;
        RECT 2463.370 137.740 2463.690 137.800 ;
        RECT 2463.385 48.520 2463.675 48.565 ;
        RECT 2464.750 48.520 2465.070 48.580 ;
        RECT 2463.385 48.380 2465.070 48.520 ;
        RECT 2463.385 48.335 2463.675 48.380 ;
        RECT 2464.750 48.320 2465.070 48.380 ;
>>>>>>> re-updated local openlane
        RECT 2464.750 2.960 2465.070 3.020 ;
        RECT 2465.210 2.960 2465.530 3.020 ;
        RECT 2464.750 2.820 2465.530 2.960 ;
        RECT 2464.750 2.760 2465.070 2.820 ;
        RECT 2465.210 2.760 2465.530 2.820 ;
      LAYER via ;
        RECT 1819.860 1604.160 1820.120 1604.420 ;
        RECT 2463.400 1593.960 2463.660 1594.220 ;
        RECT 2463.400 1545.340 2463.660 1545.600 ;
        RECT 2463.400 1497.400 2463.660 1497.660 ;
        RECT 2463.400 1448.780 2463.660 1449.040 ;
        RECT 2463.400 1400.840 2463.660 1401.100 ;
        RECT 2463.400 1352.220 2463.660 1352.480 ;
        RECT 2463.400 1304.280 2463.660 1304.540 ;
        RECT 2463.400 1255.660 2463.660 1255.920 ;
        RECT 2463.400 1207.380 2463.660 1207.640 ;
        RECT 2463.400 1110.820 2463.660 1111.080 ;
        RECT 2464.320 1110.820 2464.580 1111.080 ;
        RECT 2463.400 1014.260 2463.660 1014.520 ;
        RECT 2464.320 1014.260 2464.580 1014.520 ;
        RECT 2463.400 917.700 2463.660 917.960 ;
        RECT 2464.320 917.700 2464.580 917.960 ;
        RECT 2463.400 772.520 2463.660 772.780 ;
        RECT 2464.320 772.520 2464.580 772.780 ;
        RECT 2463.400 675.620 2463.660 675.880 ;
        RECT 2463.400 628.020 2463.660 628.280 ;
        RECT 2463.400 579.400 2463.660 579.660 ;
        RECT 2463.400 531.460 2463.660 531.720 ;
        RECT 2463.400 482.840 2463.660 483.100 ;
        RECT 2463.400 434.900 2463.660 435.160 ;
        RECT 2463.400 385.940 2463.660 386.200 ;
        RECT 2463.400 338.000 2463.660 338.260 ;
        RECT 2463.400 192.820 2463.660 193.080 ;
        RECT 2463.400 145.560 2463.660 145.820 ;
        RECT 2463.400 137.740 2463.660 138.000 ;
        RECT 2464.780 48.320 2465.040 48.580 ;
        RECT 2464.780 2.760 2465.040 3.020 ;
        RECT 2465.240 2.760 2465.500 3.020 ;
      LAYER met2 ;
        RECT 1818.010 1700.410 1818.290 1704.000 ;
        RECT 1818.010 1700.270 1819.600 1700.410 ;
        RECT 1818.010 1700.000 1818.290 1700.270 ;
        RECT 1819.460 1677.970 1819.600 1700.270 ;
        RECT 1819.460 1677.830 1820.060 1677.970 ;
        RECT 1819.920 1604.450 1820.060 1677.830 ;
        RECT 1819.860 1604.130 1820.120 1604.450 ;
        RECT 2463.400 1593.930 2463.660 1594.250 ;
        RECT 2463.460 1545.630 2463.600 1593.930 ;
        RECT 2463.400 1545.310 2463.660 1545.630 ;
        RECT 2463.400 1497.370 2463.660 1497.690 ;
        RECT 2463.460 1449.070 2463.600 1497.370 ;
        RECT 2463.400 1448.750 2463.660 1449.070 ;
        RECT 2463.400 1400.810 2463.660 1401.130 ;
        RECT 2463.460 1352.510 2463.600 1400.810 ;
        RECT 2463.400 1352.190 2463.660 1352.510 ;
        RECT 2463.400 1304.250 2463.660 1304.570 ;
        RECT 2463.460 1255.950 2463.600 1304.250 ;
        RECT 2463.400 1255.630 2463.660 1255.950 ;
        RECT 2463.400 1207.350 2463.660 1207.670 ;
        RECT 2463.460 1159.245 2463.600 1207.350 ;
        RECT 2463.390 1158.875 2463.670 1159.245 ;
        RECT 2464.310 1158.875 2464.590 1159.245 ;
        RECT 2464.380 1111.110 2464.520 1158.875 ;
        RECT 2463.400 1110.790 2463.660 1111.110 ;
        RECT 2464.320 1110.790 2464.580 1111.110 ;
        RECT 2463.460 1062.685 2463.600 1110.790 ;
        RECT 2463.390 1062.315 2463.670 1062.685 ;
        RECT 2464.310 1062.315 2464.590 1062.685 ;
        RECT 2464.380 1014.550 2464.520 1062.315 ;
        RECT 2463.400 1014.230 2463.660 1014.550 ;
        RECT 2464.320 1014.230 2464.580 1014.550 ;
        RECT 2463.460 966.125 2463.600 1014.230 ;
        RECT 2463.390 965.755 2463.670 966.125 ;
        RECT 2464.310 965.755 2464.590 966.125 ;
        RECT 2464.380 917.990 2464.520 965.755 ;
        RECT 2463.400 917.670 2463.660 917.990 ;
        RECT 2464.320 917.670 2464.580 917.990 ;
        RECT 2463.460 869.565 2463.600 917.670 ;
        RECT 2463.390 869.195 2463.670 869.565 ;
        RECT 2464.310 869.195 2464.590 869.565 ;
        RECT 2464.380 821.285 2464.520 869.195 ;
        RECT 2463.390 820.915 2463.670 821.285 ;
        RECT 2464.310 820.915 2464.590 821.285 ;
        RECT 2463.460 772.810 2463.600 820.915 ;
        RECT 2463.400 772.490 2463.660 772.810 ;
        RECT 2464.320 772.490 2464.580 772.810 ;
        RECT 2464.380 724.725 2464.520 772.490 ;
        RECT 2463.390 724.355 2463.670 724.725 ;
        RECT 2464.310 724.355 2464.590 724.725 ;
        RECT 2463.460 675.910 2463.600 724.355 ;
        RECT 2463.400 675.590 2463.660 675.910 ;
        RECT 2463.400 627.990 2463.660 628.310 ;
        RECT 2463.460 579.690 2463.600 627.990 ;
        RECT 2463.400 579.370 2463.660 579.690 ;
        RECT 2463.400 531.430 2463.660 531.750 ;
        RECT 2463.460 483.130 2463.600 531.430 ;
        RECT 2463.400 482.810 2463.660 483.130 ;
        RECT 2463.400 434.870 2463.660 435.190 ;
        RECT 2463.460 386.230 2463.600 434.870 ;
        RECT 2463.400 385.910 2463.660 386.230 ;
        RECT 2463.400 337.970 2463.660 338.290 ;
        RECT 2463.460 290.885 2463.600 337.970 ;
        RECT 2463.390 290.515 2463.670 290.885 ;
        RECT 2463.390 289.835 2463.670 290.205 ;
        RECT 2463.460 193.110 2463.600 289.835 ;
        RECT 2463.400 192.790 2463.660 193.110 ;
        RECT 2463.400 145.530 2463.660 145.850 ;
        RECT 2463.460 138.030 2463.600 145.530 ;
        RECT 2463.400 137.710 2463.660 138.030 ;
        RECT 2464.780 48.290 2465.040 48.610 ;
        RECT 2464.840 48.010 2464.980 48.290 ;
        RECT 2464.840 47.870 2465.440 48.010 ;
        RECT 2465.300 3.050 2465.440 47.870 ;
        RECT 2464.780 2.730 2465.040 3.050 ;
        RECT 2465.240 2.730 2465.500 3.050 ;
        RECT 2464.840 2.400 2464.980 2.730 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 2463.390 1158.920 2463.670 1159.200 ;
        RECT 2464.310 1158.920 2464.590 1159.200 ;
        RECT 2463.390 1062.360 2463.670 1062.640 ;
        RECT 2464.310 1062.360 2464.590 1062.640 ;
        RECT 2463.390 965.800 2463.670 966.080 ;
        RECT 2464.310 965.800 2464.590 966.080 ;
        RECT 2463.390 869.240 2463.670 869.520 ;
        RECT 2464.310 869.240 2464.590 869.520 ;
        RECT 2463.390 820.960 2463.670 821.240 ;
        RECT 2464.310 820.960 2464.590 821.240 ;
        RECT 2463.390 724.400 2463.670 724.680 ;
        RECT 2464.310 724.400 2464.590 724.680 ;
        RECT 2463.390 290.560 2463.670 290.840 ;
        RECT 2463.390 289.880 2463.670 290.160 ;
      LAYER met3 ;
        RECT 2463.365 1159.210 2463.695 1159.225 ;
        RECT 2464.285 1159.210 2464.615 1159.225 ;
        RECT 2463.365 1158.910 2464.615 1159.210 ;
        RECT 2463.365 1158.895 2463.695 1158.910 ;
        RECT 2464.285 1158.895 2464.615 1158.910 ;
        RECT 2463.365 1062.650 2463.695 1062.665 ;
        RECT 2464.285 1062.650 2464.615 1062.665 ;
        RECT 2463.365 1062.350 2464.615 1062.650 ;
        RECT 2463.365 1062.335 2463.695 1062.350 ;
        RECT 2464.285 1062.335 2464.615 1062.350 ;
        RECT 2463.365 966.090 2463.695 966.105 ;
        RECT 2464.285 966.090 2464.615 966.105 ;
        RECT 2463.365 965.790 2464.615 966.090 ;
        RECT 2463.365 965.775 2463.695 965.790 ;
        RECT 2464.285 965.775 2464.615 965.790 ;
        RECT 2463.365 869.530 2463.695 869.545 ;
        RECT 2464.285 869.530 2464.615 869.545 ;
        RECT 2463.365 869.230 2464.615 869.530 ;
        RECT 2463.365 869.215 2463.695 869.230 ;
        RECT 2464.285 869.215 2464.615 869.230 ;
        RECT 2463.365 821.250 2463.695 821.265 ;
        RECT 2464.285 821.250 2464.615 821.265 ;
        RECT 2463.365 820.950 2464.615 821.250 ;
        RECT 2463.365 820.935 2463.695 820.950 ;
        RECT 2464.285 820.935 2464.615 820.950 ;
        RECT 2463.365 724.690 2463.695 724.705 ;
        RECT 2464.285 724.690 2464.615 724.705 ;
        RECT 2463.365 724.390 2464.615 724.690 ;
        RECT 2463.365 724.375 2463.695 724.390 ;
        RECT 2464.285 724.375 2464.615 724.390 ;
        RECT 2463.365 290.850 2463.695 290.865 ;
        RECT 2463.150 290.535 2463.695 290.850 ;
        RECT 2463.150 290.185 2463.450 290.535 ;
        RECT 2463.150 289.870 2463.695 290.185 ;
        RECT 2463.365 289.855 2463.695 289.870 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 0.300 ;
=======
      LAYER li1 ;
        RECT 1825.425 19.125 1825.595 19.975 ;
      LAYER mcon ;
        RECT 1825.425 19.805 1825.595 19.975 ;
      LAYER met1 ;
        RECT 1825.365 19.960 1825.655 20.005 ;
        RECT 2482.690 19.960 2483.010 20.020 ;
        RECT 1825.365 19.820 2483.010 19.960 ;
        RECT 1825.365 19.775 1825.655 19.820 ;
        RECT 2482.690 19.760 2483.010 19.820 ;
        RECT 1821.210 19.280 1821.530 19.340 ;
        RECT 1825.365 19.280 1825.655 19.325 ;
        RECT 1821.210 19.140 1825.655 19.280 ;
        RECT 1821.210 19.080 1821.530 19.140 ;
        RECT 1825.365 19.095 1825.655 19.140 ;
      LAYER via ;
        RECT 2482.720 19.760 2482.980 20.020 ;
        RECT 1821.240 19.080 1821.500 19.340 ;
      LAYER met2 ;
        RECT 1820.310 1700.410 1820.590 1704.000 ;
        RECT 1820.310 1700.270 1821.440 1700.410 ;
        RECT 1820.310 1700.000 1820.590 1700.270 ;
        RECT 1821.300 19.370 1821.440 1700.270 ;
        RECT 2482.720 19.730 2482.980 20.050 ;
        RECT 1821.240 19.050 1821.500 19.370 ;
        RECT 2482.780 2.400 2482.920 19.730 ;
=======
      LAYER met1 ;
        RECT 1823.050 1683.920 1823.370 1683.980 ;
        RECT 1827.650 1683.920 1827.970 1683.980 ;
        RECT 1823.050 1683.780 1827.970 1683.920 ;
        RECT 1823.050 1683.720 1823.370 1683.780 ;
        RECT 1827.650 1683.720 1827.970 1683.780 ;
        RECT 1827.650 1521.400 1827.970 1521.460 ;
        RECT 2477.170 1521.400 2477.490 1521.460 ;
        RECT 1827.650 1521.260 2477.490 1521.400 ;
        RECT 1827.650 1521.200 1827.970 1521.260 ;
        RECT 2477.170 1521.200 2477.490 1521.260 ;
      LAYER via ;
        RECT 1823.080 1683.720 1823.340 1683.980 ;
        RECT 1827.680 1683.720 1827.940 1683.980 ;
        RECT 1827.680 1521.200 1827.940 1521.460 ;
        RECT 2477.200 1521.200 2477.460 1521.460 ;
      LAYER met2 ;
        RECT 1823.070 1700.000 1823.350 1704.000 ;
        RECT 1823.140 1684.010 1823.280 1700.000 ;
        RECT 1823.080 1683.690 1823.340 1684.010 ;
        RECT 1827.680 1683.690 1827.940 1684.010 ;
        RECT 1827.740 1521.490 1827.880 1683.690 ;
        RECT 1827.680 1521.170 1827.940 1521.490 ;
        RECT 2477.200 1521.170 2477.460 1521.490 ;
        RECT 2477.260 16.730 2477.400 1521.170 ;
        RECT 2477.260 16.590 2482.920 16.730 ;
        RECT 2482.780 2.400 2482.920 16.590 ;
>>>>>>> re-updated local openlane
        RECT 2482.570 -4.800 2483.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 0.300 ;
=======
      LAYER met1 ;
        RECT 1826.730 1514.600 1827.050 1514.660 ;
        RECT 2497.870 1514.600 2498.190 1514.660 ;
        RECT 1826.730 1514.460 2498.190 1514.600 ;
        RECT 1826.730 1514.400 1827.050 1514.460 ;
        RECT 2497.870 1514.400 2498.190 1514.460 ;
      LAYER via ;
        RECT 1826.760 1514.400 1827.020 1514.660 ;
        RECT 2497.900 1514.400 2498.160 1514.660 ;
      LAYER met2 ;
        RECT 1827.670 1700.410 1827.950 1704.000 ;
        RECT 1826.820 1700.270 1827.950 1700.410 ;
        RECT 1826.820 1514.690 1826.960 1700.270 ;
        RECT 1827.670 1700.000 1827.950 1700.270 ;
        RECT 1826.760 1514.370 1827.020 1514.690 ;
        RECT 2497.900 1514.370 2498.160 1514.690 ;
        RECT 2497.960 16.730 2498.100 1514.370 ;
        RECT 2497.960 16.590 2500.860 16.730 ;
        RECT 2500.720 2.400 2500.860 16.590 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 0.300 ;
=======
      LAYER li1 ;
        RECT 1847.965 1684.445 1848.135 1685.635 ;
        RECT 1866.365 1684.445 1869.755 1684.615 ;
        RECT 1869.585 1683.765 1869.755 1684.445 ;
        RECT 1938.585 1683.765 1939.675 1683.935 ;
      LAYER mcon ;
        RECT 1847.965 1685.465 1848.135 1685.635 ;
        RECT 1939.505 1683.765 1939.675 1683.935 ;
      LAYER met1 ;
        RECT 1829.950 1685.620 1830.270 1685.680 ;
        RECT 1847.905 1685.620 1848.195 1685.665 ;
        RECT 1829.950 1685.480 1848.195 1685.620 ;
        RECT 1829.950 1685.420 1830.270 1685.480 ;
        RECT 1847.905 1685.435 1848.195 1685.480 ;
        RECT 1847.905 1684.600 1848.195 1684.645 ;
        RECT 1866.305 1684.600 1866.595 1684.645 ;
        RECT 1847.905 1684.460 1866.595 1684.600 ;
        RECT 1847.905 1684.415 1848.195 1684.460 ;
        RECT 1866.305 1684.415 1866.595 1684.460 ;
        RECT 1869.525 1683.920 1869.815 1683.965 ;
        RECT 1938.525 1683.920 1938.815 1683.965 ;
        RECT 1869.525 1683.780 1938.815 1683.920 ;
        RECT 1869.525 1683.735 1869.815 1683.780 ;
        RECT 1938.525 1683.735 1938.815 1683.780 ;
        RECT 1939.445 1683.920 1939.735 1683.965 ;
        RECT 1969.790 1683.920 1970.110 1683.980 ;
        RECT 1939.445 1683.780 1970.110 1683.920 ;
        RECT 1939.445 1683.735 1939.735 1683.780 ;
        RECT 1969.790 1683.720 1970.110 1683.780 ;
        RECT 1969.790 15.200 1970.110 15.260 ;
        RECT 2518.110 15.200 2518.430 15.260 ;
        RECT 1969.790 15.060 2518.430 15.200 ;
        RECT 1969.790 15.000 1970.110 15.060 ;
        RECT 2518.110 15.000 2518.430 15.060 ;
      LAYER via ;
        RECT 1829.980 1685.420 1830.240 1685.680 ;
        RECT 1969.820 1683.720 1970.080 1683.980 ;
        RECT 1969.820 15.000 1970.080 15.260 ;
        RECT 2518.140 15.000 2518.400 15.260 ;
      LAYER met2 ;
        RECT 1829.970 1700.000 1830.250 1704.000 ;
        RECT 1830.040 1685.710 1830.180 1700.000 ;
        RECT 1829.980 1685.390 1830.240 1685.710 ;
        RECT 1969.820 1683.690 1970.080 1684.010 ;
        RECT 1969.880 15.290 1970.020 1683.690 ;
        RECT 1969.820 14.970 1970.080 15.290 ;
        RECT 2518.140 14.970 2518.400 15.290 ;
        RECT 2518.200 2.400 2518.340 14.970 ;
=======
      LAYER met1 ;
        RECT 1832.710 1684.260 1833.030 1684.320 ;
        RECT 1835.010 1684.260 1835.330 1684.320 ;
        RECT 1832.710 1684.120 1835.330 1684.260 ;
        RECT 1832.710 1684.060 1833.030 1684.120 ;
        RECT 1835.010 1684.060 1835.330 1684.120 ;
        RECT 1835.010 79.460 1835.330 79.520 ;
        RECT 2512.130 79.460 2512.450 79.520 ;
        RECT 1835.010 79.320 2512.450 79.460 ;
        RECT 1835.010 79.260 1835.330 79.320 ;
        RECT 2512.130 79.260 2512.450 79.320 ;
        RECT 2512.130 19.280 2512.450 19.340 ;
        RECT 2518.110 19.280 2518.430 19.340 ;
        RECT 2512.130 19.140 2518.430 19.280 ;
        RECT 2512.130 19.080 2512.450 19.140 ;
        RECT 2518.110 19.080 2518.430 19.140 ;
      LAYER via ;
        RECT 1832.740 1684.060 1833.000 1684.320 ;
        RECT 1835.040 1684.060 1835.300 1684.320 ;
        RECT 1835.040 79.260 1835.300 79.520 ;
        RECT 2512.160 79.260 2512.420 79.520 ;
        RECT 2512.160 19.080 2512.420 19.340 ;
        RECT 2518.140 19.080 2518.400 19.340 ;
      LAYER met2 ;
        RECT 1832.730 1700.000 1833.010 1704.000 ;
        RECT 1832.800 1684.350 1832.940 1700.000 ;
        RECT 1832.740 1684.030 1833.000 1684.350 ;
        RECT 1835.040 1684.030 1835.300 1684.350 ;
        RECT 1835.100 79.550 1835.240 1684.030 ;
        RECT 1835.040 79.230 1835.300 79.550 ;
        RECT 2512.160 79.230 2512.420 79.550 ;
        RECT 2512.220 19.370 2512.360 79.230 ;
        RECT 2512.160 19.050 2512.420 19.370 ;
        RECT 2518.140 19.050 2518.400 19.370 ;
        RECT 2518.200 2.400 2518.340 19.050 ;
>>>>>>> re-updated local openlane
        RECT 2517.990 -4.800 2518.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2535.930 -4.800 2536.490 0.300 ;
=======
        RECT 1834.570 1700.410 1834.850 1704.000 ;
        RECT 1834.570 1700.270 1835.240 1700.410 ;
        RECT 1834.570 1700.000 1834.850 1700.270 ;
        RECT 1835.100 19.565 1835.240 1700.270 ;
        RECT 1835.030 19.195 1835.310 19.565 ;
        RECT 2536.070 19.195 2536.350 19.565 ;
        RECT 2536.140 2.400 2536.280 19.195 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
      LAYER via2 ;
        RECT 1835.030 19.240 1835.310 19.520 ;
        RECT 2536.070 19.240 2536.350 19.520 ;
      LAYER met3 ;
        RECT 1835.005 19.530 1835.335 19.545 ;
        RECT 2536.045 19.530 2536.375 19.545 ;
        RECT 1835.005 19.230 2536.375 19.530 ;
        RECT 1835.005 19.215 1835.335 19.230 ;
        RECT 2536.045 19.215 2536.375 19.230 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1837.310 1684.260 1837.630 1684.320 ;
        RECT 1841.910 1684.260 1842.230 1684.320 ;
        RECT 1837.310 1684.120 1842.230 1684.260 ;
        RECT 1837.310 1684.060 1837.630 1684.120 ;
        RECT 1841.910 1684.060 1842.230 1684.120 ;
        RECT 1841.910 1507.460 1842.230 1507.520 ;
        RECT 2532.370 1507.460 2532.690 1507.520 ;
        RECT 1841.910 1507.320 2532.690 1507.460 ;
        RECT 1841.910 1507.260 1842.230 1507.320 ;
        RECT 2532.370 1507.260 2532.690 1507.320 ;
        RECT 2532.370 62.120 2532.690 62.180 ;
        RECT 2536.050 62.120 2536.370 62.180 ;
        RECT 2532.370 61.980 2536.370 62.120 ;
        RECT 2532.370 61.920 2532.690 61.980 ;
        RECT 2536.050 61.920 2536.370 61.980 ;
      LAYER via ;
        RECT 1837.340 1684.060 1837.600 1684.320 ;
        RECT 1841.940 1684.060 1842.200 1684.320 ;
        RECT 1841.940 1507.260 1842.200 1507.520 ;
        RECT 2532.400 1507.260 2532.660 1507.520 ;
        RECT 2532.400 61.920 2532.660 62.180 ;
        RECT 2536.080 61.920 2536.340 62.180 ;
      LAYER met2 ;
        RECT 1837.330 1700.000 1837.610 1704.000 ;
        RECT 1837.400 1684.350 1837.540 1700.000 ;
        RECT 1837.340 1684.030 1837.600 1684.350 ;
        RECT 1841.940 1684.030 1842.200 1684.350 ;
        RECT 1842.000 1507.550 1842.140 1684.030 ;
        RECT 1841.940 1507.230 1842.200 1507.550 ;
        RECT 2532.400 1507.230 2532.660 1507.550 ;
        RECT 2532.460 62.210 2532.600 1507.230 ;
        RECT 2532.400 61.890 2532.660 62.210 ;
        RECT 2536.080 61.890 2536.340 62.210 ;
        RECT 2536.140 2.400 2536.280 61.890 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 0.300 ;
=======
      LAYER li1 ;
        RECT 1848.885 1683.765 1849.055 1685.975 ;
        RECT 1870.505 1683.085 1870.675 1684.615 ;
      LAYER mcon ;
        RECT 1848.885 1685.805 1849.055 1685.975 ;
        RECT 1870.505 1684.445 1870.675 1684.615 ;
      LAYER met1 ;
        RECT 1839.610 1685.960 1839.930 1686.020 ;
        RECT 1848.825 1685.960 1849.115 1686.005 ;
        RECT 1839.610 1685.820 1849.115 1685.960 ;
        RECT 1839.610 1685.760 1839.930 1685.820 ;
        RECT 1848.825 1685.775 1849.115 1685.820 ;
        RECT 1870.445 1684.600 1870.735 1684.645 ;
        RECT 2004.290 1684.600 2004.610 1684.660 ;
        RECT 1870.445 1684.460 2004.610 1684.600 ;
        RECT 1870.445 1684.415 1870.735 1684.460 ;
        RECT 2004.290 1684.400 2004.610 1684.460 ;
        RECT 1848.825 1683.920 1849.115 1683.965 ;
        RECT 1848.825 1683.780 1869.280 1683.920 ;
        RECT 1848.825 1683.735 1849.115 1683.780 ;
        RECT 1869.140 1683.240 1869.280 1683.780 ;
        RECT 1870.445 1683.240 1870.735 1683.285 ;
        RECT 1869.140 1683.100 1870.735 1683.240 ;
        RECT 1870.445 1683.055 1870.735 1683.100 ;
        RECT 2004.290 15.540 2004.610 15.600 ;
        RECT 2553.990 15.540 2554.310 15.600 ;
        RECT 2004.290 15.400 2554.310 15.540 ;
        RECT 2004.290 15.340 2004.610 15.400 ;
        RECT 2553.990 15.340 2554.310 15.400 ;
      LAYER via ;
        RECT 1839.640 1685.760 1839.900 1686.020 ;
        RECT 2004.320 1684.400 2004.580 1684.660 ;
        RECT 2004.320 15.340 2004.580 15.600 ;
        RECT 2554.020 15.340 2554.280 15.600 ;
      LAYER met2 ;
        RECT 1839.630 1700.000 1839.910 1704.000 ;
        RECT 1839.700 1686.050 1839.840 1700.000 ;
        RECT 1839.640 1685.730 1839.900 1686.050 ;
        RECT 2004.320 1684.370 2004.580 1684.690 ;
        RECT 2004.380 15.630 2004.520 1684.370 ;
        RECT 2004.320 15.310 2004.580 15.630 ;
        RECT 2554.020 15.310 2554.280 15.630 ;
        RECT 2554.080 2.400 2554.220 15.310 ;
=======
      LAYER met1 ;
        RECT 1842.370 1683.920 1842.690 1683.980 ;
        RECT 1847.430 1683.920 1847.750 1683.980 ;
        RECT 1842.370 1683.780 1847.750 1683.920 ;
        RECT 1842.370 1683.720 1842.690 1683.780 ;
        RECT 1847.430 1683.720 1847.750 1683.780 ;
        RECT 1847.430 1500.660 1847.750 1500.720 ;
        RECT 2553.070 1500.660 2553.390 1500.720 ;
        RECT 1847.430 1500.520 2553.390 1500.660 ;
        RECT 1847.430 1500.460 1847.750 1500.520 ;
        RECT 2553.070 1500.460 2553.390 1500.520 ;
      LAYER via ;
        RECT 1842.400 1683.720 1842.660 1683.980 ;
        RECT 1847.460 1683.720 1847.720 1683.980 ;
        RECT 1847.460 1500.460 1847.720 1500.720 ;
        RECT 2553.100 1500.460 2553.360 1500.720 ;
      LAYER met2 ;
        RECT 1842.390 1700.000 1842.670 1704.000 ;
        RECT 1842.460 1684.010 1842.600 1700.000 ;
        RECT 1842.400 1683.690 1842.660 1684.010 ;
        RECT 1847.460 1683.690 1847.720 1684.010 ;
        RECT 1847.520 1500.750 1847.660 1683.690 ;
        RECT 1847.460 1500.430 1847.720 1500.750 ;
        RECT 2553.100 1500.430 2553.360 1500.750 ;
        RECT 2553.160 61.610 2553.300 1500.430 ;
        RECT 2553.160 61.470 2554.220 61.610 ;
        RECT 2554.080 2.400 2554.220 61.470 ;
>>>>>>> re-updated local openlane
        RECT 2553.870 -4.800 2554.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 0.300 ;
=======
      LAYER met1 ;
        RECT 1847.890 1479.920 1848.210 1479.980 ;
        RECT 2566.870 1479.920 2567.190 1479.980 ;
        RECT 1847.890 1479.780 2567.190 1479.920 ;
        RECT 1847.890 1479.720 1848.210 1479.780 ;
        RECT 2566.870 1479.720 2567.190 1479.780 ;
        RECT 2566.870 62.120 2567.190 62.180 ;
        RECT 2571.930 62.120 2572.250 62.180 ;
        RECT 2566.870 61.980 2572.250 62.120 ;
        RECT 2566.870 61.920 2567.190 61.980 ;
        RECT 2571.930 61.920 2572.250 61.980 ;
      LAYER via ;
        RECT 1847.920 1479.720 1848.180 1479.980 ;
        RECT 2566.900 1479.720 2567.160 1479.980 ;
        RECT 2566.900 61.920 2567.160 62.180 ;
        RECT 2571.960 61.920 2572.220 62.180 ;
      LAYER met2 ;
        RECT 1846.990 1700.410 1847.270 1704.000 ;
        RECT 1846.990 1700.270 1848.120 1700.410 ;
        RECT 1846.990 1700.000 1847.270 1700.270 ;
        RECT 1847.980 1480.010 1848.120 1700.270 ;
        RECT 1847.920 1479.690 1848.180 1480.010 ;
        RECT 2566.900 1479.690 2567.160 1480.010 ;
        RECT 2566.960 62.210 2567.100 1479.690 ;
        RECT 2566.900 61.890 2567.160 62.210 ;
        RECT 2571.960 61.890 2572.220 62.210 ;
        RECT 2572.020 2.400 2572.160 61.890 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 0.300 ;
=======
      LAYER li1 ;
        RECT 2587.645 766.105 2587.815 814.215 ;
        RECT 2587.645 669.545 2587.815 717.655 ;
        RECT 2587.645 572.645 2587.815 620.755 ;
        RECT 2587.645 476.085 2587.815 524.195 ;
        RECT 2587.645 282.965 2587.815 331.075 ;
        RECT 2587.645 186.405 2587.815 234.515 ;
        RECT 2587.645 89.845 2587.815 137.955 ;
      LAYER mcon ;
        RECT 2587.645 814.045 2587.815 814.215 ;
        RECT 2587.645 717.485 2587.815 717.655 ;
        RECT 2587.645 620.585 2587.815 620.755 ;
        RECT 2587.645 524.025 2587.815 524.195 ;
        RECT 2587.645 330.905 2587.815 331.075 ;
        RECT 2587.645 234.345 2587.815 234.515 ;
        RECT 2587.645 137.785 2587.815 137.955 ;
      LAYER met1 ;
        RECT 1852.030 1684.940 1852.350 1685.000 ;
        RECT 1855.250 1684.940 1855.570 1685.000 ;
        RECT 1852.030 1684.800 1855.570 1684.940 ;
        RECT 1852.030 1684.740 1852.350 1684.800 ;
        RECT 1855.250 1684.740 1855.570 1684.800 ;
        RECT 1855.250 886.620 1855.570 886.680 ;
        RECT 2587.570 886.620 2587.890 886.680 ;
        RECT 1855.250 886.480 2587.890 886.620 ;
        RECT 1855.250 886.420 1855.570 886.480 ;
        RECT 2587.570 886.420 2587.890 886.480 ;
        RECT 2587.570 814.200 2587.890 814.260 ;
        RECT 2587.375 814.060 2587.890 814.200 ;
        RECT 2587.570 814.000 2587.890 814.060 ;
        RECT 2587.570 766.260 2587.890 766.320 ;
        RECT 2587.375 766.120 2587.890 766.260 ;
        RECT 2587.570 766.060 2587.890 766.120 ;
        RECT 2587.570 717.640 2587.890 717.700 ;
        RECT 2587.375 717.500 2587.890 717.640 ;
        RECT 2587.570 717.440 2587.890 717.500 ;
        RECT 2587.570 669.700 2587.890 669.760 ;
        RECT 2587.375 669.560 2587.890 669.700 ;
        RECT 2587.570 669.500 2587.890 669.560 ;
        RECT 2587.570 620.740 2587.890 620.800 ;
        RECT 2587.375 620.600 2587.890 620.740 ;
        RECT 2587.570 620.540 2587.890 620.600 ;
        RECT 2587.570 572.800 2587.890 572.860 ;
        RECT 2587.375 572.660 2587.890 572.800 ;
        RECT 2587.570 572.600 2587.890 572.660 ;
        RECT 2587.570 524.180 2587.890 524.240 ;
        RECT 2587.375 524.040 2587.890 524.180 ;
        RECT 2587.570 523.980 2587.890 524.040 ;
        RECT 2587.570 476.240 2587.890 476.300 ;
        RECT 2587.375 476.100 2587.890 476.240 ;
        RECT 2587.570 476.040 2587.890 476.100 ;
        RECT 2587.570 331.060 2587.890 331.120 ;
        RECT 2587.375 330.920 2587.890 331.060 ;
        RECT 2587.570 330.860 2587.890 330.920 ;
        RECT 2587.570 283.120 2587.890 283.180 ;
        RECT 2587.375 282.980 2587.890 283.120 ;
        RECT 2587.570 282.920 2587.890 282.980 ;
        RECT 2587.570 234.500 2587.890 234.560 ;
        RECT 2587.375 234.360 2587.890 234.500 ;
        RECT 2587.570 234.300 2587.890 234.360 ;
        RECT 2587.570 186.560 2587.890 186.620 ;
        RECT 2587.375 186.420 2587.890 186.560 ;
        RECT 2587.570 186.360 2587.890 186.420 ;
        RECT 2587.570 137.940 2587.890 138.000 ;
        RECT 2587.375 137.800 2587.890 137.940 ;
        RECT 2587.570 137.740 2587.890 137.800 ;
        RECT 2587.570 90.000 2587.890 90.060 ;
        RECT 2587.375 89.860 2587.890 90.000 ;
        RECT 2587.570 89.800 2587.890 89.860 ;
        RECT 2587.570 62.260 2587.890 62.520 ;
        RECT 2587.660 61.780 2587.800 62.260 ;
        RECT 2589.410 61.780 2589.730 61.840 ;
        RECT 2587.660 61.640 2589.730 61.780 ;
        RECT 2589.410 61.580 2589.730 61.640 ;
        RECT 2589.410 47.980 2589.730 48.240 ;
        RECT 2589.500 47.560 2589.640 47.980 ;
        RECT 2589.410 47.300 2589.730 47.560 ;
      LAYER via ;
        RECT 1852.060 1684.740 1852.320 1685.000 ;
        RECT 1855.280 1684.740 1855.540 1685.000 ;
        RECT 1855.280 886.420 1855.540 886.680 ;
        RECT 2587.600 886.420 2587.860 886.680 ;
        RECT 2587.600 814.000 2587.860 814.260 ;
        RECT 2587.600 766.060 2587.860 766.320 ;
        RECT 2587.600 717.440 2587.860 717.700 ;
        RECT 2587.600 669.500 2587.860 669.760 ;
        RECT 2587.600 620.540 2587.860 620.800 ;
        RECT 2587.600 572.600 2587.860 572.860 ;
        RECT 2587.600 523.980 2587.860 524.240 ;
        RECT 2587.600 476.040 2587.860 476.300 ;
        RECT 2587.600 330.860 2587.860 331.120 ;
        RECT 2587.600 282.920 2587.860 283.180 ;
        RECT 2587.600 234.300 2587.860 234.560 ;
        RECT 2587.600 186.360 2587.860 186.620 ;
        RECT 2587.600 137.740 2587.860 138.000 ;
        RECT 2587.600 89.800 2587.860 90.060 ;
        RECT 2587.600 62.260 2587.860 62.520 ;
        RECT 2589.440 61.580 2589.700 61.840 ;
        RECT 2589.440 47.980 2589.700 48.240 ;
        RECT 2589.440 47.300 2589.700 47.560 ;
      LAYER met2 ;
        RECT 1852.050 1700.000 1852.330 1704.000 ;
        RECT 1852.120 1685.030 1852.260 1700.000 ;
        RECT 1852.060 1684.710 1852.320 1685.030 ;
        RECT 1855.280 1684.710 1855.540 1685.030 ;
        RECT 1855.340 886.710 1855.480 1684.710 ;
        RECT 1855.280 886.390 1855.540 886.710 ;
        RECT 2587.600 886.390 2587.860 886.710 ;
        RECT 2587.660 821.965 2587.800 886.390 ;
        RECT 2587.590 821.595 2587.870 821.965 ;
        RECT 2587.590 820.915 2587.870 821.285 ;
        RECT 2587.660 814.290 2587.800 820.915 ;
        RECT 2587.600 813.970 2587.860 814.290 ;
        RECT 2587.600 766.030 2587.860 766.350 ;
        RECT 2587.660 717.730 2587.800 766.030 ;
        RECT 2587.600 717.410 2587.860 717.730 ;
        RECT 2587.600 669.470 2587.860 669.790 ;
        RECT 2587.660 620.830 2587.800 669.470 ;
        RECT 2587.600 620.510 2587.860 620.830 ;
        RECT 2587.600 572.570 2587.860 572.890 ;
        RECT 2587.660 524.270 2587.800 572.570 ;
        RECT 2587.600 523.950 2587.860 524.270 ;
        RECT 2587.600 476.010 2587.860 476.330 ;
        RECT 2587.660 331.150 2587.800 476.010 ;
        RECT 2587.600 330.830 2587.860 331.150 ;
        RECT 2587.600 282.890 2587.860 283.210 ;
        RECT 2587.660 234.590 2587.800 282.890 ;
        RECT 2587.600 234.270 2587.860 234.590 ;
        RECT 2587.600 186.330 2587.860 186.650 ;
        RECT 2587.660 138.030 2587.800 186.330 ;
        RECT 2587.600 137.710 2587.860 138.030 ;
        RECT 2587.600 89.770 2587.860 90.090 ;
        RECT 2587.660 62.550 2587.800 89.770 ;
        RECT 2587.600 62.230 2587.860 62.550 ;
        RECT 2589.440 61.550 2589.700 61.870 ;
        RECT 2589.500 48.270 2589.640 61.550 ;
        RECT 2589.440 47.950 2589.700 48.270 ;
        RECT 2589.440 47.270 2589.700 47.590 ;
        RECT 2589.500 2.400 2589.640 47.270 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 2587.590 821.640 2587.870 821.920 ;
        RECT 2587.590 820.960 2587.870 821.240 ;
      LAYER met3 ;
        RECT 2587.565 821.930 2587.895 821.945 ;
        RECT 2587.565 821.630 2588.570 821.930 ;
        RECT 2587.565 821.615 2587.895 821.630 ;
        RECT 2587.565 821.250 2587.895 821.265 ;
        RECT 2588.270 821.250 2588.570 821.630 ;
        RECT 2587.565 820.950 2588.570 821.250 ;
        RECT 2587.565 820.935 2587.895 820.950 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1367.190 1678.140 1367.510 1678.200 ;
        RECT 1371.790 1678.140 1372.110 1678.200 ;
        RECT 1367.190 1678.000 1372.110 1678.140 ;
        RECT 1367.190 1677.940 1367.510 1678.000 ;
        RECT 1371.790 1677.940 1372.110 1678.000 ;
        RECT 823.470 37.640 823.790 37.700 ;
        RECT 1367.190 37.640 1367.510 37.700 ;
        RECT 823.470 37.500 1367.510 37.640 ;
        RECT 823.470 37.440 823.790 37.500 ;
        RECT 1367.190 37.440 1367.510 37.500 ;
      LAYER via ;
        RECT 1367.220 1677.940 1367.480 1678.200 ;
        RECT 1371.820 1677.940 1372.080 1678.200 ;
        RECT 823.500 37.440 823.760 37.700 ;
        RECT 1367.220 37.440 1367.480 37.700 ;
      LAYER met2 ;
        RECT 1372.730 1700.410 1373.010 1704.000 ;
        RECT 1371.880 1700.270 1373.010 1700.410 ;
        RECT 1371.880 1678.230 1372.020 1700.270 ;
        RECT 1372.730 1700.000 1373.010 1700.270 ;
        RECT 1367.220 1677.910 1367.480 1678.230 ;
        RECT 1371.820 1677.910 1372.080 1678.230 ;
        RECT 1367.280 37.730 1367.420 1677.910 ;
        RECT 823.500 37.410 823.760 37.730 ;
        RECT 1367.220 37.410 1367.480 37.730 ;
        RECT 823.560 2.400 823.700 37.410 ;
        RECT 823.350 -4.800 823.910 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1200.690 40.320 1200.970 40.600 ;
        RECT 1203.450 40.320 1203.730 40.600 ;
      LAYER met3 ;
        RECT 1200.665 40.610 1200.995 40.625 ;
        RECT 1203.425 40.610 1203.755 40.625 ;
        RECT 1200.665 40.310 1203.755 40.610 ;
        RECT 1200.665 40.295 1200.995 40.310 ;
        RECT 1203.425 40.295 1203.755 40.310 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 0.300 ;
=======
      LAYER li1 ;
        RECT 1858.545 17.085 1858.715 18.955 ;
      LAYER mcon ;
        RECT 1858.545 18.785 1858.715 18.955 ;
      LAYER met1 ;
        RECT 1853.870 1686.640 1854.190 1686.700 ;
        RECT 1855.710 1686.640 1856.030 1686.700 ;
        RECT 1853.870 1686.500 1856.030 1686.640 ;
        RECT 1853.870 1686.440 1854.190 1686.500 ;
        RECT 1855.710 1686.440 1856.030 1686.500 ;
        RECT 1855.710 18.940 1856.030 19.000 ;
        RECT 1858.485 18.940 1858.775 18.985 ;
        RECT 1855.710 18.800 1858.775 18.940 ;
        RECT 1855.710 18.740 1856.030 18.800 ;
        RECT 1858.485 18.755 1858.775 18.800 ;
        RECT 2607.350 17.580 2607.670 17.640 ;
        RECT 1873.740 17.440 2607.670 17.580 ;
        RECT 1858.485 17.240 1858.775 17.285 ;
        RECT 1873.740 17.240 1873.880 17.440 ;
        RECT 2607.350 17.380 2607.670 17.440 ;
        RECT 1858.485 17.100 1873.880 17.240 ;
        RECT 1858.485 17.055 1858.775 17.100 ;
      LAYER via ;
        RECT 1853.900 1686.440 1854.160 1686.700 ;
        RECT 1855.740 1686.440 1856.000 1686.700 ;
        RECT 1855.740 18.740 1856.000 19.000 ;
        RECT 2607.380 17.380 2607.640 17.640 ;
      LAYER met2 ;
        RECT 1853.890 1700.000 1854.170 1704.000 ;
        RECT 1853.960 1686.730 1854.100 1700.000 ;
        RECT 1853.900 1686.410 1854.160 1686.730 ;
        RECT 1855.740 1686.410 1856.000 1686.730 ;
        RECT 1855.800 19.030 1855.940 1686.410 ;
        RECT 1855.740 18.710 1856.000 19.030 ;
        RECT 2607.380 17.350 2607.640 17.670 ;
        RECT 2607.440 2.400 2607.580 17.350 ;
=======
      LAYER met1 ;
        RECT 1856.630 1666.240 1856.950 1666.300 ;
        RECT 2601.370 1666.240 2601.690 1666.300 ;
        RECT 1856.630 1666.100 2601.690 1666.240 ;
        RECT 1856.630 1666.040 1856.950 1666.100 ;
        RECT 2601.370 1666.040 2601.690 1666.100 ;
        RECT 2601.370 36.280 2601.690 36.340 ;
        RECT 2607.350 36.280 2607.670 36.340 ;
        RECT 2601.370 36.140 2607.670 36.280 ;
        RECT 2601.370 36.080 2601.690 36.140 ;
        RECT 2607.350 36.080 2607.670 36.140 ;
      LAYER via ;
        RECT 1856.660 1666.040 1856.920 1666.300 ;
        RECT 2601.400 1666.040 2601.660 1666.300 ;
        RECT 2601.400 36.080 2601.660 36.340 ;
        RECT 2607.380 36.080 2607.640 36.340 ;
      LAYER met2 ;
        RECT 1856.650 1700.000 1856.930 1704.000 ;
        RECT 1856.720 1666.330 1856.860 1700.000 ;
        RECT 1856.660 1666.010 1856.920 1666.330 ;
        RECT 2601.400 1666.010 2601.660 1666.330 ;
        RECT 2601.460 36.370 2601.600 1666.010 ;
        RECT 2601.400 36.050 2601.660 36.370 ;
        RECT 2607.380 36.050 2607.640 36.370 ;
        RECT 2607.440 2.400 2607.580 36.050 ;
>>>>>>> re-updated local openlane
        RECT 2607.230 -4.800 2607.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 0.300 ;
=======
      LAYER li1 ;
        RECT 1869.125 1685.125 1869.295 1686.655 ;
        RECT 1870.505 1685.125 1870.675 1686.655 ;
        RECT 2087.165 16.405 2087.335 18.615 ;
      LAYER mcon ;
        RECT 1869.125 1686.485 1869.295 1686.655 ;
        RECT 1870.505 1686.485 1870.675 1686.655 ;
        RECT 2087.165 18.445 2087.335 18.615 ;
      LAYER met1 ;
        RECT 1869.065 1686.640 1869.355 1686.685 ;
        RECT 1870.445 1686.640 1870.735 1686.685 ;
        RECT 1869.065 1686.500 1870.735 1686.640 ;
        RECT 1869.065 1686.455 1869.355 1686.500 ;
        RECT 1870.445 1686.455 1870.735 1686.500 ;
        RECT 1858.470 1685.280 1858.790 1685.340 ;
        RECT 1869.065 1685.280 1869.355 1685.325 ;
        RECT 1858.470 1685.140 1869.355 1685.280 ;
        RECT 1858.470 1685.080 1858.790 1685.140 ;
        RECT 1869.065 1685.095 1869.355 1685.140 ;
        RECT 1870.445 1685.095 1870.735 1685.325 ;
        RECT 2038.790 1685.280 2039.110 1685.340 ;
        RECT 1890.760 1685.140 2039.110 1685.280 ;
        RECT 1870.520 1684.940 1870.660 1685.095 ;
        RECT 1890.760 1684.940 1890.900 1685.140 ;
        RECT 2038.790 1685.080 2039.110 1685.140 ;
        RECT 1870.520 1684.800 1890.900 1684.940 ;
        RECT 2039.250 18.600 2039.570 18.660 ;
        RECT 2087.105 18.600 2087.395 18.645 ;
        RECT 2039.250 18.460 2087.395 18.600 ;
        RECT 2039.250 18.400 2039.570 18.460 ;
        RECT 2087.105 18.415 2087.395 18.460 ;
        RECT 2087.105 16.560 2087.395 16.605 ;
        RECT 2625.290 16.560 2625.610 16.620 ;
        RECT 2087.105 16.420 2625.610 16.560 ;
        RECT 2087.105 16.375 2087.395 16.420 ;
        RECT 2625.290 16.360 2625.610 16.420 ;
      LAYER via ;
        RECT 1858.500 1685.080 1858.760 1685.340 ;
        RECT 2038.820 1685.080 2039.080 1685.340 ;
        RECT 2039.280 18.400 2039.540 18.660 ;
        RECT 2625.320 16.360 2625.580 16.620 ;
      LAYER met2 ;
        RECT 1858.490 1700.000 1858.770 1704.000 ;
        RECT 1858.560 1685.370 1858.700 1700.000 ;
        RECT 1858.500 1685.050 1858.760 1685.370 ;
        RECT 2038.820 1685.050 2039.080 1685.370 ;
        RECT 2038.880 18.770 2039.020 1685.050 ;
        RECT 2038.880 18.690 2039.480 18.770 ;
        RECT 2038.880 18.630 2039.540 18.690 ;
        RECT 2039.280 18.370 2039.540 18.630 ;
        RECT 2625.320 16.330 2625.580 16.650 ;
        RECT 2625.380 2.400 2625.520 16.330 ;
=======
      LAYER met1 ;
        RECT 1858.470 1683.920 1858.790 1683.980 ;
        RECT 1861.690 1683.920 1862.010 1683.980 ;
        RECT 1858.470 1683.780 1862.010 1683.920 ;
        RECT 1858.470 1683.720 1858.790 1683.780 ;
        RECT 1861.690 1683.720 1862.010 1683.780 ;
        RECT 1858.470 1645.500 1858.790 1645.560 ;
        RECT 2622.070 1645.500 2622.390 1645.560 ;
        RECT 1858.470 1645.360 2622.390 1645.500 ;
        RECT 1858.470 1645.300 1858.790 1645.360 ;
        RECT 2622.070 1645.300 2622.390 1645.360 ;
        RECT 2622.070 72.660 2622.390 72.720 ;
        RECT 2625.290 72.660 2625.610 72.720 ;
        RECT 2622.070 72.520 2625.610 72.660 ;
        RECT 2622.070 72.460 2622.390 72.520 ;
        RECT 2625.290 72.460 2625.610 72.520 ;
      LAYER via ;
        RECT 1858.500 1683.720 1858.760 1683.980 ;
        RECT 1861.720 1683.720 1861.980 1683.980 ;
        RECT 1858.500 1645.300 1858.760 1645.560 ;
        RECT 2622.100 1645.300 2622.360 1645.560 ;
        RECT 2622.100 72.460 2622.360 72.720 ;
        RECT 2625.320 72.460 2625.580 72.720 ;
      LAYER met2 ;
        RECT 1861.710 1700.000 1861.990 1704.000 ;
        RECT 1861.780 1684.010 1861.920 1700.000 ;
        RECT 1858.500 1683.690 1858.760 1684.010 ;
        RECT 1861.720 1683.690 1861.980 1684.010 ;
        RECT 1858.560 1645.590 1858.700 1683.690 ;
        RECT 1858.500 1645.270 1858.760 1645.590 ;
        RECT 2622.100 1645.270 2622.360 1645.590 ;
        RECT 2622.160 72.750 2622.300 1645.270 ;
        RECT 2622.100 72.430 2622.360 72.750 ;
        RECT 2625.320 72.430 2625.580 72.750 ;
        RECT 2625.380 2.400 2625.520 72.430 ;
>>>>>>> re-updated local openlane
        RECT 2625.170 -4.800 2625.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1863.530 1686.640 1863.850 1686.700 ;
        RECT 1868.590 1686.640 1868.910 1686.700 ;
        RECT 1863.530 1686.500 1868.910 1686.640 ;
        RECT 1863.530 1686.440 1863.850 1686.500 ;
        RECT 1868.590 1686.440 1868.910 1686.500 ;
        RECT 1868.590 51.920 1868.910 51.980 ;
        RECT 2642.770 51.920 2643.090 51.980 ;
        RECT 1868.590 51.780 2643.090 51.920 ;
        RECT 1868.590 51.720 1868.910 51.780 ;
        RECT 2642.770 51.720 2643.090 51.780 ;
      LAYER via ;
        RECT 1863.560 1686.440 1863.820 1686.700 ;
        RECT 1868.620 1686.440 1868.880 1686.700 ;
        RECT 1868.620 51.720 1868.880 51.980 ;
        RECT 2642.800 51.720 2643.060 51.980 ;
      LAYER met2 ;
        RECT 1863.550 1700.000 1863.830 1704.000 ;
        RECT 1863.620 1686.730 1863.760 1700.000 ;
        RECT 1863.560 1686.410 1863.820 1686.730 ;
        RECT 1868.620 1686.410 1868.880 1686.730 ;
        RECT 1868.680 52.010 1868.820 1686.410 ;
        RECT 1868.620 51.690 1868.880 52.010 ;
        RECT 2642.800 51.690 2643.060 52.010 ;
        RECT 2642.860 3.130 2643.000 51.690 ;
        RECT 2642.860 2.990 2643.460 3.130 ;
        RECT 2643.320 2.400 2643.460 2.990 ;
=======
      LAYER li1 ;
        RECT 2642.845 48.365 2643.015 96.475 ;
      LAYER mcon ;
        RECT 2642.845 96.305 2643.015 96.475 ;
      LAYER met1 ;
        RECT 1867.670 1638.700 1867.990 1638.760 ;
        RECT 2642.770 1638.700 2643.090 1638.760 ;
        RECT 1867.670 1638.560 2643.090 1638.700 ;
        RECT 1867.670 1638.500 1867.990 1638.560 ;
        RECT 2642.770 1638.500 2643.090 1638.560 ;
        RECT 2642.770 96.460 2643.090 96.520 ;
        RECT 2642.575 96.320 2643.090 96.460 ;
        RECT 2642.770 96.260 2643.090 96.320 ;
        RECT 2642.785 48.520 2643.075 48.565 ;
        RECT 2643.230 48.520 2643.550 48.580 ;
        RECT 2642.785 48.380 2643.550 48.520 ;
        RECT 2642.785 48.335 2643.075 48.380 ;
        RECT 2643.230 48.320 2643.550 48.380 ;
        RECT 2643.230 2.960 2643.550 3.020 ;
        RECT 2643.690 2.960 2644.010 3.020 ;
        RECT 2643.230 2.820 2644.010 2.960 ;
        RECT 2643.230 2.760 2643.550 2.820 ;
        RECT 2643.690 2.760 2644.010 2.820 ;
      LAYER via ;
        RECT 1867.700 1638.500 1867.960 1638.760 ;
        RECT 2642.800 1638.500 2643.060 1638.760 ;
        RECT 2642.800 96.260 2643.060 96.520 ;
        RECT 2643.260 48.320 2643.520 48.580 ;
        RECT 2643.260 2.760 2643.520 3.020 ;
        RECT 2643.720 2.760 2643.980 3.020 ;
      LAYER met2 ;
        RECT 1866.310 1700.410 1866.590 1704.000 ;
        RECT 1866.310 1700.270 1867.900 1700.410 ;
        RECT 1866.310 1700.000 1866.590 1700.270 ;
        RECT 1867.760 1638.790 1867.900 1700.270 ;
        RECT 1867.700 1638.470 1867.960 1638.790 ;
        RECT 2642.800 1638.470 2643.060 1638.790 ;
        RECT 2642.860 96.550 2643.000 1638.470 ;
        RECT 2642.800 96.230 2643.060 96.550 ;
        RECT 2643.260 48.290 2643.520 48.610 ;
        RECT 2643.320 48.010 2643.460 48.290 ;
        RECT 2643.320 47.870 2643.920 48.010 ;
        RECT 2643.780 3.050 2643.920 47.870 ;
        RECT 2643.260 2.730 2643.520 3.050 ;
        RECT 2643.720 2.730 2643.980 3.050 ;
        RECT 2643.320 2.400 2643.460 2.730 ;
>>>>>>> re-updated local openlane
        RECT 2643.110 -4.800 2643.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 0.300 ;
=======
      LAYER li1 ;
        RECT 1893.965 1684.785 1894.135 1685.975 ;
      LAYER mcon ;
        RECT 1893.965 1685.805 1894.135 1685.975 ;
      LAYER met1 ;
        RECT 1868.130 1685.960 1868.450 1686.020 ;
        RECT 1893.905 1685.960 1894.195 1686.005 ;
        RECT 1868.130 1685.820 1894.195 1685.960 ;
        RECT 1868.130 1685.760 1868.450 1685.820 ;
        RECT 1893.905 1685.775 1894.195 1685.820 ;
        RECT 1893.905 1684.940 1894.195 1684.985 ;
        RECT 2039.250 1684.940 2039.570 1685.000 ;
        RECT 1893.905 1684.800 2039.570 1684.940 ;
        RECT 1893.905 1684.755 1894.195 1684.800 ;
        RECT 2039.250 1684.740 2039.570 1684.800 ;
        RECT 2054.890 20.300 2055.210 20.360 ;
        RECT 2661.170 20.300 2661.490 20.360 ;
        RECT 2054.890 20.160 2661.490 20.300 ;
        RECT 2054.890 20.100 2055.210 20.160 ;
        RECT 2661.170 20.100 2661.490 20.160 ;
      LAYER via ;
        RECT 1868.160 1685.760 1868.420 1686.020 ;
        RECT 2039.280 1684.740 2039.540 1685.000 ;
        RECT 2054.920 20.100 2055.180 20.360 ;
        RECT 2661.200 20.100 2661.460 20.360 ;
=======
      LAYER met1 ;
        RECT 1871.350 1683.920 1871.670 1683.980 ;
        RECT 1875.030 1683.920 1875.350 1683.980 ;
        RECT 1871.350 1683.780 1875.350 1683.920 ;
        RECT 1871.350 1683.720 1871.670 1683.780 ;
        RECT 1875.030 1683.720 1875.350 1683.780 ;
        RECT 1875.030 1487.060 1875.350 1487.120 ;
        RECT 2656.570 1487.060 2656.890 1487.120 ;
        RECT 1875.030 1486.920 2656.890 1487.060 ;
        RECT 1875.030 1486.860 1875.350 1486.920 ;
        RECT 2656.570 1486.860 2656.890 1486.920 ;
        RECT 2656.570 62.120 2656.890 62.180 ;
        RECT 2661.170 62.120 2661.490 62.180 ;
        RECT 2656.570 61.980 2661.490 62.120 ;
        RECT 2656.570 61.920 2656.890 61.980 ;
        RECT 2661.170 61.920 2661.490 61.980 ;
      LAYER via ;
        RECT 1871.380 1683.720 1871.640 1683.980 ;
        RECT 1875.060 1683.720 1875.320 1683.980 ;
        RECT 1875.060 1486.860 1875.320 1487.120 ;
        RECT 2656.600 1486.860 2656.860 1487.120 ;
        RECT 2656.600 61.920 2656.860 62.180 ;
        RECT 2661.200 61.920 2661.460 62.180 ;
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1871.370 1700.000 1871.650 1704.000 ;
        RECT 1871.440 1684.010 1871.580 1700.000 ;
        RECT 1871.380 1683.690 1871.640 1684.010 ;
        RECT 1875.060 1683.690 1875.320 1684.010 ;
        RECT 1875.120 1487.150 1875.260 1683.690 ;
        RECT 1875.060 1486.830 1875.320 1487.150 ;
        RECT 2656.600 1486.830 2656.860 1487.150 ;
        RECT 2656.660 62.210 2656.800 1486.830 ;
        RECT 2656.600 61.890 2656.860 62.210 ;
        RECT 2661.200 61.890 2661.460 62.210 ;
        RECT 2661.260 2.400 2661.400 61.890 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 2039.270 20.600 2039.550 20.880 ;
        RECT 2054.910 20.600 2055.190 20.880 ;
      LAYER met3 ;
        RECT 2039.245 20.890 2039.575 20.905 ;
        RECT 2054.885 20.890 2055.215 20.905 ;
        RECT 2039.245 20.590 2055.215 20.890 ;
        RECT 2039.245 20.575 2039.575 20.590 ;
        RECT 2054.885 20.575 2055.215 20.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1874.110 1683.580 1874.430 1683.640 ;
        RECT 1876.410 1683.580 1876.730 1683.640 ;
        RECT 1874.110 1683.440 1876.730 1683.580 ;
        RECT 1874.110 1683.380 1874.430 1683.440 ;
        RECT 1876.410 1683.380 1876.730 1683.440 ;
        RECT 1876.410 17.240 1876.730 17.300 ;
        RECT 2678.650 17.240 2678.970 17.300 ;
        RECT 1876.410 17.100 2678.970 17.240 ;
        RECT 1876.410 17.040 1876.730 17.100 ;
        RECT 2678.650 17.040 2678.970 17.100 ;
      LAYER via ;
        RECT 1874.140 1683.380 1874.400 1683.640 ;
        RECT 1876.440 1683.380 1876.700 1683.640 ;
        RECT 1876.440 17.040 1876.700 17.300 ;
        RECT 2678.680 17.040 2678.940 17.300 ;
      LAYER met2 ;
        RECT 1873.210 1700.410 1873.490 1704.000 ;
        RECT 1873.210 1700.270 1874.340 1700.410 ;
        RECT 1873.210 1700.000 1873.490 1700.270 ;
        RECT 1874.200 1683.670 1874.340 1700.270 ;
        RECT 1874.140 1683.350 1874.400 1683.670 ;
        RECT 1876.440 1683.350 1876.700 1683.670 ;
        RECT 1876.500 17.330 1876.640 1683.350 ;
        RECT 1876.440 17.010 1876.700 17.330 ;
        RECT 2678.680 17.010 2678.940 17.330 ;
        RECT 2678.740 2.400 2678.880 17.010 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 2677.345 1442.025 2677.515 1473.135 ;
        RECT 2677.345 766.105 2677.515 814.215 ;
        RECT 2677.345 669.545 2677.515 717.655 ;
        RECT 2677.345 572.645 2677.515 620.755 ;
        RECT 2677.345 476.085 2677.515 524.195 ;
        RECT 2677.345 379.525 2677.515 427.635 ;
        RECT 2677.345 282.965 2677.515 331.075 ;
        RECT 2677.345 186.405 2677.515 234.515 ;
        RECT 2677.345 48.365 2677.515 137.955 ;
      LAYER mcon ;
        RECT 2677.345 1472.965 2677.515 1473.135 ;
        RECT 2677.345 814.045 2677.515 814.215 ;
        RECT 2677.345 717.485 2677.515 717.655 ;
        RECT 2677.345 620.585 2677.515 620.755 ;
        RECT 2677.345 524.025 2677.515 524.195 ;
        RECT 2677.345 427.465 2677.515 427.635 ;
        RECT 2677.345 330.905 2677.515 331.075 ;
        RECT 2677.345 234.345 2677.515 234.515 ;
        RECT 2677.345 137.785 2677.515 137.955 ;
      LAYER met1 ;
        RECT 1875.490 1473.120 1875.810 1473.180 ;
        RECT 2677.285 1473.120 2677.575 1473.165 ;
        RECT 1875.490 1472.980 2677.575 1473.120 ;
        RECT 1875.490 1472.920 1875.810 1472.980 ;
        RECT 2677.285 1472.935 2677.575 1472.980 ;
        RECT 2677.270 1442.180 2677.590 1442.240 ;
        RECT 2677.075 1442.040 2677.590 1442.180 ;
        RECT 2677.270 1441.980 2677.590 1442.040 ;
        RECT 2677.270 1345.620 2677.590 1345.680 ;
        RECT 2678.190 1345.620 2678.510 1345.680 ;
        RECT 2677.270 1345.480 2678.510 1345.620 ;
        RECT 2677.270 1345.420 2677.590 1345.480 ;
        RECT 2678.190 1345.420 2678.510 1345.480 ;
        RECT 2677.270 1249.060 2677.590 1249.120 ;
        RECT 2678.190 1249.060 2678.510 1249.120 ;
        RECT 2677.270 1248.920 2678.510 1249.060 ;
        RECT 2677.270 1248.860 2677.590 1248.920 ;
        RECT 2678.190 1248.860 2678.510 1248.920 ;
        RECT 2677.270 1152.500 2677.590 1152.560 ;
        RECT 2678.190 1152.500 2678.510 1152.560 ;
        RECT 2677.270 1152.360 2678.510 1152.500 ;
        RECT 2677.270 1152.300 2677.590 1152.360 ;
        RECT 2678.190 1152.300 2678.510 1152.360 ;
        RECT 2677.270 1007.320 2677.590 1007.380 ;
        RECT 2678.190 1007.320 2678.510 1007.380 ;
        RECT 2677.270 1007.180 2678.510 1007.320 ;
        RECT 2677.270 1007.120 2677.590 1007.180 ;
        RECT 2678.190 1007.120 2678.510 1007.180 ;
        RECT 2677.270 910.760 2677.590 910.820 ;
        RECT 2678.190 910.760 2678.510 910.820 ;
        RECT 2677.270 910.620 2678.510 910.760 ;
        RECT 2677.270 910.560 2677.590 910.620 ;
        RECT 2678.190 910.560 2678.510 910.620 ;
        RECT 2677.270 814.200 2677.590 814.260 ;
        RECT 2677.075 814.060 2677.590 814.200 ;
        RECT 2677.270 814.000 2677.590 814.060 ;
        RECT 2677.270 766.260 2677.590 766.320 ;
        RECT 2677.075 766.120 2677.590 766.260 ;
        RECT 2677.270 766.060 2677.590 766.120 ;
        RECT 2677.270 717.640 2677.590 717.700 ;
        RECT 2677.075 717.500 2677.590 717.640 ;
        RECT 2677.270 717.440 2677.590 717.500 ;
        RECT 2677.270 669.700 2677.590 669.760 ;
        RECT 2677.075 669.560 2677.590 669.700 ;
        RECT 2677.270 669.500 2677.590 669.560 ;
        RECT 2677.270 620.740 2677.590 620.800 ;
        RECT 2677.075 620.600 2677.590 620.740 ;
        RECT 2677.270 620.540 2677.590 620.600 ;
        RECT 2677.270 572.800 2677.590 572.860 ;
        RECT 2677.075 572.660 2677.590 572.800 ;
        RECT 2677.270 572.600 2677.590 572.660 ;
        RECT 2677.270 524.180 2677.590 524.240 ;
        RECT 2677.075 524.040 2677.590 524.180 ;
        RECT 2677.270 523.980 2677.590 524.040 ;
        RECT 2677.270 476.240 2677.590 476.300 ;
        RECT 2677.075 476.100 2677.590 476.240 ;
        RECT 2677.270 476.040 2677.590 476.100 ;
        RECT 2677.270 427.620 2677.590 427.680 ;
        RECT 2677.075 427.480 2677.590 427.620 ;
        RECT 2677.270 427.420 2677.590 427.480 ;
        RECT 2677.270 379.680 2677.590 379.740 ;
        RECT 2677.075 379.540 2677.590 379.680 ;
        RECT 2677.270 379.480 2677.590 379.540 ;
        RECT 2677.270 331.060 2677.590 331.120 ;
        RECT 2677.075 330.920 2677.590 331.060 ;
        RECT 2677.270 330.860 2677.590 330.920 ;
        RECT 2677.270 283.120 2677.590 283.180 ;
        RECT 2677.075 282.980 2677.590 283.120 ;
        RECT 2677.270 282.920 2677.590 282.980 ;
        RECT 2677.270 234.500 2677.590 234.560 ;
        RECT 2677.075 234.360 2677.590 234.500 ;
        RECT 2677.270 234.300 2677.590 234.360 ;
        RECT 2677.270 186.560 2677.590 186.620 ;
        RECT 2677.075 186.420 2677.590 186.560 ;
        RECT 2677.270 186.360 2677.590 186.420 ;
        RECT 2677.270 137.940 2677.590 138.000 ;
        RECT 2677.075 137.800 2677.590 137.940 ;
        RECT 2677.270 137.740 2677.590 137.800 ;
        RECT 2677.285 48.520 2677.575 48.565 ;
        RECT 2678.650 48.520 2678.970 48.580 ;
        RECT 2677.285 48.380 2678.970 48.520 ;
        RECT 2677.285 48.335 2677.575 48.380 ;
        RECT 2678.650 48.320 2678.970 48.380 ;
      LAYER via ;
        RECT 1875.520 1472.920 1875.780 1473.180 ;
        RECT 2677.300 1441.980 2677.560 1442.240 ;
        RECT 2677.300 1345.420 2677.560 1345.680 ;
        RECT 2678.220 1345.420 2678.480 1345.680 ;
        RECT 2677.300 1248.860 2677.560 1249.120 ;
        RECT 2678.220 1248.860 2678.480 1249.120 ;
        RECT 2677.300 1152.300 2677.560 1152.560 ;
        RECT 2678.220 1152.300 2678.480 1152.560 ;
        RECT 2677.300 1007.120 2677.560 1007.380 ;
        RECT 2678.220 1007.120 2678.480 1007.380 ;
        RECT 2677.300 910.560 2677.560 910.820 ;
        RECT 2678.220 910.560 2678.480 910.820 ;
        RECT 2677.300 814.000 2677.560 814.260 ;
        RECT 2677.300 766.060 2677.560 766.320 ;
        RECT 2677.300 717.440 2677.560 717.700 ;
        RECT 2677.300 669.500 2677.560 669.760 ;
        RECT 2677.300 620.540 2677.560 620.800 ;
        RECT 2677.300 572.600 2677.560 572.860 ;
        RECT 2677.300 523.980 2677.560 524.240 ;
        RECT 2677.300 476.040 2677.560 476.300 ;
        RECT 2677.300 427.420 2677.560 427.680 ;
        RECT 2677.300 379.480 2677.560 379.740 ;
        RECT 2677.300 330.860 2677.560 331.120 ;
        RECT 2677.300 282.920 2677.560 283.180 ;
        RECT 2677.300 234.300 2677.560 234.560 ;
        RECT 2677.300 186.360 2677.560 186.620 ;
        RECT 2677.300 137.740 2677.560 138.000 ;
        RECT 2678.680 48.320 2678.940 48.580 ;
      LAYER met2 ;
        RECT 1875.970 1700.410 1876.250 1704.000 ;
        RECT 1875.580 1700.270 1876.250 1700.410 ;
        RECT 1875.580 1473.210 1875.720 1700.270 ;
        RECT 1875.970 1700.000 1876.250 1700.270 ;
        RECT 1875.520 1472.890 1875.780 1473.210 ;
        RECT 2677.300 1441.950 2677.560 1442.270 ;
        RECT 2677.360 1393.845 2677.500 1441.950 ;
        RECT 2677.290 1393.475 2677.570 1393.845 ;
        RECT 2678.210 1393.475 2678.490 1393.845 ;
        RECT 2678.280 1345.710 2678.420 1393.475 ;
        RECT 2677.300 1345.390 2677.560 1345.710 ;
        RECT 2678.220 1345.390 2678.480 1345.710 ;
        RECT 2677.360 1297.285 2677.500 1345.390 ;
        RECT 2677.290 1296.915 2677.570 1297.285 ;
        RECT 2678.210 1296.915 2678.490 1297.285 ;
        RECT 2678.280 1249.150 2678.420 1296.915 ;
        RECT 2677.300 1248.830 2677.560 1249.150 ;
        RECT 2678.220 1248.830 2678.480 1249.150 ;
        RECT 2677.360 1200.725 2677.500 1248.830 ;
        RECT 2677.290 1200.355 2677.570 1200.725 ;
        RECT 2678.210 1200.355 2678.490 1200.725 ;
        RECT 2678.280 1152.590 2678.420 1200.355 ;
        RECT 2677.300 1152.270 2677.560 1152.590 ;
        RECT 2678.220 1152.270 2678.480 1152.590 ;
        RECT 2677.360 1104.165 2677.500 1152.270 ;
        RECT 2677.290 1103.795 2677.570 1104.165 ;
        RECT 2678.210 1103.795 2678.490 1104.165 ;
        RECT 2678.280 1055.885 2678.420 1103.795 ;
        RECT 2677.290 1055.515 2677.570 1055.885 ;
        RECT 2678.210 1055.515 2678.490 1055.885 ;
        RECT 2677.360 1007.410 2677.500 1055.515 ;
        RECT 2677.300 1007.090 2677.560 1007.410 ;
        RECT 2678.220 1007.090 2678.480 1007.410 ;
        RECT 2678.280 959.325 2678.420 1007.090 ;
        RECT 2677.290 958.955 2677.570 959.325 ;
        RECT 2678.210 958.955 2678.490 959.325 ;
        RECT 2677.360 910.850 2677.500 958.955 ;
        RECT 2677.300 910.530 2677.560 910.850 ;
        RECT 2678.220 910.530 2678.480 910.850 ;
        RECT 2678.280 862.765 2678.420 910.530 ;
        RECT 2677.290 862.395 2677.570 862.765 ;
        RECT 2678.210 862.395 2678.490 862.765 ;
        RECT 2677.360 814.290 2677.500 862.395 ;
        RECT 2677.300 813.970 2677.560 814.290 ;
        RECT 2677.300 766.030 2677.560 766.350 ;
        RECT 2677.360 717.730 2677.500 766.030 ;
        RECT 2677.300 717.410 2677.560 717.730 ;
        RECT 2677.300 669.470 2677.560 669.790 ;
        RECT 2677.360 620.830 2677.500 669.470 ;
        RECT 2677.300 620.510 2677.560 620.830 ;
        RECT 2677.300 572.570 2677.560 572.890 ;
        RECT 2677.360 524.270 2677.500 572.570 ;
        RECT 2677.300 523.950 2677.560 524.270 ;
        RECT 2677.300 476.010 2677.560 476.330 ;
        RECT 2677.360 427.710 2677.500 476.010 ;
        RECT 2677.300 427.390 2677.560 427.710 ;
        RECT 2677.300 379.450 2677.560 379.770 ;
        RECT 2677.360 331.150 2677.500 379.450 ;
        RECT 2677.300 330.830 2677.560 331.150 ;
        RECT 2677.300 282.890 2677.560 283.210 ;
        RECT 2677.360 234.590 2677.500 282.890 ;
        RECT 2677.300 234.270 2677.560 234.590 ;
        RECT 2677.300 186.330 2677.560 186.650 ;
        RECT 2677.360 138.030 2677.500 186.330 ;
        RECT 2677.300 137.710 2677.560 138.030 ;
        RECT 2678.680 48.290 2678.940 48.610 ;
        RECT 2678.740 2.400 2678.880 48.290 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
      LAYER via2 ;
        RECT 2677.290 1393.520 2677.570 1393.800 ;
        RECT 2678.210 1393.520 2678.490 1393.800 ;
        RECT 2677.290 1296.960 2677.570 1297.240 ;
        RECT 2678.210 1296.960 2678.490 1297.240 ;
        RECT 2677.290 1200.400 2677.570 1200.680 ;
        RECT 2678.210 1200.400 2678.490 1200.680 ;
        RECT 2677.290 1103.840 2677.570 1104.120 ;
        RECT 2678.210 1103.840 2678.490 1104.120 ;
        RECT 2677.290 1055.560 2677.570 1055.840 ;
        RECT 2678.210 1055.560 2678.490 1055.840 ;
        RECT 2677.290 959.000 2677.570 959.280 ;
        RECT 2678.210 959.000 2678.490 959.280 ;
        RECT 2677.290 862.440 2677.570 862.720 ;
        RECT 2678.210 862.440 2678.490 862.720 ;
      LAYER met3 ;
        RECT 2677.265 1393.810 2677.595 1393.825 ;
        RECT 2678.185 1393.810 2678.515 1393.825 ;
        RECT 2677.265 1393.510 2678.515 1393.810 ;
        RECT 2677.265 1393.495 2677.595 1393.510 ;
        RECT 2678.185 1393.495 2678.515 1393.510 ;
        RECT 2677.265 1297.250 2677.595 1297.265 ;
        RECT 2678.185 1297.250 2678.515 1297.265 ;
        RECT 2677.265 1296.950 2678.515 1297.250 ;
        RECT 2677.265 1296.935 2677.595 1296.950 ;
        RECT 2678.185 1296.935 2678.515 1296.950 ;
        RECT 2677.265 1200.690 2677.595 1200.705 ;
        RECT 2678.185 1200.690 2678.515 1200.705 ;
        RECT 2677.265 1200.390 2678.515 1200.690 ;
        RECT 2677.265 1200.375 2677.595 1200.390 ;
        RECT 2678.185 1200.375 2678.515 1200.390 ;
        RECT 2677.265 1104.130 2677.595 1104.145 ;
        RECT 2678.185 1104.130 2678.515 1104.145 ;
        RECT 2677.265 1103.830 2678.515 1104.130 ;
        RECT 2677.265 1103.815 2677.595 1103.830 ;
        RECT 2678.185 1103.815 2678.515 1103.830 ;
        RECT 2677.265 1055.850 2677.595 1055.865 ;
        RECT 2678.185 1055.850 2678.515 1055.865 ;
        RECT 2677.265 1055.550 2678.515 1055.850 ;
        RECT 2677.265 1055.535 2677.595 1055.550 ;
        RECT 2678.185 1055.535 2678.515 1055.550 ;
        RECT 2677.265 959.290 2677.595 959.305 ;
        RECT 2678.185 959.290 2678.515 959.305 ;
        RECT 2677.265 958.990 2678.515 959.290 ;
        RECT 2677.265 958.975 2677.595 958.990 ;
        RECT 2678.185 958.975 2678.515 958.990 ;
        RECT 2677.265 862.730 2677.595 862.745 ;
        RECT 2678.185 862.730 2678.515 862.745 ;
        RECT 2677.265 862.430 2678.515 862.730 ;
        RECT 2677.265 862.415 2677.595 862.430 ;
        RECT 2678.185 862.415 2678.515 862.430 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 0.300 ;
=======
      LAYER li1 ;
        RECT 1939.045 1685.465 1939.215 1690.735 ;
      LAYER mcon ;
        RECT 1939.045 1690.565 1939.215 1690.735 ;
      LAYER met1 ;
        RECT 1879.170 1690.720 1879.490 1690.780 ;
        RECT 1938.985 1690.720 1939.275 1690.765 ;
        RECT 1879.170 1690.580 1939.275 1690.720 ;
        RECT 1879.170 1690.520 1879.490 1690.580 ;
        RECT 1938.985 1690.535 1939.275 1690.580 ;
        RECT 1938.985 1685.620 1939.275 1685.665 ;
        RECT 2073.290 1685.620 2073.610 1685.680 ;
        RECT 1938.985 1685.480 2073.610 1685.620 ;
        RECT 1938.985 1685.435 1939.275 1685.480 ;
        RECT 2073.290 1685.420 2073.610 1685.480 ;
      LAYER via ;
        RECT 1879.200 1690.520 1879.460 1690.780 ;
        RECT 2073.320 1685.420 2073.580 1685.680 ;
      LAYER met2 ;
        RECT 1877.810 1700.410 1878.090 1704.000 ;
        RECT 1877.810 1700.270 1879.400 1700.410 ;
        RECT 1877.810 1700.000 1878.090 1700.270 ;
        RECT 1879.260 1690.810 1879.400 1700.270 ;
        RECT 1879.200 1690.490 1879.460 1690.810 ;
        RECT 2073.320 1685.390 2073.580 1685.710 ;
        RECT 2073.380 20.245 2073.520 1685.390 ;
        RECT 2073.310 19.875 2073.590 20.245 ;
        RECT 2696.610 19.875 2696.890 20.245 ;
        RECT 2696.680 2.400 2696.820 19.875 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
      LAYER via2 ;
        RECT 2073.310 19.920 2073.590 20.200 ;
        RECT 2696.610 19.920 2696.890 20.200 ;
      LAYER met3 ;
        RECT 2073.285 20.210 2073.615 20.225 ;
        RECT 2696.585 20.210 2696.915 20.225 ;
        RECT 2073.285 19.910 2696.915 20.210 ;
        RECT 2073.285 19.895 2073.615 19.910 ;
        RECT 2696.585 19.895 2696.915 19.910 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1881.930 1466.320 1882.250 1466.380 ;
        RECT 2691.070 1466.320 2691.390 1466.380 ;
        RECT 1881.930 1466.180 2691.390 1466.320 ;
        RECT 1881.930 1466.120 1882.250 1466.180 ;
        RECT 2691.070 1466.120 2691.390 1466.180 ;
        RECT 2691.070 62.120 2691.390 62.180 ;
        RECT 2696.590 62.120 2696.910 62.180 ;
        RECT 2691.070 61.980 2696.910 62.120 ;
        RECT 2691.070 61.920 2691.390 61.980 ;
        RECT 2696.590 61.920 2696.910 61.980 ;
      LAYER via ;
        RECT 1881.960 1466.120 1882.220 1466.380 ;
        RECT 2691.100 1466.120 2691.360 1466.380 ;
        RECT 2691.100 61.920 2691.360 62.180 ;
        RECT 2696.620 61.920 2696.880 62.180 ;
      LAYER met2 ;
        RECT 1881.030 1700.410 1881.310 1704.000 ;
        RECT 1881.030 1700.270 1882.160 1700.410 ;
        RECT 1881.030 1700.000 1881.310 1700.270 ;
        RECT 1882.020 1466.410 1882.160 1700.270 ;
        RECT 1881.960 1466.090 1882.220 1466.410 ;
        RECT 2691.100 1466.090 2691.360 1466.410 ;
        RECT 2691.160 62.210 2691.300 1466.090 ;
        RECT 2691.100 61.890 2691.360 62.210 ;
        RECT 2696.620 61.890 2696.880 62.210 ;
        RECT 2696.680 2.400 2696.820 61.890 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 0.300 ;
=======
      LAYER met1 ;
        RECT 1885.610 1684.940 1885.930 1685.000 ;
        RECT 1890.210 1684.940 1890.530 1685.000 ;
        RECT 1885.610 1684.800 1890.530 1684.940 ;
        RECT 1885.610 1684.740 1885.930 1684.800 ;
        RECT 1890.210 1684.740 1890.530 1684.800 ;
        RECT 1890.210 18.940 1890.530 19.000 ;
        RECT 2714.530 18.940 2714.850 19.000 ;
        RECT 1890.210 18.800 2714.850 18.940 ;
        RECT 1890.210 18.740 1890.530 18.800 ;
        RECT 2714.530 18.740 2714.850 18.800 ;
      LAYER via ;
        RECT 1885.640 1684.740 1885.900 1685.000 ;
        RECT 1890.240 1684.740 1890.500 1685.000 ;
        RECT 1890.240 18.740 1890.500 19.000 ;
        RECT 2714.560 18.740 2714.820 19.000 ;
      LAYER met2 ;
        RECT 1885.630 1700.000 1885.910 1704.000 ;
        RECT 1885.700 1685.030 1885.840 1700.000 ;
        RECT 1885.640 1684.710 1885.900 1685.030 ;
        RECT 1890.240 1684.710 1890.500 1685.030 ;
        RECT 1890.300 19.030 1890.440 1684.710 ;
        RECT 1890.240 18.710 1890.500 19.030 ;
        RECT 2714.560 18.710 2714.820 19.030 ;
        RECT 2714.620 2.400 2714.760 18.710 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1883.330 18.560 1883.610 18.840 ;
        RECT 2714.550 18.560 2714.830 18.840 ;
      LAYER met3 ;
        RECT 1883.305 18.850 1883.635 18.865 ;
        RECT 2714.525 18.850 2714.855 18.865 ;
        RECT 1883.305 18.550 2714.855 18.850 ;
        RECT 1883.305 18.535 1883.635 18.550 ;
        RECT 2714.525 18.535 2714.855 18.550 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1890.670 1690.040 1890.990 1690.100 ;
        RECT 1897.110 1690.040 1897.430 1690.100 ;
        RECT 1890.670 1689.900 1897.430 1690.040 ;
        RECT 1890.670 1689.840 1890.990 1689.900 ;
        RECT 1897.110 1689.840 1897.430 1689.900 ;
        RECT 1897.110 18.600 1897.430 18.660 ;
        RECT 2732.470 18.600 2732.790 18.660 ;
        RECT 1897.110 18.460 2732.790 18.600 ;
        RECT 1897.110 18.400 1897.430 18.460 ;
        RECT 2732.470 18.400 2732.790 18.460 ;
      LAYER via ;
        RECT 1890.700 1689.840 1890.960 1690.100 ;
        RECT 1897.140 1689.840 1897.400 1690.100 ;
        RECT 1897.140 18.400 1897.400 18.660 ;
        RECT 2732.500 18.400 2732.760 18.660 ;
      LAYER met2 ;
        RECT 1890.690 1700.000 1890.970 1704.000 ;
        RECT 1890.760 1690.130 1890.900 1700.000 ;
        RECT 1890.700 1689.810 1890.960 1690.130 ;
        RECT 1897.140 1689.810 1897.400 1690.130 ;
        RECT 1897.200 18.690 1897.340 1689.810 ;
        RECT 1897.140 18.370 1897.400 18.690 ;
        RECT 2732.500 18.370 2732.760 18.690 ;
        RECT 2732.560 2.400 2732.700 18.370 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1887.470 1686.600 1887.750 1686.880 ;
        RECT 1897.590 1686.600 1897.870 1686.880 ;
      LAYER met3 ;
        RECT 1887.445 1686.890 1887.775 1686.905 ;
        RECT 1897.565 1686.890 1897.895 1686.905 ;
        RECT 1887.445 1686.590 1897.895 1686.890 ;
        RECT 1887.445 1686.575 1887.775 1686.590 ;
        RECT 1897.565 1686.575 1897.895 1686.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1895.270 1683.920 1895.590 1683.980 ;
        RECT 1896.650 1683.920 1896.970 1683.980 ;
        RECT 1895.270 1683.780 1896.970 1683.920 ;
        RECT 1895.270 1683.720 1895.590 1683.780 ;
        RECT 1896.650 1683.720 1896.970 1683.780 ;
        RECT 1896.650 18.260 1896.970 18.320 ;
        RECT 2750.410 18.260 2750.730 18.320 ;
        RECT 1896.650 18.120 2750.730 18.260 ;
        RECT 1896.650 18.060 1896.970 18.120 ;
        RECT 2750.410 18.060 2750.730 18.120 ;
      LAYER via ;
        RECT 1895.300 1683.720 1895.560 1683.980 ;
        RECT 1896.680 1683.720 1896.940 1683.980 ;
        RECT 1896.680 18.060 1896.940 18.320 ;
        RECT 2750.440 18.060 2750.700 18.320 ;
      LAYER met2 ;
        RECT 1895.290 1700.000 1895.570 1704.000 ;
        RECT 1895.360 1684.010 1895.500 1700.000 ;
        RECT 1895.300 1683.690 1895.560 1684.010 ;
        RECT 1896.680 1683.690 1896.940 1684.010 ;
        RECT 1896.740 18.350 1896.880 1683.690 ;
        RECT 1896.680 18.030 1896.940 18.350 ;
        RECT 2750.440 18.030 2750.700 18.350 ;
        RECT 2750.500 2.400 2750.640 18.030 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1900.330 1684.940 1900.650 1685.000 ;
        RECT 1904.010 1684.940 1904.330 1685.000 ;
        RECT 1900.330 1684.800 1904.330 1684.940 ;
        RECT 1900.330 1684.740 1900.650 1684.800 ;
        RECT 1904.010 1684.740 1904.330 1684.800 ;
        RECT 1904.010 17.920 1904.330 17.980 ;
        RECT 2767.890 17.920 2768.210 17.980 ;
        RECT 1904.010 17.780 2768.210 17.920 ;
        RECT 1904.010 17.720 1904.330 17.780 ;
        RECT 2767.890 17.720 2768.210 17.780 ;
      LAYER via ;
        RECT 1900.360 1684.740 1900.620 1685.000 ;
        RECT 1904.040 1684.740 1904.300 1685.000 ;
        RECT 1904.040 17.720 1904.300 17.980 ;
        RECT 2767.920 17.720 2768.180 17.980 ;
      LAYER met2 ;
        RECT 1900.350 1700.000 1900.630 1704.000 ;
        RECT 1900.420 1685.030 1900.560 1700.000 ;
        RECT 1900.360 1684.710 1900.620 1685.030 ;
        RECT 1904.040 1684.710 1904.300 1685.030 ;
        RECT 1904.100 18.010 1904.240 1684.710 ;
        RECT 1904.040 17.690 1904.300 18.010 ;
        RECT 2767.920 17.690 2768.180 18.010 ;
        RECT 2767.980 2.400 2768.120 17.690 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1373.630 1678.140 1373.950 1678.200 ;
        RECT 1376.390 1678.140 1376.710 1678.200 ;
        RECT 1373.630 1678.000 1376.710 1678.140 ;
        RECT 1373.630 1677.940 1373.950 1678.000 ;
        RECT 1376.390 1677.940 1376.710 1678.000 ;
        RECT 840.950 37.300 841.270 37.360 ;
        RECT 1373.630 37.300 1373.950 37.360 ;
        RECT 840.950 37.160 1373.950 37.300 ;
        RECT 840.950 37.100 841.270 37.160 ;
        RECT 1373.630 37.100 1373.950 37.160 ;
      LAYER via ;
        RECT 1373.660 1677.940 1373.920 1678.200 ;
        RECT 1376.420 1677.940 1376.680 1678.200 ;
        RECT 840.980 37.100 841.240 37.360 ;
        RECT 1373.660 37.100 1373.920 37.360 ;
      LAYER met2 ;
        RECT 1377.790 1700.410 1378.070 1704.000 ;
        RECT 1376.480 1700.270 1378.070 1700.410 ;
        RECT 1376.480 1678.230 1376.620 1700.270 ;
        RECT 1377.790 1700.000 1378.070 1700.270 ;
        RECT 1373.660 1677.910 1373.920 1678.230 ;
        RECT 1376.420 1677.910 1376.680 1678.230 ;
        RECT 1373.720 37.390 1373.860 1677.910 ;
        RECT 840.980 37.070 841.240 37.390 ;
        RECT 1373.660 37.070 1373.920 37.390 ;
        RECT 841.040 2.400 841.180 37.070 ;
        RECT 840.830 -4.800 841.390 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1904.930 1684.260 1905.250 1684.320 ;
        RECT 1910.450 1684.260 1910.770 1684.320 ;
        RECT 1904.930 1684.120 1910.770 1684.260 ;
        RECT 1904.930 1684.060 1905.250 1684.120 ;
        RECT 1910.450 1684.060 1910.770 1684.120 ;
      LAYER via ;
        RECT 1904.960 1684.060 1905.220 1684.320 ;
        RECT 1910.480 1684.060 1910.740 1684.320 ;
      LAYER met2 ;
        RECT 1904.950 1700.000 1905.230 1704.000 ;
        RECT 1905.020 1684.350 1905.160 1700.000 ;
        RECT 1904.960 1684.030 1905.220 1684.350 ;
        RECT 1910.480 1684.030 1910.740 1684.350 ;
        RECT 1910.540 20.245 1910.680 1684.030 ;
        RECT 1910.470 19.875 1910.750 20.245 ;
        RECT 2785.850 19.875 2786.130 20.245 ;
        RECT 2785.920 2.400 2786.060 19.875 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
      LAYER via2 ;
        RECT 1910.470 19.920 1910.750 20.200 ;
        RECT 2785.850 19.920 2786.130 20.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1904.005 18.170 1904.335 18.185 ;
        RECT 2785.825 18.170 2786.155 18.185 ;
        RECT 1904.005 17.870 2786.155 18.170 ;
        RECT 1904.005 17.855 1904.335 17.870 ;
        RECT 2785.825 17.855 2786.155 17.870 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1910.445 20.210 1910.775 20.225 ;
        RECT 2785.825 20.210 2786.155 20.225 ;
        RECT 1910.445 19.910 2786.155 20.210 ;
        RECT 1910.445 19.895 1910.775 19.910 ;
        RECT 2785.825 19.895 2786.155 19.910 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 0.300 ;
=======
      LAYER met1 ;
        RECT 2142.290 19.620 2142.610 19.680 ;
        RECT 2803.770 19.620 2804.090 19.680 ;
        RECT 2142.290 19.480 2804.090 19.620 ;
        RECT 2142.290 19.420 2142.610 19.480 ;
        RECT 2803.770 19.420 2804.090 19.480 ;
      LAYER via ;
        RECT 2142.320 19.420 2142.580 19.680 ;
        RECT 2803.800 19.420 2804.060 19.680 ;
=======
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1910.010 1700.410 1910.290 1704.000 ;
        RECT 1910.010 1700.270 1911.140 1700.410 ;
        RECT 1910.010 1700.000 1910.290 1700.270 ;
        RECT 1911.000 19.565 1911.140 1700.270 ;
        RECT 1910.930 19.195 1911.210 19.565 ;
        RECT 2803.790 19.195 2804.070 19.565 ;
        RECT 2803.860 2.400 2804.000 19.195 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
      LAYER via2 ;
        RECT 1910.930 19.240 1911.210 19.520 ;
        RECT 2803.790 19.240 2804.070 19.520 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1906.765 1688.930 1907.095 1688.945 ;
        RECT 2142.285 1688.930 2142.615 1688.945 ;
        RECT 1906.765 1688.630 2142.615 1688.930 ;
        RECT 1906.765 1688.615 1907.095 1688.630 ;
        RECT 2142.285 1688.615 2142.615 1688.630 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1910.905 19.530 1911.235 19.545 ;
        RECT 2803.765 19.530 2804.095 19.545 ;
        RECT 1910.905 19.230 2804.095 19.530 ;
        RECT 1910.905 19.215 1911.235 19.230 ;
        RECT 2803.765 19.215 2804.095 19.230 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 0.300 ;
=======
      LAYER met1 ;
        RECT 1915.510 1678.140 1915.830 1678.200 ;
        RECT 1917.810 1678.140 1918.130 1678.200 ;
        RECT 1915.510 1678.000 1918.130 1678.140 ;
        RECT 1915.510 1677.940 1915.830 1678.000 ;
        RECT 1917.810 1677.940 1918.130 1678.000 ;
        RECT 1917.350 17.580 1917.670 17.640 ;
        RECT 2821.710 17.580 2822.030 17.640 ;
        RECT 1917.350 17.440 2822.030 17.580 ;
        RECT 1917.350 17.380 1917.670 17.440 ;
        RECT 2821.710 17.380 2822.030 17.440 ;
      LAYER via ;
        RECT 1915.540 1677.940 1915.800 1678.200 ;
        RECT 1917.840 1677.940 1918.100 1678.200 ;
        RECT 1917.380 17.380 1917.640 17.640 ;
        RECT 2821.740 17.380 2822.000 17.640 ;
      LAYER met2 ;
        RECT 1914.610 1700.410 1914.890 1704.000 ;
        RECT 1914.610 1700.270 1915.740 1700.410 ;
        RECT 1914.610 1700.000 1914.890 1700.270 ;
        RECT 1915.600 1678.230 1915.740 1700.270 ;
        RECT 1915.540 1677.910 1915.800 1678.230 ;
        RECT 1917.840 1677.910 1918.100 1678.230 ;
        RECT 1917.900 24.890 1918.040 1677.910 ;
        RECT 1917.440 24.750 1918.040 24.890 ;
        RECT 1917.440 17.670 1917.580 24.750 ;
        RECT 1917.380 17.350 1917.640 17.670 ;
        RECT 2821.740 17.350 2822.000 17.670 ;
        RECT 2821.800 2.400 2821.940 17.350 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1916.910 44.400 1917.190 44.680 ;
        RECT 2821.730 44.400 2822.010 44.680 ;
      LAYER met3 ;
        RECT 1916.885 44.690 1917.215 44.705 ;
        RECT 2821.705 44.690 2822.035 44.705 ;
        RECT 1916.885 44.390 2822.035 44.690 ;
        RECT 1916.885 44.375 1917.215 44.390 ;
        RECT 2821.705 44.375 2822.035 44.390 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 0.300 ;
=======
      LAYER li1 ;
        RECT 2183.765 17.765 2183.935 18.615 ;
      LAYER mcon ;
        RECT 2183.765 18.445 2183.935 18.615 ;
      LAYER met1 ;
        RECT 2183.705 18.600 2183.995 18.645 ;
        RECT 2839.190 18.600 2839.510 18.660 ;
        RECT 2183.705 18.460 2839.510 18.600 ;
        RECT 2183.705 18.415 2183.995 18.460 ;
        RECT 2839.190 18.400 2839.510 18.460 ;
        RECT 2149.190 17.920 2149.510 17.980 ;
        RECT 2183.705 17.920 2183.995 17.965 ;
        RECT 2149.190 17.780 2183.995 17.920 ;
        RECT 2149.190 17.720 2149.510 17.780 ;
        RECT 2183.705 17.735 2183.995 17.780 ;
      LAYER via ;
        RECT 2839.220 18.400 2839.480 18.660 ;
        RECT 2149.220 17.720 2149.480 17.980 ;
      LAYER met2 ;
        RECT 1916.450 1700.000 1916.730 1704.000 ;
        RECT 1916.520 1688.285 1916.660 1700.000 ;
        RECT 1916.450 1687.915 1916.730 1688.285 ;
        RECT 2149.210 1687.915 2149.490 1688.285 ;
        RECT 2149.280 18.010 2149.420 1687.915 ;
        RECT 2839.220 18.370 2839.480 18.690 ;
        RECT 2149.220 17.690 2149.480 18.010 ;
        RECT 2839.280 2.400 2839.420 18.370 ;
=======
      LAYER met1 ;
        RECT 1919.650 1684.260 1919.970 1684.320 ;
        RECT 1924.250 1684.260 1924.570 1684.320 ;
        RECT 1919.650 1684.120 1924.570 1684.260 ;
        RECT 1919.650 1684.060 1919.970 1684.120 ;
        RECT 1924.250 1684.060 1924.570 1684.120 ;
      LAYER via ;
        RECT 1919.680 1684.060 1919.940 1684.320 ;
        RECT 1924.280 1684.060 1924.540 1684.320 ;
      LAYER met2 ;
        RECT 1919.670 1700.000 1919.950 1704.000 ;
        RECT 1919.740 1684.350 1919.880 1700.000 ;
        RECT 1919.680 1684.030 1919.940 1684.350 ;
        RECT 1924.280 1684.030 1924.540 1684.350 ;
        RECT 1924.340 18.885 1924.480 1684.030 ;
        RECT 1924.270 18.515 1924.550 18.885 ;
        RECT 2839.210 18.515 2839.490 18.885 ;
        RECT 2839.280 2.400 2839.420 18.515 ;
>>>>>>> re-updated local openlane
        RECT 2839.070 -4.800 2839.630 2.400 ;
      LAYER via2 ;
        RECT 1924.270 18.560 1924.550 18.840 ;
        RECT 2839.210 18.560 2839.490 18.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1916.425 1688.250 1916.755 1688.265 ;
        RECT 2149.185 1688.250 2149.515 1688.265 ;
        RECT 1916.425 1687.950 2149.515 1688.250 ;
        RECT 1916.425 1687.935 1916.755 1687.950 ;
        RECT 2149.185 1687.935 2149.515 1687.950 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1924.245 18.850 1924.575 18.865 ;
        RECT 2839.185 18.850 2839.515 18.865 ;
        RECT 1924.245 18.550 2839.515 18.850 ;
        RECT 1924.245 18.535 1924.575 18.550 ;
        RECT 2839.185 18.535 2839.515 18.550 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1920.110 1632.240 1920.430 1632.300 ;
        RECT 1924.710 1632.240 1925.030 1632.300 ;
        RECT 1920.110 1632.100 1925.030 1632.240 ;
        RECT 1920.110 1632.040 1920.430 1632.100 ;
        RECT 1924.710 1632.040 1925.030 1632.100 ;
      LAYER via ;
        RECT 1920.140 1632.040 1920.400 1632.300 ;
        RECT 1924.740 1632.040 1925.000 1632.300 ;
=======
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1924.270 1700.410 1924.550 1704.000 ;
        RECT 1924.270 1700.270 1924.940 1700.410 ;
        RECT 1924.270 1700.000 1924.550 1700.270 ;
        RECT 1924.800 18.205 1924.940 1700.270 ;
        RECT 1924.730 17.835 1925.010 18.205 ;
        RECT 2857.150 17.835 2857.430 18.205 ;
        RECT 2857.220 2.400 2857.360 17.835 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
      LAYER via2 ;
        RECT 1924.730 17.880 1925.010 18.160 ;
        RECT 2857.150 17.880 2857.430 18.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1924.705 17.490 1925.035 17.505 ;
        RECT 2857.125 17.490 2857.455 17.505 ;
        RECT 1924.705 17.190 2857.455 17.490 ;
        RECT 1924.705 17.175 1925.035 17.190 ;
        RECT 2857.125 17.175 2857.455 17.190 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1924.705 18.170 1925.035 18.185 ;
        RECT 2857.125 18.170 2857.455 18.185 ;
        RECT 1924.705 17.870 2857.455 18.170 ;
        RECT 1924.705 17.855 1925.035 17.870 ;
        RECT 2857.125 17.855 2857.455 17.870 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 0.300 ;
=======
      LAYER li1 ;
        RECT 2183.305 18.785 2184.395 18.955 ;
        RECT 2183.305 18.445 2183.475 18.785 ;
        RECT 2184.225 17.765 2184.395 18.785 ;
      LAYER met1 ;
        RECT 2180.010 18.600 2180.330 18.660 ;
        RECT 2183.245 18.600 2183.535 18.645 ;
        RECT 2180.010 18.460 2183.535 18.600 ;
        RECT 2180.010 18.400 2180.330 18.460 ;
        RECT 2183.245 18.415 2183.535 18.460 ;
        RECT 2184.165 17.920 2184.455 17.965 ;
        RECT 2875.070 17.920 2875.390 17.980 ;
        RECT 2184.165 17.780 2875.390 17.920 ;
        RECT 2184.165 17.735 2184.455 17.780 ;
        RECT 2875.070 17.720 2875.390 17.780 ;
      LAYER via ;
        RECT 2180.040 18.400 2180.300 18.660 ;
        RECT 2875.100 17.720 2875.360 17.980 ;
      LAYER met2 ;
        RECT 1926.110 1700.000 1926.390 1704.000 ;
        RECT 1926.180 1687.605 1926.320 1700.000 ;
        RECT 1926.110 1687.235 1926.390 1687.605 ;
        RECT 2176.810 1687.235 2177.090 1687.605 ;
        RECT 2176.880 26.250 2177.020 1687.235 ;
        RECT 2176.880 26.110 2180.240 26.250 ;
        RECT 2180.100 18.690 2180.240 26.110 ;
        RECT 2180.040 18.370 2180.300 18.690 ;
        RECT 2875.100 17.690 2875.360 18.010 ;
        RECT 2875.160 2.400 2875.300 17.690 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
      LAYER via2 ;
        RECT 1926.110 1687.280 1926.390 1687.560 ;
        RECT 2176.810 1687.280 2177.090 1687.560 ;
      LAYER met3 ;
        RECT 1926.085 1687.570 1926.415 1687.585 ;
        RECT 2176.785 1687.570 2177.115 1687.585 ;
        RECT 1926.085 1687.270 2177.115 1687.570 ;
        RECT 1926.085 1687.255 1926.415 1687.270 ;
        RECT 2176.785 1687.255 2177.115 1687.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1929.310 1683.920 1929.630 1683.980 ;
        RECT 1931.610 1683.920 1931.930 1683.980 ;
        RECT 1929.310 1683.780 1931.930 1683.920 ;
        RECT 1929.310 1683.720 1929.630 1683.780 ;
        RECT 1931.610 1683.720 1931.930 1683.780 ;
        RECT 1931.610 17.240 1931.930 17.300 ;
        RECT 2875.070 17.240 2875.390 17.300 ;
        RECT 1931.610 17.100 2875.390 17.240 ;
        RECT 1931.610 17.040 1931.930 17.100 ;
        RECT 2875.070 17.040 2875.390 17.100 ;
      LAYER via ;
        RECT 1929.340 1683.720 1929.600 1683.980 ;
        RECT 1931.640 1683.720 1931.900 1683.980 ;
        RECT 1931.640 17.040 1931.900 17.300 ;
        RECT 2875.100 17.040 2875.360 17.300 ;
      LAYER met2 ;
        RECT 1929.330 1700.000 1929.610 1704.000 ;
        RECT 1929.400 1684.010 1929.540 1700.000 ;
        RECT 1929.340 1683.690 1929.600 1684.010 ;
        RECT 1931.640 1683.690 1931.900 1684.010 ;
        RECT 1931.700 17.330 1931.840 1683.690 ;
        RECT 1931.640 17.010 1931.900 17.330 ;
        RECT 2875.100 17.010 2875.360 17.330 ;
        RECT 2875.160 2.400 2875.300 17.010 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1933.910 1685.280 1934.230 1685.340 ;
        RECT 1938.510 1685.280 1938.830 1685.340 ;
        RECT 1933.910 1685.140 1938.830 1685.280 ;
        RECT 1933.910 1685.080 1934.230 1685.140 ;
        RECT 1938.510 1685.080 1938.830 1685.140 ;
      LAYER via ;
        RECT 1933.940 1685.080 1934.200 1685.340 ;
        RECT 1938.540 1685.080 1938.800 1685.340 ;
      LAYER met2 ;
        RECT 1933.930 1700.000 1934.210 1704.000 ;
        RECT 1934.000 1685.370 1934.140 1700.000 ;
        RECT 1933.940 1685.050 1934.200 1685.370 ;
        RECT 1938.540 1685.050 1938.800 1685.370 ;
        RECT 1938.600 17.525 1938.740 1685.050 ;
        RECT 1938.530 17.155 1938.810 17.525 ;
        RECT 2893.030 17.155 2893.310 17.525 ;
        RECT 2893.100 2.400 2893.240 17.155 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 1938.530 17.200 1938.810 17.480 ;
        RECT 2893.030 17.200 2893.310 17.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1931.605 16.810 1931.935 16.825 ;
        RECT 2893.005 16.810 2893.335 16.825 ;
        RECT 1931.605 16.510 2893.335 16.810 ;
        RECT 1931.605 16.495 1931.935 16.510 ;
        RECT 2893.005 16.495 2893.335 16.510 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1938.505 17.490 1938.835 17.505 ;
        RECT 2893.005 17.490 2893.335 17.505 ;
        RECT 1938.505 17.190 2893.335 17.490 ;
        RECT 1938.505 17.175 1938.835 17.190 ;
        RECT 2893.005 17.175 2893.335 17.190 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1938.970 1683.920 1939.290 1683.980 ;
        RECT 1945.410 1683.920 1945.730 1683.980 ;
        RECT 1938.970 1683.780 1945.730 1683.920 ;
        RECT 1938.970 1683.720 1939.290 1683.780 ;
        RECT 1945.410 1683.720 1945.730 1683.780 ;
      LAYER via ;
        RECT 1939.000 1683.720 1939.260 1683.980 ;
        RECT 1945.440 1683.720 1945.700 1683.980 ;
      LAYER met2 ;
        RECT 1938.990 1700.000 1939.270 1704.000 ;
        RECT 1939.060 1684.010 1939.200 1700.000 ;
        RECT 1939.000 1683.690 1939.260 1684.010 ;
        RECT 1945.440 1683.690 1945.700 1684.010 ;
        RECT 1945.500 16.845 1945.640 1683.690 ;
        RECT 1945.430 16.475 1945.710 16.845 ;
        RECT 2910.970 16.475 2911.250 16.845 ;
        RECT 2911.040 2.400 2911.180 16.475 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 1945.430 16.520 1945.710 16.800 ;
        RECT 2910.970 16.520 2911.250 16.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1935.745 1686.890 1936.075 1686.905 ;
        RECT 2218.185 1686.890 2218.515 1686.905 ;
        RECT 1935.745 1686.590 2218.515 1686.890 ;
        RECT 1935.745 1686.575 1936.075 1686.590 ;
        RECT 2218.185 1686.575 2218.515 1686.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1945.405 16.810 1945.735 16.825 ;
        RECT 2910.945 16.810 2911.275 16.825 ;
        RECT 1945.405 16.510 2911.275 16.810 ;
        RECT 1945.405 16.495 1945.735 16.510 ;
        RECT 2910.945 16.495 2911.275 16.510 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 0.300 ;
=======
      LAYER met1 ;
        RECT 858.890 37.300 859.210 37.360 ;
        RECT 1381.910 37.300 1382.230 37.360 ;
        RECT 858.890 37.160 1382.230 37.300 ;
        RECT 858.890 37.100 859.210 37.160 ;
        RECT 1381.910 37.100 1382.230 37.160 ;
      LAYER via ;
        RECT 858.920 37.100 859.180 37.360 ;
        RECT 1381.940 37.100 1382.200 37.360 ;
      LAYER met2 ;
        RECT 1381.470 1700.410 1381.750 1704.000 ;
        RECT 1381.470 1700.270 1382.140 1700.410 ;
        RECT 1381.470 1700.000 1381.750 1700.270 ;
        RECT 1382.000 37.390 1382.140 1700.270 ;
        RECT 858.920 37.070 859.180 37.390 ;
        RECT 1381.940 37.070 1382.200 37.390 ;
        RECT 858.980 2.400 859.120 37.070 ;
        RECT 858.770 -4.800 859.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1381.985 1442.025 1382.155 1490.475 ;
        RECT 1381.985 1297.185 1382.155 1318.095 ;
        RECT 1381.985 1035.045 1382.155 1083.155 ;
        RECT 1381.985 945.285 1382.155 993.395 ;
        RECT 1381.985 655.605 1382.155 703.715 ;
        RECT 1381.985 469.285 1382.155 517.395 ;
        RECT 1382.445 372.725 1382.615 420.835 ;
        RECT 1381.985 241.485 1382.155 289.595 ;
        RECT 1381.985 192.525 1382.155 234.515 ;
      LAYER mcon ;
        RECT 1381.985 1490.305 1382.155 1490.475 ;
        RECT 1381.985 1317.925 1382.155 1318.095 ;
        RECT 1381.985 1082.985 1382.155 1083.155 ;
        RECT 1381.985 993.225 1382.155 993.395 ;
        RECT 1381.985 703.545 1382.155 703.715 ;
        RECT 1381.985 517.225 1382.155 517.395 ;
        RECT 1382.445 420.665 1382.615 420.835 ;
        RECT 1381.985 289.425 1382.155 289.595 ;
        RECT 1381.985 234.345 1382.155 234.515 ;
      LAYER met1 ;
        RECT 1381.910 1490.460 1382.230 1490.520 ;
        RECT 1381.715 1490.320 1382.230 1490.460 ;
        RECT 1381.910 1490.260 1382.230 1490.320 ;
        RECT 1381.925 1442.180 1382.215 1442.225 ;
        RECT 1382.830 1442.180 1383.150 1442.240 ;
        RECT 1381.925 1442.040 1383.150 1442.180 ;
        RECT 1381.925 1441.995 1382.215 1442.040 ;
        RECT 1382.830 1441.980 1383.150 1442.040 ;
        RECT 1382.370 1352.760 1382.690 1352.820 ;
        RECT 1382.830 1352.760 1383.150 1352.820 ;
        RECT 1382.370 1352.620 1383.150 1352.760 ;
        RECT 1382.370 1352.560 1382.690 1352.620 ;
        RECT 1382.830 1352.560 1383.150 1352.620 ;
        RECT 1381.910 1318.080 1382.230 1318.140 ;
        RECT 1381.715 1317.940 1382.230 1318.080 ;
        RECT 1381.910 1317.880 1382.230 1317.940 ;
        RECT 1381.910 1297.340 1382.230 1297.400 ;
        RECT 1381.715 1297.200 1382.230 1297.340 ;
        RECT 1381.910 1297.140 1382.230 1297.200 ;
        RECT 1382.370 1241.920 1382.690 1241.980 ;
        RECT 1383.290 1241.920 1383.610 1241.980 ;
        RECT 1382.370 1241.780 1383.610 1241.920 ;
        RECT 1382.370 1241.720 1382.690 1241.780 ;
        RECT 1383.290 1241.720 1383.610 1241.780 ;
        RECT 1381.910 1090.280 1382.230 1090.340 ;
        RECT 1382.830 1090.280 1383.150 1090.340 ;
        RECT 1381.910 1090.140 1383.150 1090.280 ;
        RECT 1381.910 1090.080 1382.230 1090.140 ;
        RECT 1382.830 1090.080 1383.150 1090.140 ;
        RECT 1381.910 1083.140 1382.230 1083.200 ;
        RECT 1381.715 1083.000 1382.230 1083.140 ;
        RECT 1381.910 1082.940 1382.230 1083.000 ;
        RECT 1381.925 1035.200 1382.215 1035.245 ;
        RECT 1382.370 1035.200 1382.690 1035.260 ;
        RECT 1381.925 1035.060 1382.690 1035.200 ;
        RECT 1381.925 1035.015 1382.215 1035.060 ;
        RECT 1382.370 1035.000 1382.690 1035.060 ;
        RECT 1381.910 993.380 1382.230 993.440 ;
        RECT 1381.715 993.240 1382.230 993.380 ;
        RECT 1381.910 993.180 1382.230 993.240 ;
        RECT 1381.925 945.440 1382.215 945.485 ;
        RECT 1382.370 945.440 1382.690 945.500 ;
        RECT 1381.925 945.300 1382.690 945.440 ;
        RECT 1381.925 945.255 1382.215 945.300 ;
        RECT 1382.370 945.240 1382.690 945.300 ;
        RECT 1381.910 758.920 1382.230 759.180 ;
        RECT 1382.000 758.440 1382.140 758.920 ;
        RECT 1382.370 758.440 1382.690 758.500 ;
        RECT 1382.000 758.300 1382.690 758.440 ;
        RECT 1382.370 758.240 1382.690 758.300 ;
        RECT 1381.910 710.160 1382.230 710.220 ;
        RECT 1383.290 710.160 1383.610 710.220 ;
        RECT 1381.910 710.020 1383.610 710.160 ;
        RECT 1381.910 709.960 1382.230 710.020 ;
        RECT 1383.290 709.960 1383.610 710.020 ;
        RECT 1381.925 703.700 1382.215 703.745 ;
        RECT 1383.290 703.700 1383.610 703.760 ;
        RECT 1381.925 703.560 1383.610 703.700 ;
        RECT 1381.925 703.515 1382.215 703.560 ;
        RECT 1383.290 703.500 1383.610 703.560 ;
        RECT 1381.910 655.760 1382.230 655.820 ;
        RECT 1381.715 655.620 1382.230 655.760 ;
        RECT 1381.910 655.560 1382.230 655.620 ;
        RECT 1381.910 517.380 1382.230 517.440 ;
        RECT 1381.715 517.240 1382.230 517.380 ;
        RECT 1381.910 517.180 1382.230 517.240 ;
        RECT 1381.925 469.440 1382.215 469.485 ;
        RECT 1382.370 469.440 1382.690 469.500 ;
        RECT 1381.925 469.300 1382.690 469.440 ;
        RECT 1381.925 469.255 1382.215 469.300 ;
        RECT 1382.370 469.240 1382.690 469.300 ;
        RECT 1382.370 420.820 1382.690 420.880 ;
        RECT 1382.175 420.680 1382.690 420.820 ;
        RECT 1382.370 420.620 1382.690 420.680 ;
        RECT 1382.370 372.880 1382.690 372.940 ;
        RECT 1382.175 372.740 1382.690 372.880 ;
        RECT 1382.370 372.680 1382.690 372.740 ;
        RECT 1382.370 338.540 1382.690 338.600 ;
        RECT 1382.000 338.400 1382.690 338.540 ;
        RECT 1382.000 337.920 1382.140 338.400 ;
        RECT 1382.370 338.340 1382.690 338.400 ;
        RECT 1381.910 337.660 1382.230 337.920 ;
        RECT 1381.910 289.580 1382.230 289.640 ;
        RECT 1381.715 289.440 1382.230 289.580 ;
        RECT 1381.910 289.380 1382.230 289.440 ;
        RECT 1381.910 241.640 1382.230 241.700 ;
        RECT 1381.715 241.500 1382.230 241.640 ;
        RECT 1381.910 241.440 1382.230 241.500 ;
        RECT 1381.910 234.500 1382.230 234.560 ;
        RECT 1381.715 234.360 1382.230 234.500 ;
        RECT 1381.910 234.300 1382.230 234.360 ;
        RECT 1381.925 192.680 1382.215 192.725 ;
        RECT 1382.830 192.680 1383.150 192.740 ;
        RECT 1381.925 192.540 1383.150 192.680 ;
        RECT 1381.925 192.495 1382.215 192.540 ;
        RECT 1382.830 192.480 1383.150 192.540 ;
        RECT 1381.450 145.080 1381.770 145.140 ;
        RECT 1382.830 145.080 1383.150 145.140 ;
        RECT 1381.450 144.940 1383.150 145.080 ;
        RECT 1381.450 144.880 1381.770 144.940 ;
        RECT 1382.830 144.880 1383.150 144.940 ;
        RECT 1381.450 120.940 1381.770 121.000 ;
        RECT 1382.370 120.940 1382.690 121.000 ;
        RECT 1381.450 120.800 1382.690 120.940 ;
        RECT 1381.450 120.740 1381.770 120.800 ;
        RECT 1382.370 120.740 1382.690 120.800 ;
        RECT 858.890 36.960 859.210 37.020 ;
        RECT 1382.370 36.960 1382.690 37.020 ;
        RECT 858.890 36.820 1382.690 36.960 ;
        RECT 858.890 36.760 859.210 36.820 ;
        RECT 1382.370 36.760 1382.690 36.820 ;
      LAYER via ;
        RECT 1381.940 1490.260 1382.200 1490.520 ;
        RECT 1382.860 1441.980 1383.120 1442.240 ;
        RECT 1382.400 1352.560 1382.660 1352.820 ;
        RECT 1382.860 1352.560 1383.120 1352.820 ;
        RECT 1381.940 1317.880 1382.200 1318.140 ;
        RECT 1381.940 1297.140 1382.200 1297.400 ;
        RECT 1382.400 1241.720 1382.660 1241.980 ;
        RECT 1383.320 1241.720 1383.580 1241.980 ;
        RECT 1381.940 1090.080 1382.200 1090.340 ;
        RECT 1382.860 1090.080 1383.120 1090.340 ;
        RECT 1381.940 1082.940 1382.200 1083.200 ;
        RECT 1382.400 1035.000 1382.660 1035.260 ;
        RECT 1381.940 993.180 1382.200 993.440 ;
        RECT 1382.400 945.240 1382.660 945.500 ;
        RECT 1381.940 758.920 1382.200 759.180 ;
        RECT 1382.400 758.240 1382.660 758.500 ;
        RECT 1381.940 709.960 1382.200 710.220 ;
        RECT 1383.320 709.960 1383.580 710.220 ;
        RECT 1383.320 703.500 1383.580 703.760 ;
        RECT 1381.940 655.560 1382.200 655.820 ;
        RECT 1381.940 517.180 1382.200 517.440 ;
        RECT 1382.400 469.240 1382.660 469.500 ;
        RECT 1382.400 420.620 1382.660 420.880 ;
        RECT 1382.400 372.680 1382.660 372.940 ;
        RECT 1382.400 338.340 1382.660 338.600 ;
        RECT 1381.940 337.660 1382.200 337.920 ;
        RECT 1381.940 289.380 1382.200 289.640 ;
        RECT 1381.940 241.440 1382.200 241.700 ;
        RECT 1381.940 234.300 1382.200 234.560 ;
        RECT 1382.860 192.480 1383.120 192.740 ;
        RECT 1381.480 144.880 1381.740 145.140 ;
        RECT 1382.860 144.880 1383.120 145.140 ;
        RECT 1381.480 120.740 1381.740 121.000 ;
        RECT 1382.400 120.740 1382.660 121.000 ;
        RECT 858.920 36.760 859.180 37.020 ;
        RECT 1382.400 36.760 1382.660 37.020 ;
      LAYER met2 ;
        RECT 1382.390 1700.000 1382.670 1704.000 ;
        RECT 1382.460 1691.570 1382.600 1700.000 ;
        RECT 1382.000 1691.430 1382.600 1691.570 ;
        RECT 1382.000 1690.890 1382.140 1691.430 ;
        RECT 1382.000 1690.750 1382.600 1690.890 ;
        RECT 1382.460 1556.250 1382.600 1690.750 ;
        RECT 1381.540 1556.110 1382.600 1556.250 ;
        RECT 1381.540 1514.770 1381.680 1556.110 ;
        RECT 1381.540 1514.630 1382.140 1514.770 ;
        RECT 1382.000 1490.550 1382.140 1514.630 ;
        RECT 1381.940 1490.230 1382.200 1490.550 ;
        RECT 1382.860 1441.950 1383.120 1442.270 ;
        RECT 1382.920 1352.850 1383.060 1441.950 ;
        RECT 1382.400 1352.530 1382.660 1352.850 ;
        RECT 1382.860 1352.530 1383.120 1352.850 ;
        RECT 1382.460 1345.450 1382.600 1352.530 ;
        RECT 1382.000 1345.310 1382.600 1345.450 ;
        RECT 1382.000 1318.170 1382.140 1345.310 ;
        RECT 1381.940 1317.850 1382.200 1318.170 ;
        RECT 1381.940 1297.110 1382.200 1297.430 ;
        RECT 1382.000 1274.050 1382.140 1297.110 ;
        RECT 1381.540 1273.910 1382.140 1274.050 ;
        RECT 1381.540 1249.005 1381.680 1273.910 ;
        RECT 1381.470 1248.635 1381.750 1249.005 ;
        RECT 1382.390 1248.635 1382.670 1249.005 ;
        RECT 1382.460 1242.010 1382.600 1248.635 ;
        RECT 1382.400 1241.690 1382.660 1242.010 ;
        RECT 1383.320 1241.690 1383.580 1242.010 ;
        RECT 1383.380 1193.925 1383.520 1241.690 ;
        RECT 1382.390 1193.555 1382.670 1193.925 ;
        RECT 1383.310 1193.555 1383.590 1193.925 ;
        RECT 1382.460 1173.410 1382.600 1193.555 ;
        RECT 1382.000 1173.270 1382.600 1173.410 ;
        RECT 1382.000 1146.325 1382.140 1173.270 ;
        RECT 1381.930 1145.955 1382.210 1146.325 ;
        RECT 1382.390 1145.275 1382.670 1145.645 ;
        RECT 1382.460 1097.250 1382.600 1145.275 ;
        RECT 1382.460 1097.110 1383.060 1097.250 ;
        RECT 1382.920 1090.370 1383.060 1097.110 ;
        RECT 1381.940 1090.050 1382.200 1090.370 ;
        RECT 1382.860 1090.050 1383.120 1090.370 ;
        RECT 1382.000 1083.230 1382.140 1090.050 ;
        RECT 1381.940 1082.910 1382.200 1083.230 ;
        RECT 1382.400 1034.970 1382.660 1035.290 ;
        RECT 1382.460 1011.570 1382.600 1034.970 ;
        RECT 1382.000 1011.430 1382.600 1011.570 ;
        RECT 1382.000 993.470 1382.140 1011.430 ;
        RECT 1381.940 993.150 1382.200 993.470 ;
        RECT 1382.400 945.210 1382.660 945.530 ;
        RECT 1382.460 944.930 1382.600 945.210 ;
        RECT 1382.460 944.790 1383.060 944.930 ;
        RECT 1382.920 885.770 1383.060 944.790 ;
        RECT 1382.460 885.630 1383.060 885.770 ;
        RECT 1382.460 831.370 1382.600 885.630 ;
        RECT 1382.000 831.230 1382.600 831.370 ;
        RECT 1382.000 759.210 1382.140 831.230 ;
        RECT 1381.940 758.890 1382.200 759.210 ;
        RECT 1382.400 758.210 1382.660 758.530 ;
        RECT 1382.460 734.810 1382.600 758.210 ;
        RECT 1382.000 734.670 1382.600 734.810 ;
        RECT 1382.000 710.250 1382.140 734.670 ;
        RECT 1381.940 709.930 1382.200 710.250 ;
        RECT 1383.320 709.930 1383.580 710.250 ;
        RECT 1383.380 703.790 1383.520 709.930 ;
        RECT 1383.320 703.470 1383.580 703.790 ;
        RECT 1381.940 655.530 1382.200 655.850 ;
        RECT 1382.000 596.770 1382.140 655.530 ;
        RECT 1382.000 596.630 1382.600 596.770 ;
        RECT 1382.460 532.285 1382.600 596.630 ;
        RECT 1382.390 531.915 1382.670 532.285 ;
        RECT 1381.930 531.235 1382.210 531.605 ;
        RECT 1382.000 517.470 1382.140 531.235 ;
        RECT 1381.940 517.150 1382.200 517.470 ;
        RECT 1382.400 469.210 1382.660 469.530 ;
        RECT 1382.460 420.910 1382.600 469.210 ;
        RECT 1382.400 420.590 1382.660 420.910 ;
        RECT 1382.400 372.650 1382.660 372.970 ;
        RECT 1382.460 338.630 1382.600 372.650 ;
        RECT 1382.400 338.310 1382.660 338.630 ;
        RECT 1381.940 337.630 1382.200 337.950 ;
        RECT 1382.000 289.670 1382.140 337.630 ;
        RECT 1381.940 289.350 1382.200 289.670 ;
        RECT 1381.940 241.410 1382.200 241.730 ;
        RECT 1382.000 234.590 1382.140 241.410 ;
        RECT 1381.940 234.270 1382.200 234.590 ;
        RECT 1382.860 192.450 1383.120 192.770 ;
        RECT 1382.920 145.170 1383.060 192.450 ;
        RECT 1381.480 144.850 1381.740 145.170 ;
        RECT 1382.860 144.850 1383.120 145.170 ;
        RECT 1381.540 121.030 1381.680 144.850 ;
        RECT 1381.480 120.710 1381.740 121.030 ;
        RECT 1382.400 120.710 1382.660 121.030 ;
        RECT 1382.460 37.050 1382.600 120.710 ;
        RECT 858.920 36.730 859.180 37.050 ;
        RECT 1382.400 36.730 1382.660 37.050 ;
        RECT 858.980 2.400 859.120 36.730 ;
        RECT 858.770 -4.800 859.330 2.400 ;
      LAYER via2 ;
        RECT 1381.470 1248.680 1381.750 1248.960 ;
        RECT 1382.390 1248.680 1382.670 1248.960 ;
        RECT 1382.390 1193.600 1382.670 1193.880 ;
        RECT 1383.310 1193.600 1383.590 1193.880 ;
        RECT 1381.930 1146.000 1382.210 1146.280 ;
        RECT 1382.390 1145.320 1382.670 1145.600 ;
        RECT 1382.390 531.960 1382.670 532.240 ;
        RECT 1381.930 531.280 1382.210 531.560 ;
      LAYER met3 ;
        RECT 1381.445 1248.970 1381.775 1248.985 ;
        RECT 1382.365 1248.970 1382.695 1248.985 ;
        RECT 1381.445 1248.670 1382.695 1248.970 ;
        RECT 1381.445 1248.655 1381.775 1248.670 ;
        RECT 1382.365 1248.655 1382.695 1248.670 ;
        RECT 1382.365 1193.890 1382.695 1193.905 ;
        RECT 1383.285 1193.890 1383.615 1193.905 ;
        RECT 1382.365 1193.590 1383.615 1193.890 ;
        RECT 1382.365 1193.575 1382.695 1193.590 ;
        RECT 1383.285 1193.575 1383.615 1193.590 ;
        RECT 1381.905 1146.290 1382.235 1146.305 ;
        RECT 1381.905 1145.975 1382.450 1146.290 ;
        RECT 1382.150 1145.625 1382.450 1145.975 ;
        RECT 1382.150 1145.310 1382.695 1145.625 ;
        RECT 1382.365 1145.295 1382.695 1145.310 ;
        RECT 1382.365 532.250 1382.695 532.265 ;
        RECT 1382.150 531.935 1382.695 532.250 ;
        RECT 1382.150 531.585 1382.450 531.935 ;
        RECT 1381.905 531.270 1382.450 531.585 ;
        RECT 1381.905 531.255 1382.235 531.270 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 0.300 ;
=======
      LAYER li1 ;
        RECT 1383.365 593.045 1383.535 627.895 ;
        RECT 1382.905 469.285 1383.075 496.995 ;
        RECT 1383.365 372.725 1383.535 420.835 ;
        RECT 1382.905 179.605 1383.075 227.715 ;
      LAYER mcon ;
        RECT 1383.365 627.725 1383.535 627.895 ;
        RECT 1382.905 496.825 1383.075 496.995 ;
        RECT 1383.365 420.665 1383.535 420.835 ;
        RECT 1382.905 227.545 1383.075 227.715 ;
      LAYER met1 ;
        RECT 1382.830 1678.480 1383.150 1678.540 ;
        RECT 1386.050 1678.480 1386.370 1678.540 ;
        RECT 1382.830 1678.340 1386.370 1678.480 ;
        RECT 1382.830 1678.280 1383.150 1678.340 ;
        RECT 1386.050 1678.280 1386.370 1678.340 ;
        RECT 1382.830 1607.900 1383.150 1608.160 ;
        RECT 1382.920 1607.420 1383.060 1607.900 ;
        RECT 1383.290 1607.420 1383.610 1607.480 ;
        RECT 1382.920 1607.280 1383.610 1607.420 ;
        RECT 1383.290 1607.220 1383.610 1607.280 ;
        RECT 1383.290 1593.620 1383.610 1593.880 ;
        RECT 1383.380 1593.200 1383.520 1593.620 ;
        RECT 1383.290 1592.940 1383.610 1593.200 ;
        RECT 1383.290 1159.300 1383.610 1159.360 ;
        RECT 1384.210 1159.300 1384.530 1159.360 ;
        RECT 1383.290 1159.160 1384.530 1159.300 ;
        RECT 1383.290 1159.100 1383.610 1159.160 ;
        RECT 1384.210 1159.100 1384.530 1159.160 ;
        RECT 1383.290 966.180 1383.610 966.240 ;
        RECT 1384.210 966.180 1384.530 966.240 ;
        RECT 1383.290 966.040 1384.530 966.180 ;
        RECT 1383.290 965.980 1383.610 966.040 ;
        RECT 1384.210 965.980 1384.530 966.040 ;
        RECT 1383.290 627.880 1383.610 627.940 ;
        RECT 1383.095 627.740 1383.610 627.880 ;
        RECT 1383.290 627.680 1383.610 627.740 ;
        RECT 1383.290 593.200 1383.610 593.260 ;
        RECT 1383.095 593.060 1383.610 593.200 ;
        RECT 1383.290 593.000 1383.610 593.060 ;
        RECT 1382.845 496.980 1383.135 497.025 ;
        RECT 1383.290 496.980 1383.610 497.040 ;
        RECT 1382.845 496.840 1383.610 496.980 ;
        RECT 1382.845 496.795 1383.135 496.840 ;
        RECT 1383.290 496.780 1383.610 496.840 ;
        RECT 1382.830 469.440 1383.150 469.500 ;
        RECT 1382.635 469.300 1383.150 469.440 ;
        RECT 1382.830 469.240 1383.150 469.300 ;
        RECT 1382.830 427.960 1383.150 428.020 ;
        RECT 1383.290 427.960 1383.610 428.020 ;
        RECT 1382.830 427.820 1383.610 427.960 ;
        RECT 1382.830 427.760 1383.150 427.820 ;
        RECT 1383.290 427.760 1383.610 427.820 ;
        RECT 1383.290 420.820 1383.610 420.880 ;
        RECT 1383.095 420.680 1383.610 420.820 ;
        RECT 1383.290 420.620 1383.610 420.680 ;
        RECT 1383.290 372.880 1383.610 372.940 ;
        RECT 1383.095 372.740 1383.610 372.880 ;
        RECT 1383.290 372.680 1383.610 372.740 ;
        RECT 1382.845 227.700 1383.135 227.745 ;
        RECT 1383.750 227.700 1384.070 227.760 ;
        RECT 1382.845 227.560 1384.070 227.700 ;
        RECT 1382.845 227.515 1383.135 227.560 ;
        RECT 1383.750 227.500 1384.070 227.560 ;
        RECT 1382.830 179.760 1383.150 179.820 ;
        RECT 1382.635 179.620 1383.150 179.760 ;
        RECT 1382.830 179.560 1383.150 179.620 ;
        RECT 876.830 36.960 877.150 37.020 ;
        RECT 1383.290 36.960 1383.610 37.020 ;
        RECT 876.830 36.820 1383.610 36.960 ;
        RECT 876.830 36.760 877.150 36.820 ;
        RECT 1383.290 36.760 1383.610 36.820 ;
      LAYER via ;
        RECT 1382.860 1678.280 1383.120 1678.540 ;
        RECT 1386.080 1678.280 1386.340 1678.540 ;
        RECT 1382.860 1607.900 1383.120 1608.160 ;
        RECT 1383.320 1607.220 1383.580 1607.480 ;
        RECT 1383.320 1593.620 1383.580 1593.880 ;
        RECT 1383.320 1592.940 1383.580 1593.200 ;
        RECT 1383.320 1159.100 1383.580 1159.360 ;
        RECT 1384.240 1159.100 1384.500 1159.360 ;
        RECT 1383.320 965.980 1383.580 966.240 ;
        RECT 1384.240 965.980 1384.500 966.240 ;
        RECT 1383.320 627.680 1383.580 627.940 ;
        RECT 1383.320 593.000 1383.580 593.260 ;
        RECT 1383.320 496.780 1383.580 497.040 ;
        RECT 1382.860 469.240 1383.120 469.500 ;
        RECT 1382.860 427.760 1383.120 428.020 ;
        RECT 1383.320 427.760 1383.580 428.020 ;
        RECT 1383.320 420.620 1383.580 420.880 ;
        RECT 1383.320 372.680 1383.580 372.940 ;
        RECT 1383.780 227.500 1384.040 227.760 ;
        RECT 1382.860 179.560 1383.120 179.820 ;
        RECT 876.860 36.760 877.120 37.020 ;
        RECT 1383.320 36.760 1383.580 37.020 ;
      LAYER met2 ;
        RECT 1386.530 1700.410 1386.810 1704.000 ;
        RECT 1386.140 1700.270 1386.810 1700.410 ;
        RECT 1386.140 1678.570 1386.280 1700.270 ;
        RECT 1386.530 1700.000 1386.810 1700.270 ;
        RECT 1382.860 1678.250 1383.120 1678.570 ;
        RECT 1386.080 1678.250 1386.340 1678.570 ;
        RECT 1382.920 1608.190 1383.060 1678.250 ;
        RECT 1382.860 1607.870 1383.120 1608.190 ;
        RECT 1383.320 1607.190 1383.580 1607.510 ;
        RECT 1383.380 1593.910 1383.520 1607.190 ;
        RECT 1383.320 1593.590 1383.580 1593.910 ;
        RECT 1383.320 1592.910 1383.580 1593.230 ;
        RECT 1383.380 1463.090 1383.520 1592.910 ;
        RECT 1382.920 1462.950 1383.520 1463.090 ;
        RECT 1382.920 1462.410 1383.060 1462.950 ;
        RECT 1382.920 1462.270 1383.520 1462.410 ;
        RECT 1383.380 1366.530 1383.520 1462.270 ;
        RECT 1382.920 1366.390 1383.520 1366.530 ;
        RECT 1382.920 1365.850 1383.060 1366.390 ;
        RECT 1382.920 1365.710 1383.520 1365.850 ;
        RECT 1383.380 1269.970 1383.520 1365.710 ;
        RECT 1382.920 1269.830 1383.520 1269.970 ;
        RECT 1382.920 1269.290 1383.060 1269.830 ;
        RECT 1382.920 1269.150 1383.520 1269.290 ;
        RECT 1383.380 1207.525 1383.520 1269.150 ;
        RECT 1383.310 1207.155 1383.590 1207.525 ;
        RECT 1384.230 1207.155 1384.510 1207.525 ;
        RECT 1384.300 1159.390 1384.440 1207.155 ;
        RECT 1383.320 1159.070 1383.580 1159.390 ;
        RECT 1384.240 1159.070 1384.500 1159.390 ;
        RECT 1383.380 1014.405 1383.520 1159.070 ;
        RECT 1383.310 1014.035 1383.590 1014.405 ;
        RECT 1384.230 1014.035 1384.510 1014.405 ;
        RECT 1384.300 966.270 1384.440 1014.035 ;
        RECT 1383.320 965.950 1383.580 966.270 ;
        RECT 1384.240 965.950 1384.500 966.270 ;
        RECT 1383.380 883.730 1383.520 965.950 ;
        RECT 1382.920 883.590 1383.520 883.730 ;
        RECT 1382.920 883.050 1383.060 883.590 ;
        RECT 1382.920 882.910 1383.520 883.050 ;
        RECT 1383.380 787.170 1383.520 882.910 ;
        RECT 1382.920 787.030 1383.520 787.170 ;
        RECT 1382.920 785.810 1383.060 787.030 ;
        RECT 1382.920 785.670 1383.520 785.810 ;
        RECT 1383.380 627.970 1383.520 785.670 ;
        RECT 1383.320 627.650 1383.580 627.970 ;
        RECT 1383.320 592.970 1383.580 593.290 ;
        RECT 1383.380 497.070 1383.520 592.970 ;
        RECT 1383.320 496.750 1383.580 497.070 ;
        RECT 1382.860 469.210 1383.120 469.530 ;
        RECT 1382.920 428.050 1383.060 469.210 ;
        RECT 1382.860 427.730 1383.120 428.050 ;
        RECT 1383.320 427.730 1383.580 428.050 ;
        RECT 1383.380 420.910 1383.520 427.730 ;
        RECT 1383.320 420.590 1383.580 420.910 ;
        RECT 1383.320 372.650 1383.580 372.970 ;
        RECT 1383.380 235.125 1383.520 372.650 ;
        RECT 1383.310 234.755 1383.590 235.125 ;
        RECT 1383.770 234.075 1384.050 234.445 ;
        RECT 1383.840 227.790 1383.980 234.075 ;
        RECT 1383.780 227.470 1384.040 227.790 ;
        RECT 1382.860 179.530 1383.120 179.850 ;
        RECT 1382.920 144.570 1383.060 179.530 ;
        RECT 1382.920 144.430 1383.520 144.570 ;
        RECT 1383.380 37.050 1383.520 144.430 ;
        RECT 876.860 36.730 877.120 37.050 ;
        RECT 1383.320 36.730 1383.580 37.050 ;
        RECT 876.920 2.400 877.060 36.730 ;
        RECT 876.710 -4.800 877.270 2.400 ;
      LAYER via2 ;
        RECT 1383.310 1207.200 1383.590 1207.480 ;
        RECT 1384.230 1207.200 1384.510 1207.480 ;
        RECT 1383.310 1014.080 1383.590 1014.360 ;
        RECT 1384.230 1014.080 1384.510 1014.360 ;
        RECT 1383.310 234.800 1383.590 235.080 ;
        RECT 1383.770 234.120 1384.050 234.400 ;
      LAYER met3 ;
        RECT 1383.285 1207.490 1383.615 1207.505 ;
        RECT 1384.205 1207.490 1384.535 1207.505 ;
        RECT 1383.285 1207.190 1384.535 1207.490 ;
        RECT 1383.285 1207.175 1383.615 1207.190 ;
        RECT 1384.205 1207.175 1384.535 1207.190 ;
        RECT 1383.285 1014.370 1383.615 1014.385 ;
        RECT 1384.205 1014.370 1384.535 1014.385 ;
        RECT 1383.285 1014.070 1384.535 1014.370 ;
        RECT 1383.285 1014.055 1383.615 1014.070 ;
        RECT 1384.205 1014.055 1384.535 1014.070 ;
        RECT 1383.285 235.090 1383.615 235.105 ;
        RECT 1383.070 234.775 1383.615 235.090 ;
        RECT 1383.070 234.410 1383.370 234.775 ;
        RECT 1383.745 234.410 1384.075 234.425 ;
        RECT 1383.070 234.110 1384.075 234.410 ;
        RECT 1383.745 234.095 1384.075 234.110 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1387.430 759.260 1387.750 759.520 ;
        RECT 1387.520 758.840 1387.660 759.260 ;
        RECT 1387.430 758.580 1387.750 758.840 ;
        RECT 876.830 36.620 877.150 36.680 ;
        RECT 1387.430 36.620 1387.750 36.680 ;
        RECT 876.830 36.480 1387.750 36.620 ;
        RECT 876.830 36.420 877.150 36.480 ;
        RECT 1387.430 36.420 1387.750 36.480 ;
      LAYER via ;
        RECT 1387.460 759.260 1387.720 759.520 ;
        RECT 1387.460 758.580 1387.720 758.840 ;
        RECT 876.860 36.420 877.120 36.680 ;
        RECT 1387.460 36.420 1387.720 36.680 ;
      LAYER met2 ;
        RECT 1387.450 1700.000 1387.730 1704.000 ;
        RECT 1387.520 759.550 1387.660 1700.000 ;
        RECT 1387.460 759.230 1387.720 759.550 ;
        RECT 1387.460 758.550 1387.720 758.870 ;
        RECT 1387.520 36.710 1387.660 758.550 ;
        RECT 876.860 36.390 877.120 36.710 ;
        RECT 1387.460 36.390 1387.720 36.710 ;
        RECT 876.920 2.400 877.060 36.390 ;
        RECT 876.710 -4.800 877.270 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 0.300 ;
=======
      LAYER met1 ;
        RECT 1387.890 1678.140 1388.210 1678.200 ;
        RECT 1391.110 1678.140 1391.430 1678.200 ;
        RECT 1387.890 1678.000 1391.430 1678.140 ;
        RECT 1387.890 1677.940 1388.210 1678.000 ;
        RECT 1391.110 1677.940 1391.430 1678.000 ;
        RECT 1387.890 759.260 1388.210 759.520 ;
        RECT 1387.980 758.840 1388.120 759.260 ;
        RECT 1387.890 758.580 1388.210 758.840 ;
        RECT 1387.890 620.540 1388.210 620.800 ;
        RECT 1387.980 620.120 1388.120 620.540 ;
        RECT 1387.890 619.860 1388.210 620.120 ;
        RECT 894.770 36.280 895.090 36.340 ;
        RECT 1387.890 36.280 1388.210 36.340 ;
        RECT 894.770 36.140 1388.210 36.280 ;
        RECT 894.770 36.080 895.090 36.140 ;
        RECT 1387.890 36.080 1388.210 36.140 ;
      LAYER via ;
        RECT 1387.920 1677.940 1388.180 1678.200 ;
        RECT 1391.140 1677.940 1391.400 1678.200 ;
        RECT 1387.920 759.260 1388.180 759.520 ;
        RECT 1387.920 758.580 1388.180 758.840 ;
        RECT 1387.920 620.540 1388.180 620.800 ;
        RECT 1387.920 619.860 1388.180 620.120 ;
        RECT 894.800 36.080 895.060 36.340 ;
        RECT 1387.920 36.080 1388.180 36.340 ;
      LAYER met2 ;
        RECT 1392.050 1700.410 1392.330 1704.000 ;
        RECT 1391.200 1700.270 1392.330 1700.410 ;
        RECT 1391.200 1678.230 1391.340 1700.270 ;
        RECT 1392.050 1700.000 1392.330 1700.270 ;
        RECT 1387.920 1677.910 1388.180 1678.230 ;
        RECT 1391.140 1677.910 1391.400 1678.230 ;
        RECT 1387.980 759.550 1388.120 1677.910 ;
        RECT 1387.920 759.230 1388.180 759.550 ;
        RECT 1387.920 758.550 1388.180 758.870 ;
        RECT 1387.980 620.830 1388.120 758.550 ;
        RECT 1387.920 620.510 1388.180 620.830 ;
        RECT 1387.920 619.830 1388.180 620.150 ;
        RECT 1387.980 36.370 1388.120 619.830 ;
        RECT 894.800 36.050 895.060 36.370 ;
        RECT 1387.920 36.050 1388.180 36.370 ;
        RECT 894.860 2.400 895.000 36.050 ;
        RECT 894.650 -4.800 895.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 0.300 ;
=======
      LAYER met1 ;
        RECT 912.710 35.940 913.030 36.000 ;
        RECT 1394.790 35.940 1395.110 36.000 ;
        RECT 912.710 35.800 1395.110 35.940 ;
        RECT 912.710 35.740 913.030 35.800 ;
        RECT 1394.790 35.740 1395.110 35.800 ;
      LAYER via ;
        RECT 912.740 35.740 913.000 36.000 ;
        RECT 1394.820 35.740 1395.080 36.000 ;
      LAYER met2 ;
        RECT 1397.110 1700.410 1397.390 1704.000 ;
        RECT 1395.800 1700.270 1397.390 1700.410 ;
        RECT 1395.800 1678.140 1395.940 1700.270 ;
        RECT 1397.110 1700.000 1397.390 1700.270 ;
        RECT 1394.880 1678.000 1395.940 1678.140 ;
        RECT 1394.880 36.030 1395.020 1678.000 ;
        RECT 912.740 35.710 913.000 36.030 ;
        RECT 1394.820 35.710 1395.080 36.030 ;
        RECT 912.800 2.400 912.940 35.710 ;
        RECT 912.590 -4.800 913.150 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 0.300 ;
=======
      LAYER met1 ;
        RECT 930.190 35.940 930.510 36.000 ;
        RECT 1401.690 35.940 1402.010 36.000 ;
        RECT 930.190 35.800 1402.010 35.940 ;
        RECT 930.190 35.740 930.510 35.800 ;
        RECT 1401.690 35.740 1402.010 35.800 ;
      LAYER via ;
        RECT 930.220 35.740 930.480 36.000 ;
        RECT 1401.720 35.740 1401.980 36.000 ;
      LAYER met2 ;
        RECT 1400.790 1700.410 1401.070 1704.000 ;
        RECT 1400.790 1700.270 1401.920 1700.410 ;
        RECT 1400.790 1700.000 1401.070 1700.270 ;
        RECT 1401.780 36.030 1401.920 1700.270 ;
        RECT 930.220 35.710 930.480 36.030 ;
        RECT 1401.720 35.710 1401.980 36.030 ;
        RECT 930.280 2.400 930.420 35.710 ;
        RECT 930.070 -4.800 930.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1402.225 1538.925 1402.395 1563.235 ;
        RECT 1402.685 1349.545 1402.855 1400.715 ;
        RECT 1402.225 1321.325 1402.395 1338.835 ;
        RECT 1401.765 1090.125 1401.935 1104.575 ;
        RECT 1401.765 758.965 1401.935 807.075 ;
        RECT 1402.685 620.925 1402.855 669.375 ;
        RECT 1401.765 469.285 1401.935 516.715 ;
        RECT 1402.685 347.565 1402.855 386.155 ;
        RECT 1401.765 282.965 1401.935 331.075 ;
        RECT 1402.685 186.405 1402.855 258.995 ;
        RECT 1401.765 89.845 1401.935 137.955 ;
      LAYER mcon ;
        RECT 1402.225 1563.065 1402.395 1563.235 ;
        RECT 1402.685 1400.545 1402.855 1400.715 ;
        RECT 1402.225 1338.665 1402.395 1338.835 ;
        RECT 1401.765 1104.405 1401.935 1104.575 ;
        RECT 1401.765 806.905 1401.935 807.075 ;
        RECT 1402.685 669.205 1402.855 669.375 ;
        RECT 1401.765 516.545 1401.935 516.715 ;
        RECT 1402.685 385.985 1402.855 386.155 ;
        RECT 1401.765 330.905 1401.935 331.075 ;
        RECT 1402.685 258.825 1402.855 258.995 ;
        RECT 1401.765 137.785 1401.935 137.955 ;
      LAYER met1 ;
        RECT 1402.165 1563.220 1402.455 1563.265 ;
        RECT 1402.610 1563.220 1402.930 1563.280 ;
        RECT 1402.165 1563.080 1402.930 1563.220 ;
        RECT 1402.165 1563.035 1402.455 1563.080 ;
        RECT 1402.610 1563.020 1402.930 1563.080 ;
        RECT 1402.150 1539.080 1402.470 1539.140 ;
        RECT 1401.955 1538.940 1402.470 1539.080 ;
        RECT 1402.150 1538.880 1402.470 1538.940 ;
        RECT 1402.150 1448.980 1402.470 1449.040 ;
        RECT 1402.610 1448.980 1402.930 1449.040 ;
        RECT 1402.150 1448.840 1402.930 1448.980 ;
        RECT 1402.150 1448.780 1402.470 1448.840 ;
        RECT 1402.610 1448.780 1402.930 1448.840 ;
        RECT 1402.610 1400.700 1402.930 1400.760 ;
        RECT 1402.415 1400.560 1402.930 1400.700 ;
        RECT 1402.610 1400.500 1402.930 1400.560 ;
        RECT 1402.150 1349.700 1402.470 1349.760 ;
        RECT 1402.625 1349.700 1402.915 1349.745 ;
        RECT 1402.150 1349.560 1402.915 1349.700 ;
        RECT 1402.150 1349.500 1402.470 1349.560 ;
        RECT 1402.625 1349.515 1402.915 1349.560 ;
        RECT 1402.150 1338.820 1402.470 1338.880 ;
        RECT 1401.955 1338.680 1402.470 1338.820 ;
        RECT 1402.150 1338.620 1402.470 1338.680 ;
        RECT 1402.165 1321.480 1402.455 1321.525 ;
        RECT 1402.610 1321.480 1402.930 1321.540 ;
        RECT 1402.165 1321.340 1402.930 1321.480 ;
        RECT 1402.165 1321.295 1402.455 1321.340 ;
        RECT 1402.610 1321.280 1402.930 1321.340 ;
        RECT 1401.690 1152.500 1402.010 1152.560 ;
        RECT 1402.610 1152.500 1402.930 1152.560 ;
        RECT 1401.690 1152.360 1402.930 1152.500 ;
        RECT 1401.690 1152.300 1402.010 1152.360 ;
        RECT 1402.610 1152.300 1402.930 1152.360 ;
        RECT 1401.705 1104.560 1401.995 1104.605 ;
        RECT 1402.610 1104.560 1402.930 1104.620 ;
        RECT 1401.705 1104.420 1402.930 1104.560 ;
        RECT 1401.705 1104.375 1401.995 1104.420 ;
        RECT 1402.610 1104.360 1402.930 1104.420 ;
        RECT 1401.690 1090.280 1402.010 1090.340 ;
        RECT 1401.495 1090.140 1402.010 1090.280 ;
        RECT 1401.690 1090.080 1402.010 1090.140 ;
        RECT 1401.690 1028.200 1402.010 1028.460 ;
        RECT 1401.780 1027.720 1401.920 1028.200 ;
        RECT 1402.150 1027.720 1402.470 1027.780 ;
        RECT 1401.780 1027.580 1402.470 1027.720 ;
        RECT 1402.150 1027.520 1402.470 1027.580 ;
        RECT 1402.150 980.120 1402.470 980.180 ;
        RECT 1401.780 979.980 1402.470 980.120 ;
        RECT 1401.780 979.840 1401.920 979.980 ;
        RECT 1402.150 979.920 1402.470 979.980 ;
        RECT 1401.690 979.580 1402.010 979.840 ;
        RECT 1401.690 903.960 1402.010 904.020 ;
        RECT 1402.610 903.960 1402.930 904.020 ;
        RECT 1401.690 903.820 1402.930 903.960 ;
        RECT 1401.690 903.760 1402.010 903.820 ;
        RECT 1402.610 903.760 1402.930 903.820 ;
        RECT 1401.705 807.060 1401.995 807.105 ;
        RECT 1402.610 807.060 1402.930 807.120 ;
        RECT 1401.705 806.920 1402.930 807.060 ;
        RECT 1401.705 806.875 1401.995 806.920 ;
        RECT 1402.610 806.860 1402.930 806.920 ;
        RECT 1401.690 759.120 1402.010 759.180 ;
        RECT 1401.495 758.980 1402.010 759.120 ;
        RECT 1401.690 758.920 1402.010 758.980 ;
        RECT 1402.610 669.360 1402.930 669.420 ;
        RECT 1402.415 669.220 1402.930 669.360 ;
        RECT 1402.610 669.160 1402.930 669.220 ;
        RECT 1402.610 621.080 1402.930 621.140 ;
        RECT 1402.415 620.940 1402.930 621.080 ;
        RECT 1402.610 620.880 1402.930 620.940 ;
        RECT 1401.690 517.180 1402.010 517.440 ;
        RECT 1401.780 516.745 1401.920 517.180 ;
        RECT 1401.705 516.515 1401.995 516.745 ;
        RECT 1401.690 469.440 1402.010 469.500 ;
        RECT 1401.495 469.300 1402.010 469.440 ;
        RECT 1401.690 469.240 1402.010 469.300 ;
        RECT 1401.690 427.960 1402.010 428.020 ;
        RECT 1402.610 427.960 1402.930 428.020 ;
        RECT 1401.690 427.820 1402.930 427.960 ;
        RECT 1401.690 427.760 1402.010 427.820 ;
        RECT 1402.610 427.760 1402.930 427.820 ;
        RECT 1402.610 386.140 1402.930 386.200 ;
        RECT 1402.415 386.000 1402.930 386.140 ;
        RECT 1402.610 385.940 1402.930 386.000 ;
        RECT 1401.690 347.720 1402.010 347.780 ;
        RECT 1402.625 347.720 1402.915 347.765 ;
        RECT 1401.690 347.580 1402.915 347.720 ;
        RECT 1401.690 347.520 1402.010 347.580 ;
        RECT 1402.625 347.535 1402.915 347.580 ;
        RECT 1401.690 331.060 1402.010 331.120 ;
        RECT 1401.495 330.920 1402.010 331.060 ;
        RECT 1401.690 330.860 1402.010 330.920 ;
        RECT 1401.690 283.120 1402.010 283.180 ;
        RECT 1401.495 282.980 1402.010 283.120 ;
        RECT 1401.690 282.920 1402.010 282.980 ;
        RECT 1401.690 258.980 1402.010 259.040 ;
        RECT 1402.625 258.980 1402.915 259.025 ;
        RECT 1401.690 258.840 1402.915 258.980 ;
        RECT 1401.690 258.780 1402.010 258.840 ;
        RECT 1402.625 258.795 1402.915 258.840 ;
        RECT 1402.610 186.560 1402.930 186.620 ;
        RECT 1402.415 186.420 1402.930 186.560 ;
        RECT 1402.610 186.360 1402.930 186.420 ;
        RECT 1401.705 137.940 1401.995 137.985 ;
        RECT 1402.610 137.940 1402.930 138.000 ;
        RECT 1401.705 137.800 1402.930 137.940 ;
        RECT 1401.705 137.755 1401.995 137.800 ;
        RECT 1402.610 137.740 1402.930 137.800 ;
        RECT 1401.690 90.000 1402.010 90.060 ;
        RECT 1401.495 89.860 1402.010 90.000 ;
        RECT 1401.690 89.800 1402.010 89.860 ;
        RECT 930.190 35.600 930.510 35.660 ;
        RECT 1401.690 35.600 1402.010 35.660 ;
        RECT 930.190 35.460 1402.010 35.600 ;
        RECT 930.190 35.400 930.510 35.460 ;
        RECT 1401.690 35.400 1402.010 35.460 ;
      LAYER via ;
        RECT 1402.640 1563.020 1402.900 1563.280 ;
        RECT 1402.180 1538.880 1402.440 1539.140 ;
        RECT 1402.180 1448.780 1402.440 1449.040 ;
        RECT 1402.640 1448.780 1402.900 1449.040 ;
        RECT 1402.640 1400.500 1402.900 1400.760 ;
        RECT 1402.180 1349.500 1402.440 1349.760 ;
        RECT 1402.180 1338.620 1402.440 1338.880 ;
        RECT 1402.640 1321.280 1402.900 1321.540 ;
        RECT 1401.720 1152.300 1401.980 1152.560 ;
        RECT 1402.640 1152.300 1402.900 1152.560 ;
        RECT 1402.640 1104.360 1402.900 1104.620 ;
        RECT 1401.720 1090.080 1401.980 1090.340 ;
        RECT 1401.720 1028.200 1401.980 1028.460 ;
        RECT 1402.180 1027.520 1402.440 1027.780 ;
        RECT 1402.180 979.920 1402.440 980.180 ;
        RECT 1401.720 979.580 1401.980 979.840 ;
        RECT 1401.720 903.760 1401.980 904.020 ;
        RECT 1402.640 903.760 1402.900 904.020 ;
        RECT 1402.640 806.860 1402.900 807.120 ;
        RECT 1401.720 758.920 1401.980 759.180 ;
        RECT 1402.640 669.160 1402.900 669.420 ;
        RECT 1402.640 620.880 1402.900 621.140 ;
        RECT 1401.720 517.180 1401.980 517.440 ;
        RECT 1401.720 469.240 1401.980 469.500 ;
        RECT 1401.720 427.760 1401.980 428.020 ;
        RECT 1402.640 427.760 1402.900 428.020 ;
        RECT 1402.640 385.940 1402.900 386.200 ;
        RECT 1401.720 347.520 1401.980 347.780 ;
        RECT 1401.720 330.860 1401.980 331.120 ;
        RECT 1401.720 282.920 1401.980 283.180 ;
        RECT 1401.720 258.780 1401.980 259.040 ;
        RECT 1402.640 186.360 1402.900 186.620 ;
        RECT 1402.640 137.740 1402.900 138.000 ;
        RECT 1401.720 89.800 1401.980 90.060 ;
        RECT 930.220 35.400 930.480 35.660 ;
        RECT 1401.720 35.400 1401.980 35.660 ;
      LAYER met2 ;
        RECT 1401.710 1700.410 1401.990 1704.000 ;
        RECT 1401.710 1700.270 1402.840 1700.410 ;
        RECT 1401.710 1700.000 1401.990 1700.270 ;
        RECT 1402.700 1563.310 1402.840 1700.270 ;
        RECT 1402.640 1562.990 1402.900 1563.310 ;
        RECT 1402.180 1538.850 1402.440 1539.170 ;
        RECT 1402.240 1449.070 1402.380 1538.850 ;
        RECT 1402.180 1448.750 1402.440 1449.070 ;
        RECT 1402.640 1448.750 1402.900 1449.070 ;
        RECT 1402.700 1400.790 1402.840 1448.750 ;
        RECT 1402.640 1400.470 1402.900 1400.790 ;
        RECT 1402.180 1349.470 1402.440 1349.790 ;
        RECT 1402.240 1338.910 1402.380 1349.470 ;
        RECT 1402.180 1338.590 1402.440 1338.910 ;
        RECT 1402.640 1321.250 1402.900 1321.570 ;
        RECT 1402.700 1152.590 1402.840 1321.250 ;
        RECT 1401.720 1152.445 1401.980 1152.590 ;
        RECT 1402.640 1152.445 1402.900 1152.590 ;
        RECT 1401.710 1152.075 1401.990 1152.445 ;
        RECT 1402.630 1152.075 1402.910 1152.445 ;
        RECT 1402.700 1104.650 1402.840 1152.075 ;
        RECT 1402.640 1104.330 1402.900 1104.650 ;
        RECT 1401.720 1090.050 1401.980 1090.370 ;
        RECT 1401.780 1028.490 1401.920 1090.050 ;
        RECT 1401.720 1028.170 1401.980 1028.490 ;
        RECT 1402.180 1027.490 1402.440 1027.810 ;
        RECT 1402.240 980.210 1402.380 1027.490 ;
        RECT 1402.180 979.890 1402.440 980.210 ;
        RECT 1401.720 979.550 1401.980 979.870 ;
        RECT 1401.780 966.125 1401.920 979.550 ;
        RECT 1401.710 965.755 1401.990 966.125 ;
        RECT 1402.630 965.755 1402.910 966.125 ;
        RECT 1402.700 904.245 1402.840 965.755 ;
        RECT 1401.710 903.875 1401.990 904.245 ;
        RECT 1402.630 903.875 1402.910 904.245 ;
        RECT 1401.720 903.730 1401.980 903.875 ;
        RECT 1402.640 903.730 1402.900 903.875 ;
        RECT 1402.700 807.150 1402.840 903.730 ;
        RECT 1402.640 806.830 1402.900 807.150 ;
        RECT 1401.720 758.890 1401.980 759.210 ;
        RECT 1401.780 735.490 1401.920 758.890 ;
        RECT 1401.780 735.350 1402.840 735.490 ;
        RECT 1402.700 669.450 1402.840 735.350 ;
        RECT 1402.640 669.130 1402.900 669.450 ;
        RECT 1402.640 620.850 1402.900 621.170 ;
        RECT 1402.700 590.085 1402.840 620.850 ;
        RECT 1402.630 589.715 1402.910 590.085 ;
        RECT 1401.710 524.435 1401.990 524.805 ;
        RECT 1401.780 517.470 1401.920 524.435 ;
        RECT 1401.720 517.150 1401.980 517.470 ;
        RECT 1401.720 469.210 1401.980 469.530 ;
        RECT 1401.780 428.050 1401.920 469.210 ;
        RECT 1401.720 427.730 1401.980 428.050 ;
        RECT 1402.640 427.730 1402.900 428.050 ;
        RECT 1402.700 386.230 1402.840 427.730 ;
        RECT 1402.640 385.910 1402.900 386.230 ;
        RECT 1401.720 347.490 1401.980 347.810 ;
        RECT 1401.780 331.150 1401.920 347.490 ;
        RECT 1401.720 330.830 1401.980 331.150 ;
        RECT 1401.720 282.890 1401.980 283.210 ;
        RECT 1401.780 259.070 1401.920 282.890 ;
        RECT 1401.720 258.750 1401.980 259.070 ;
        RECT 1402.640 186.330 1402.900 186.650 ;
        RECT 1402.700 138.030 1402.840 186.330 ;
        RECT 1402.640 137.710 1402.900 138.030 ;
        RECT 1401.720 89.770 1401.980 90.090 ;
        RECT 1401.780 35.690 1401.920 89.770 ;
        RECT 930.220 35.370 930.480 35.690 ;
        RECT 1401.720 35.370 1401.980 35.690 ;
        RECT 930.280 2.400 930.420 35.370 ;
        RECT 930.070 -4.800 930.630 2.400 ;
      LAYER via2 ;
        RECT 1401.710 1152.120 1401.990 1152.400 ;
        RECT 1402.630 1152.120 1402.910 1152.400 ;
        RECT 1401.710 965.800 1401.990 966.080 ;
        RECT 1402.630 965.800 1402.910 966.080 ;
        RECT 1401.710 903.920 1401.990 904.200 ;
        RECT 1402.630 903.920 1402.910 904.200 ;
        RECT 1402.630 589.760 1402.910 590.040 ;
        RECT 1401.710 524.480 1401.990 524.760 ;
      LAYER met3 ;
        RECT 1401.685 1152.410 1402.015 1152.425 ;
        RECT 1402.605 1152.410 1402.935 1152.425 ;
        RECT 1401.685 1152.110 1402.935 1152.410 ;
        RECT 1401.685 1152.095 1402.015 1152.110 ;
        RECT 1402.605 1152.095 1402.935 1152.110 ;
        RECT 1401.685 966.090 1402.015 966.105 ;
        RECT 1402.605 966.090 1402.935 966.105 ;
        RECT 1401.685 965.790 1402.935 966.090 ;
        RECT 1401.685 965.775 1402.015 965.790 ;
        RECT 1402.605 965.775 1402.935 965.790 ;
        RECT 1401.685 904.210 1402.015 904.225 ;
        RECT 1402.605 904.210 1402.935 904.225 ;
        RECT 1401.685 903.910 1402.935 904.210 ;
        RECT 1401.685 903.895 1402.015 903.910 ;
        RECT 1402.605 903.895 1402.935 903.910 ;
        RECT 1401.430 590.050 1401.810 590.060 ;
        RECT 1402.605 590.050 1402.935 590.065 ;
        RECT 1401.430 589.750 1402.935 590.050 ;
        RECT 1401.430 589.740 1401.810 589.750 ;
        RECT 1402.605 589.735 1402.935 589.750 ;
        RECT 1401.685 524.780 1402.015 524.785 ;
        RECT 1401.430 524.770 1402.015 524.780 ;
        RECT 1401.430 524.470 1402.240 524.770 ;
        RECT 1401.430 524.460 1402.015 524.470 ;
        RECT 1401.685 524.455 1402.015 524.460 ;
      LAYER via3 ;
        RECT 1401.460 589.740 1401.780 590.060 ;
        RECT 1401.460 524.460 1401.780 524.780 ;
      LAYER met4 ;
        RECT 1401.455 589.735 1401.785 590.065 ;
        RECT 1401.470 524.785 1401.770 589.735 ;
        RECT 1401.455 524.455 1401.785 524.785 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1402.150 1678.140 1402.470 1678.200 ;
        RECT 1404.450 1678.140 1404.770 1678.200 ;
        RECT 1402.150 1678.000 1404.770 1678.140 ;
        RECT 1402.150 1677.940 1402.470 1678.000 ;
        RECT 1404.450 1677.940 1404.770 1678.000 ;
        RECT 948.130 35.600 948.450 35.660 ;
        RECT 1402.150 35.600 1402.470 35.660 ;
        RECT 948.130 35.460 1402.470 35.600 ;
        RECT 948.130 35.400 948.450 35.460 ;
        RECT 1402.150 35.400 1402.470 35.460 ;
      LAYER via ;
        RECT 1402.180 1677.940 1402.440 1678.200 ;
        RECT 1404.480 1677.940 1404.740 1678.200 ;
        RECT 948.160 35.400 948.420 35.660 ;
        RECT 1402.180 35.400 1402.440 35.660 ;
      LAYER met2 ;
        RECT 1405.850 1700.410 1406.130 1704.000 ;
        RECT 1404.540 1700.270 1406.130 1700.410 ;
        RECT 1404.540 1678.230 1404.680 1700.270 ;
        RECT 1405.850 1700.000 1406.130 1700.270 ;
        RECT 1402.180 1677.910 1402.440 1678.230 ;
        RECT 1404.480 1677.910 1404.740 1678.230 ;
        RECT 1402.240 35.690 1402.380 1677.910 ;
        RECT 948.160 35.370 948.420 35.690 ;
        RECT 1402.180 35.370 1402.440 35.690 ;
        RECT 948.220 2.400 948.360 35.370 ;
        RECT 948.010 -4.800 948.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1403.145 1435.225 1403.315 1573.095 ;
        RECT 1403.605 1352.605 1403.775 1411.255 ;
        RECT 1403.145 1110.525 1403.315 1125.315 ;
        RECT 1403.145 855.525 1403.315 910.775 ;
        RECT 1403.145 711.025 1403.315 787.015 ;
        RECT 1403.605 572.645 1403.775 645.235 ;
        RECT 1403.605 338.045 1403.775 386.155 ;
        RECT 1403.145 179.605 1403.315 227.715 ;
      LAYER mcon ;
        RECT 1403.145 1572.925 1403.315 1573.095 ;
        RECT 1403.605 1411.085 1403.775 1411.255 ;
        RECT 1403.145 1125.145 1403.315 1125.315 ;
        RECT 1403.145 910.605 1403.315 910.775 ;
        RECT 1403.145 786.845 1403.315 787.015 ;
        RECT 1403.605 645.065 1403.775 645.235 ;
        RECT 1403.605 385.985 1403.775 386.155 ;
        RECT 1403.145 227.545 1403.315 227.715 ;
      LAYER met1 ;
        RECT 1403.530 1678.140 1403.850 1678.200 ;
        RECT 1406.750 1678.140 1407.070 1678.200 ;
        RECT 1403.530 1678.000 1407.070 1678.140 ;
        RECT 1403.530 1677.940 1403.850 1678.000 ;
        RECT 1406.750 1677.940 1407.070 1678.000 ;
        RECT 1404.450 1621.700 1404.770 1621.760 ;
        RECT 1405.370 1621.700 1405.690 1621.760 ;
        RECT 1404.450 1621.560 1405.690 1621.700 ;
        RECT 1404.450 1621.500 1404.770 1621.560 ;
        RECT 1405.370 1621.500 1405.690 1621.560 ;
        RECT 1403.530 1580.220 1403.850 1580.280 ;
        RECT 1404.450 1580.220 1404.770 1580.280 ;
        RECT 1403.530 1580.080 1404.770 1580.220 ;
        RECT 1403.530 1580.020 1403.850 1580.080 ;
        RECT 1404.450 1580.020 1404.770 1580.080 ;
        RECT 1403.085 1573.080 1403.375 1573.125 ;
        RECT 1403.530 1573.080 1403.850 1573.140 ;
        RECT 1403.085 1572.940 1403.850 1573.080 ;
        RECT 1403.085 1572.895 1403.375 1572.940 ;
        RECT 1403.530 1572.880 1403.850 1572.940 ;
        RECT 1403.085 1435.380 1403.375 1435.425 ;
        RECT 1403.530 1435.380 1403.850 1435.440 ;
        RECT 1403.085 1435.240 1403.850 1435.380 ;
        RECT 1403.085 1435.195 1403.375 1435.240 ;
        RECT 1403.530 1435.180 1403.850 1435.240 ;
        RECT 1403.530 1411.240 1403.850 1411.300 ;
        RECT 1403.335 1411.100 1403.850 1411.240 ;
        RECT 1403.530 1411.040 1403.850 1411.100 ;
        RECT 1403.530 1352.760 1403.850 1352.820 ;
        RECT 1403.335 1352.620 1403.850 1352.760 ;
        RECT 1403.530 1352.560 1403.850 1352.620 ;
        RECT 1403.530 1318.420 1403.850 1318.480 ;
        RECT 1403.160 1318.280 1403.850 1318.420 ;
        RECT 1403.160 1317.800 1403.300 1318.280 ;
        RECT 1403.530 1318.220 1403.850 1318.280 ;
        RECT 1403.070 1317.540 1403.390 1317.800 ;
        RECT 1402.150 1259.260 1402.470 1259.320 ;
        RECT 1403.070 1259.260 1403.390 1259.320 ;
        RECT 1402.150 1259.120 1403.390 1259.260 ;
        RECT 1402.150 1259.060 1402.470 1259.120 ;
        RECT 1403.070 1259.060 1403.390 1259.120 ;
        RECT 1403.070 1125.300 1403.390 1125.360 ;
        RECT 1402.875 1125.160 1403.390 1125.300 ;
        RECT 1403.070 1125.100 1403.390 1125.160 ;
        RECT 1403.070 1110.680 1403.390 1110.740 ;
        RECT 1402.875 1110.540 1403.390 1110.680 ;
        RECT 1403.070 1110.480 1403.390 1110.540 ;
        RECT 1403.530 918.240 1403.850 918.300 ;
        RECT 1403.160 918.100 1403.850 918.240 ;
        RECT 1403.160 917.960 1403.300 918.100 ;
        RECT 1403.530 918.040 1403.850 918.100 ;
        RECT 1403.070 917.700 1403.390 917.960 ;
        RECT 1403.070 910.760 1403.390 910.820 ;
        RECT 1402.875 910.620 1403.390 910.760 ;
        RECT 1403.070 910.560 1403.390 910.620 ;
        RECT 1403.085 855.680 1403.375 855.725 ;
        RECT 1403.530 855.680 1403.850 855.740 ;
        RECT 1403.085 855.540 1403.850 855.680 ;
        RECT 1403.085 855.495 1403.375 855.540 ;
        RECT 1403.530 855.480 1403.850 855.540 ;
        RECT 1403.085 787.000 1403.375 787.045 ;
        RECT 1403.530 787.000 1403.850 787.060 ;
        RECT 1403.085 786.860 1403.850 787.000 ;
        RECT 1403.085 786.815 1403.375 786.860 ;
        RECT 1403.530 786.800 1403.850 786.860 ;
        RECT 1403.070 711.180 1403.390 711.240 ;
        RECT 1402.875 711.040 1403.390 711.180 ;
        RECT 1403.070 710.980 1403.390 711.040 ;
        RECT 1403.070 645.220 1403.390 645.280 ;
        RECT 1403.545 645.220 1403.835 645.265 ;
        RECT 1403.070 645.080 1403.835 645.220 ;
        RECT 1403.070 645.020 1403.390 645.080 ;
        RECT 1403.545 645.035 1403.835 645.080 ;
        RECT 1403.530 572.800 1403.850 572.860 ;
        RECT 1403.335 572.660 1403.850 572.800 ;
        RECT 1403.530 572.600 1403.850 572.660 ;
        RECT 1403.070 476.240 1403.390 476.300 ;
        RECT 1403.530 476.240 1403.850 476.300 ;
        RECT 1403.070 476.100 1403.850 476.240 ;
        RECT 1403.070 476.040 1403.390 476.100 ;
        RECT 1403.530 476.040 1403.850 476.100 ;
        RECT 1403.070 448.500 1403.390 448.760 ;
        RECT 1403.160 448.020 1403.300 448.500 ;
        RECT 1403.530 448.020 1403.850 448.080 ;
        RECT 1403.160 447.880 1403.850 448.020 ;
        RECT 1403.530 447.820 1403.850 447.880 ;
        RECT 1403.530 386.140 1403.850 386.200 ;
        RECT 1403.335 386.000 1403.850 386.140 ;
        RECT 1403.530 385.940 1403.850 386.000 ;
        RECT 1403.530 338.200 1403.850 338.260 ;
        RECT 1403.335 338.060 1403.850 338.200 ;
        RECT 1403.530 338.000 1403.850 338.060 ;
        RECT 1402.150 331.060 1402.470 331.120 ;
        RECT 1403.530 331.060 1403.850 331.120 ;
        RECT 1402.150 330.920 1403.850 331.060 ;
        RECT 1402.150 330.860 1402.470 330.920 ;
        RECT 1403.530 330.860 1403.850 330.920 ;
        RECT 1403.070 235.180 1403.390 235.240 ;
        RECT 1403.070 235.040 1403.760 235.180 ;
        RECT 1403.070 234.980 1403.390 235.040 ;
        RECT 1403.620 234.900 1403.760 235.040 ;
        RECT 1403.530 234.640 1403.850 234.900 ;
        RECT 1403.085 227.700 1403.375 227.745 ;
        RECT 1403.530 227.700 1403.850 227.760 ;
        RECT 1403.085 227.560 1403.850 227.700 ;
        RECT 1403.085 227.515 1403.375 227.560 ;
        RECT 1403.530 227.500 1403.850 227.560 ;
        RECT 1403.070 179.760 1403.390 179.820 ;
        RECT 1402.875 179.620 1403.390 179.760 ;
        RECT 1403.070 179.560 1403.390 179.620 ;
        RECT 1402.610 83.200 1402.930 83.260 ;
        RECT 1403.070 83.200 1403.390 83.260 ;
        RECT 1402.610 83.060 1403.390 83.200 ;
        RECT 1402.610 83.000 1402.930 83.060 ;
        RECT 1403.070 83.000 1403.390 83.060 ;
        RECT 948.130 35.260 948.450 35.320 ;
        RECT 1403.070 35.260 1403.390 35.320 ;
        RECT 948.130 35.120 1403.390 35.260 ;
        RECT 948.130 35.060 948.450 35.120 ;
        RECT 1403.070 35.060 1403.390 35.120 ;
      LAYER via ;
        RECT 1403.560 1677.940 1403.820 1678.200 ;
        RECT 1406.780 1677.940 1407.040 1678.200 ;
        RECT 1404.480 1621.500 1404.740 1621.760 ;
        RECT 1405.400 1621.500 1405.660 1621.760 ;
        RECT 1403.560 1580.020 1403.820 1580.280 ;
        RECT 1404.480 1580.020 1404.740 1580.280 ;
        RECT 1403.560 1572.880 1403.820 1573.140 ;
        RECT 1403.560 1435.180 1403.820 1435.440 ;
        RECT 1403.560 1411.040 1403.820 1411.300 ;
        RECT 1403.560 1352.560 1403.820 1352.820 ;
        RECT 1403.560 1318.220 1403.820 1318.480 ;
        RECT 1403.100 1317.540 1403.360 1317.800 ;
        RECT 1402.180 1259.060 1402.440 1259.320 ;
        RECT 1403.100 1259.060 1403.360 1259.320 ;
        RECT 1403.100 1125.100 1403.360 1125.360 ;
        RECT 1403.100 1110.480 1403.360 1110.740 ;
        RECT 1403.560 918.040 1403.820 918.300 ;
        RECT 1403.100 917.700 1403.360 917.960 ;
        RECT 1403.100 910.560 1403.360 910.820 ;
        RECT 1403.560 855.480 1403.820 855.740 ;
        RECT 1403.560 786.800 1403.820 787.060 ;
        RECT 1403.100 710.980 1403.360 711.240 ;
        RECT 1403.100 645.020 1403.360 645.280 ;
        RECT 1403.560 572.600 1403.820 572.860 ;
        RECT 1403.100 476.040 1403.360 476.300 ;
        RECT 1403.560 476.040 1403.820 476.300 ;
        RECT 1403.100 448.500 1403.360 448.760 ;
        RECT 1403.560 447.820 1403.820 448.080 ;
        RECT 1403.560 385.940 1403.820 386.200 ;
        RECT 1403.560 338.000 1403.820 338.260 ;
        RECT 1402.180 330.860 1402.440 331.120 ;
        RECT 1403.560 330.860 1403.820 331.120 ;
        RECT 1403.100 234.980 1403.360 235.240 ;
        RECT 1403.560 234.640 1403.820 234.900 ;
        RECT 1403.560 227.500 1403.820 227.760 ;
        RECT 1403.100 179.560 1403.360 179.820 ;
        RECT 1402.640 83.000 1402.900 83.260 ;
        RECT 1403.100 83.000 1403.360 83.260 ;
        RECT 948.160 35.060 948.420 35.320 ;
        RECT 1403.100 35.060 1403.360 35.320 ;
      LAYER met2 ;
        RECT 1406.770 1700.000 1407.050 1704.000 ;
        RECT 1406.840 1678.230 1406.980 1700.000 ;
        RECT 1403.560 1677.910 1403.820 1678.230 ;
        RECT 1406.780 1677.910 1407.040 1678.230 ;
        RECT 1403.620 1669.925 1403.760 1677.910 ;
        RECT 1403.550 1669.555 1403.830 1669.925 ;
        RECT 1405.390 1669.555 1405.670 1669.925 ;
        RECT 1405.460 1621.790 1405.600 1669.555 ;
        RECT 1404.480 1621.470 1404.740 1621.790 ;
        RECT 1405.400 1621.470 1405.660 1621.790 ;
        RECT 1404.540 1580.310 1404.680 1621.470 ;
        RECT 1403.560 1579.990 1403.820 1580.310 ;
        RECT 1404.480 1579.990 1404.740 1580.310 ;
        RECT 1403.620 1573.170 1403.760 1579.990 ;
        RECT 1403.560 1572.850 1403.820 1573.170 ;
        RECT 1403.560 1435.150 1403.820 1435.470 ;
        RECT 1403.620 1411.330 1403.760 1435.150 ;
        RECT 1403.560 1411.010 1403.820 1411.330 ;
        RECT 1403.560 1352.530 1403.820 1352.850 ;
        RECT 1403.620 1318.510 1403.760 1352.530 ;
        RECT 1403.560 1318.190 1403.820 1318.510 ;
        RECT 1403.100 1317.510 1403.360 1317.830 ;
        RECT 1403.160 1259.350 1403.300 1317.510 ;
        RECT 1402.180 1259.030 1402.440 1259.350 ;
        RECT 1403.100 1259.030 1403.360 1259.350 ;
        RECT 1402.240 1235.405 1402.380 1259.030 ;
        RECT 1402.170 1235.035 1402.450 1235.405 ;
        RECT 1404.470 1235.035 1404.750 1235.405 ;
        RECT 1404.540 1193.925 1404.680 1235.035 ;
        RECT 1403.550 1193.555 1403.830 1193.925 ;
        RECT 1404.470 1193.555 1404.750 1193.925 ;
        RECT 1403.620 1176.810 1403.760 1193.555 ;
        RECT 1403.160 1176.670 1403.760 1176.810 ;
        RECT 1403.160 1125.390 1403.300 1176.670 ;
        RECT 1403.100 1125.070 1403.360 1125.390 ;
        RECT 1403.100 1110.450 1403.360 1110.770 ;
        RECT 1403.160 1104.165 1403.300 1110.450 ;
        RECT 1403.090 1103.795 1403.370 1104.165 ;
        RECT 1403.550 1103.115 1403.830 1103.485 ;
        RECT 1403.620 918.330 1403.760 1103.115 ;
        RECT 1403.560 918.010 1403.820 918.330 ;
        RECT 1403.100 917.670 1403.360 917.990 ;
        RECT 1403.160 910.850 1403.300 917.670 ;
        RECT 1403.100 910.530 1403.360 910.850 ;
        RECT 1403.560 855.450 1403.820 855.770 ;
        RECT 1403.620 787.090 1403.760 855.450 ;
        RECT 1403.560 786.770 1403.820 787.090 ;
        RECT 1403.100 710.950 1403.360 711.270 ;
        RECT 1403.160 645.310 1403.300 710.950 ;
        RECT 1403.100 644.990 1403.360 645.310 ;
        RECT 1403.560 572.570 1403.820 572.890 ;
        RECT 1403.620 476.330 1403.760 572.570 ;
        RECT 1403.100 476.010 1403.360 476.330 ;
        RECT 1403.560 476.010 1403.820 476.330 ;
        RECT 1403.160 448.790 1403.300 476.010 ;
        RECT 1403.100 448.470 1403.360 448.790 ;
        RECT 1403.560 447.790 1403.820 448.110 ;
        RECT 1403.620 386.230 1403.760 447.790 ;
        RECT 1403.560 385.910 1403.820 386.230 ;
        RECT 1403.560 337.970 1403.820 338.290 ;
        RECT 1403.620 331.150 1403.760 337.970 ;
        RECT 1402.180 330.830 1402.440 331.150 ;
        RECT 1403.560 330.830 1403.820 331.150 ;
        RECT 1402.240 283.405 1402.380 330.830 ;
        RECT 1402.170 283.035 1402.450 283.405 ;
        RECT 1403.090 283.035 1403.370 283.405 ;
        RECT 1403.160 235.270 1403.300 283.035 ;
        RECT 1403.100 234.950 1403.360 235.270 ;
        RECT 1403.560 234.610 1403.820 234.930 ;
        RECT 1403.620 227.790 1403.760 234.610 ;
        RECT 1403.560 227.470 1403.820 227.790 ;
        RECT 1403.100 179.530 1403.360 179.850 ;
        RECT 1403.160 137.090 1403.300 179.530 ;
        RECT 1402.700 136.950 1403.300 137.090 ;
        RECT 1402.700 83.290 1402.840 136.950 ;
        RECT 1402.640 82.970 1402.900 83.290 ;
        RECT 1403.100 82.970 1403.360 83.290 ;
        RECT 1403.160 35.350 1403.300 82.970 ;
        RECT 948.160 35.030 948.420 35.350 ;
        RECT 1403.100 35.030 1403.360 35.350 ;
        RECT 948.220 2.400 948.360 35.030 ;
        RECT 948.010 -4.800 948.570 2.400 ;
      LAYER via2 ;
        RECT 1403.550 1669.600 1403.830 1669.880 ;
        RECT 1405.390 1669.600 1405.670 1669.880 ;
        RECT 1402.170 1235.080 1402.450 1235.360 ;
        RECT 1404.470 1235.080 1404.750 1235.360 ;
        RECT 1403.550 1193.600 1403.830 1193.880 ;
        RECT 1404.470 1193.600 1404.750 1193.880 ;
        RECT 1403.090 1103.840 1403.370 1104.120 ;
        RECT 1403.550 1103.160 1403.830 1103.440 ;
        RECT 1402.170 283.080 1402.450 283.360 ;
        RECT 1403.090 283.080 1403.370 283.360 ;
      LAYER met3 ;
        RECT 1403.525 1669.890 1403.855 1669.905 ;
        RECT 1405.365 1669.890 1405.695 1669.905 ;
        RECT 1403.525 1669.590 1405.695 1669.890 ;
        RECT 1403.525 1669.575 1403.855 1669.590 ;
        RECT 1405.365 1669.575 1405.695 1669.590 ;
        RECT 1402.145 1235.370 1402.475 1235.385 ;
        RECT 1404.445 1235.370 1404.775 1235.385 ;
        RECT 1402.145 1235.070 1404.775 1235.370 ;
        RECT 1402.145 1235.055 1402.475 1235.070 ;
        RECT 1404.445 1235.055 1404.775 1235.070 ;
        RECT 1403.525 1193.890 1403.855 1193.905 ;
        RECT 1404.445 1193.890 1404.775 1193.905 ;
        RECT 1403.525 1193.590 1404.775 1193.890 ;
        RECT 1403.525 1193.575 1403.855 1193.590 ;
        RECT 1404.445 1193.575 1404.775 1193.590 ;
        RECT 1403.065 1104.130 1403.395 1104.145 ;
        RECT 1403.065 1103.815 1403.610 1104.130 ;
        RECT 1403.310 1103.465 1403.610 1103.815 ;
        RECT 1403.310 1103.150 1403.855 1103.465 ;
        RECT 1403.525 1103.135 1403.855 1103.150 ;
        RECT 1402.145 283.370 1402.475 283.385 ;
        RECT 1403.065 283.370 1403.395 283.385 ;
        RECT 1402.145 283.070 1403.395 283.370 ;
        RECT 1402.145 283.055 1402.475 283.070 ;
        RECT 1403.065 283.055 1403.395 283.070 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 0.300 ;
=======
      LAYER met1 ;
        RECT 966.070 34.920 966.390 34.980 ;
        RECT 1409.050 34.920 1409.370 34.980 ;
        RECT 966.070 34.780 1409.370 34.920 ;
        RECT 966.070 34.720 966.390 34.780 ;
        RECT 1409.050 34.720 1409.370 34.780 ;
      LAYER via ;
        RECT 966.100 34.720 966.360 34.980 ;
        RECT 1409.080 34.720 1409.340 34.980 ;
      LAYER met2 ;
        RECT 1411.370 1700.410 1411.650 1704.000 ;
        RECT 1410.520 1700.270 1411.650 1700.410 ;
        RECT 1410.520 1678.140 1410.660 1700.270 ;
        RECT 1411.370 1700.000 1411.650 1700.270 ;
        RECT 1409.140 1678.000 1410.660 1678.140 ;
        RECT 1409.140 35.010 1409.280 1678.000 ;
        RECT 966.100 34.690 966.360 35.010 ;
        RECT 1409.080 34.690 1409.340 35.010 ;
        RECT 966.160 2.400 966.300 34.690 ;
        RECT 965.950 -4.800 966.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 0.300 ;
=======
      LAYER met1 ;
        RECT 986.310 1570.020 986.630 1570.080 ;
        RECT 1415.950 1570.020 1416.270 1570.080 ;
        RECT 986.310 1569.880 1416.270 1570.020 ;
        RECT 986.310 1569.820 986.630 1569.880 ;
        RECT 1415.950 1569.820 1416.270 1569.880 ;
      LAYER via ;
        RECT 986.340 1569.820 986.600 1570.080 ;
        RECT 1415.980 1569.820 1416.240 1570.080 ;
      LAYER met2 ;
        RECT 1416.430 1700.410 1416.710 1704.000 ;
        RECT 1416.040 1700.270 1416.710 1700.410 ;
        RECT 1416.040 1570.110 1416.180 1700.270 ;
        RECT 1416.430 1700.000 1416.710 1700.270 ;
        RECT 986.340 1569.790 986.600 1570.110 ;
        RECT 1415.980 1569.790 1416.240 1570.110 ;
        RECT 986.400 16.730 986.540 1569.790 ;
        RECT 984.100 16.590 986.540 16.730 ;
        RECT 984.100 2.400 984.240 16.590 ;
        RECT 983.890 -4.800 984.450 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 0.300 ;
=======
      LAYER met1 ;
        RECT 668.450 1548.940 668.770 1549.000 ;
        RECT 1326.710 1548.940 1327.030 1549.000 ;
        RECT 668.450 1548.800 1327.030 1548.940 ;
        RECT 668.450 1548.740 668.770 1548.800 ;
        RECT 1326.710 1548.740 1327.030 1548.800 ;
        RECT 662.930 2.960 663.250 3.020 ;
        RECT 668.450 2.960 668.770 3.020 ;
        RECT 662.930 2.820 668.770 2.960 ;
        RECT 662.930 2.760 663.250 2.820 ;
        RECT 668.450 2.760 668.770 2.820 ;
      LAYER via ;
        RECT 668.480 1548.740 668.740 1549.000 ;
        RECT 1326.740 1548.740 1327.000 1549.000 ;
        RECT 662.960 2.760 663.220 3.020 ;
        RECT 668.480 2.760 668.740 3.020 ;
      LAYER met2 ;
        RECT 1329.490 1701.090 1329.770 1704.000 ;
        RECT 1328.180 1700.950 1329.770 1701.090 ;
        RECT 1328.180 1695.650 1328.320 1700.950 ;
        RECT 1329.490 1700.000 1329.770 1700.950 ;
        RECT 1327.260 1695.510 1328.320 1695.650 ;
        RECT 1327.260 1666.410 1327.400 1695.510 ;
        RECT 1326.800 1666.270 1327.400 1666.410 ;
        RECT 1326.800 1549.030 1326.940 1666.270 ;
        RECT 668.480 1548.710 668.740 1549.030 ;
        RECT 1326.740 1548.710 1327.000 1549.030 ;
        RECT 668.540 3.050 668.680 1548.710 ;
        RECT 662.960 2.730 663.220 3.050 ;
        RECT 668.480 2.730 668.740 3.050 ;
        RECT 663.020 2.400 663.160 2.730 ;
        RECT 662.810 -4.800 663.370 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 0.300 ;
=======
      LAYER li1 ;
        RECT 1416.025 1442.025 1416.195 1449.675 ;
        RECT 1416.485 1200.625 1416.655 1207.595 ;
        RECT 1416.485 1074.825 1416.655 1097.095 ;
        RECT 1416.025 855.525 1416.195 903.975 ;
        RECT 1416.485 688.245 1416.655 717.655 ;
        RECT 1416.025 425.085 1416.195 517.395 ;
        RECT 1416.025 324.445 1416.195 414.035 ;
        RECT 1416.025 228.225 1416.195 275.995 ;
        RECT 1416.025 179.605 1416.195 227.715 ;
      LAYER mcon ;
        RECT 1416.025 1449.505 1416.195 1449.675 ;
        RECT 1416.485 1207.425 1416.655 1207.595 ;
        RECT 1416.485 1096.925 1416.655 1097.095 ;
        RECT 1416.025 903.805 1416.195 903.975 ;
        RECT 1416.485 717.485 1416.655 717.655 ;
        RECT 1416.025 517.225 1416.195 517.395 ;
        RECT 1416.025 413.865 1416.195 414.035 ;
        RECT 1416.025 275.825 1416.195 275.995 ;
        RECT 1416.025 227.545 1416.195 227.715 ;
      LAYER met1 ;
        RECT 1416.410 1635.640 1416.730 1635.700 ;
        RECT 1419.630 1635.640 1419.950 1635.700 ;
        RECT 1416.410 1635.500 1419.950 1635.640 ;
        RECT 1416.410 1635.440 1416.730 1635.500 ;
        RECT 1419.630 1635.440 1419.950 1635.500 ;
        RECT 1415.965 1449.660 1416.255 1449.705 ;
        RECT 1416.410 1449.660 1416.730 1449.720 ;
        RECT 1415.965 1449.520 1416.730 1449.660 ;
        RECT 1415.965 1449.475 1416.255 1449.520 ;
        RECT 1416.410 1449.460 1416.730 1449.520 ;
        RECT 1415.950 1442.180 1416.270 1442.240 ;
        RECT 1415.755 1442.040 1416.270 1442.180 ;
        RECT 1415.950 1441.980 1416.270 1442.040 ;
        RECT 1416.870 1297.680 1417.190 1297.740 ;
        RECT 1416.040 1297.540 1417.190 1297.680 ;
        RECT 1416.040 1297.400 1416.180 1297.540 ;
        RECT 1416.870 1297.480 1417.190 1297.540 ;
        RECT 1415.950 1297.140 1416.270 1297.400 ;
        RECT 1416.870 1249.200 1417.190 1249.460 ;
        RECT 1416.410 1249.060 1416.730 1249.120 ;
        RECT 1416.960 1249.060 1417.100 1249.200 ;
        RECT 1416.410 1248.920 1417.100 1249.060 ;
        RECT 1416.410 1248.860 1416.730 1248.920 ;
        RECT 1416.410 1207.580 1416.730 1207.640 ;
        RECT 1416.215 1207.440 1416.730 1207.580 ;
        RECT 1416.410 1207.380 1416.730 1207.440 ;
        RECT 1416.410 1200.780 1416.730 1200.840 ;
        RECT 1416.215 1200.640 1416.730 1200.780 ;
        RECT 1416.410 1200.580 1416.730 1200.640 ;
        RECT 1416.410 1152.300 1416.730 1152.560 ;
        RECT 1416.500 1151.880 1416.640 1152.300 ;
        RECT 1416.410 1151.620 1416.730 1151.880 ;
        RECT 1416.410 1145.360 1416.730 1145.420 ;
        RECT 1417.330 1145.360 1417.650 1145.420 ;
        RECT 1416.410 1145.220 1417.650 1145.360 ;
        RECT 1416.410 1145.160 1416.730 1145.220 ;
        RECT 1417.330 1145.160 1417.650 1145.220 ;
        RECT 1416.410 1097.080 1416.730 1097.140 ;
        RECT 1416.215 1096.940 1416.730 1097.080 ;
        RECT 1416.410 1096.880 1416.730 1096.940 ;
        RECT 1416.425 1074.980 1416.715 1075.025 ;
        RECT 1416.870 1074.980 1417.190 1075.040 ;
        RECT 1416.425 1074.840 1417.190 1074.980 ;
        RECT 1416.425 1074.795 1416.715 1074.840 ;
        RECT 1416.870 1074.780 1417.190 1074.840 ;
        RECT 1416.870 1048.800 1417.190 1048.860 ;
        RECT 1417.790 1048.800 1418.110 1048.860 ;
        RECT 1416.870 1048.660 1418.110 1048.800 ;
        RECT 1416.870 1048.600 1417.190 1048.660 ;
        RECT 1417.790 1048.600 1418.110 1048.660 ;
        RECT 1415.950 917.900 1416.270 917.960 ;
        RECT 1416.870 917.900 1417.190 917.960 ;
        RECT 1415.950 917.760 1417.190 917.900 ;
        RECT 1415.950 917.700 1416.270 917.760 ;
        RECT 1416.870 917.700 1417.190 917.760 ;
        RECT 1415.950 903.960 1416.270 904.020 ;
        RECT 1415.755 903.820 1416.270 903.960 ;
        RECT 1415.950 903.760 1416.270 903.820 ;
        RECT 1415.965 855.680 1416.255 855.725 ;
        RECT 1416.870 855.680 1417.190 855.740 ;
        RECT 1415.965 855.540 1417.190 855.680 ;
        RECT 1415.965 855.495 1416.255 855.540 ;
        RECT 1416.870 855.480 1417.190 855.540 ;
        RECT 1415.950 814.200 1416.270 814.260 ;
        RECT 1416.870 814.200 1417.190 814.260 ;
        RECT 1415.950 814.060 1417.190 814.200 ;
        RECT 1415.950 814.000 1416.270 814.060 ;
        RECT 1416.870 814.000 1417.190 814.060 ;
        RECT 1415.950 724.440 1416.270 724.500 ;
        RECT 1416.870 724.440 1417.190 724.500 ;
        RECT 1415.950 724.300 1417.190 724.440 ;
        RECT 1415.950 724.240 1416.270 724.300 ;
        RECT 1416.870 724.240 1417.190 724.300 ;
        RECT 1416.425 717.640 1416.715 717.685 ;
        RECT 1416.870 717.640 1417.190 717.700 ;
        RECT 1416.425 717.500 1417.190 717.640 ;
        RECT 1416.425 717.455 1416.715 717.500 ;
        RECT 1416.870 717.440 1417.190 717.500 ;
        RECT 1416.410 688.400 1416.730 688.460 ;
        RECT 1416.215 688.260 1416.730 688.400 ;
        RECT 1416.410 688.200 1416.730 688.260 ;
        RECT 1416.410 525.340 1416.730 525.600 ;
        RECT 1416.500 524.920 1416.640 525.340 ;
        RECT 1416.410 524.660 1416.730 524.920 ;
        RECT 1415.965 517.380 1416.255 517.425 ;
        RECT 1416.410 517.380 1416.730 517.440 ;
        RECT 1415.965 517.240 1416.730 517.380 ;
        RECT 1415.965 517.195 1416.255 517.240 ;
        RECT 1416.410 517.180 1416.730 517.240 ;
        RECT 1415.950 425.240 1416.270 425.300 ;
        RECT 1415.755 425.100 1416.270 425.240 ;
        RECT 1415.950 425.040 1416.270 425.100 ;
        RECT 1415.950 414.020 1416.270 414.080 ;
        RECT 1415.755 413.880 1416.270 414.020 ;
        RECT 1415.950 413.820 1416.270 413.880 ;
        RECT 1415.965 324.600 1416.255 324.645 ;
        RECT 1416.410 324.600 1416.730 324.660 ;
        RECT 1415.965 324.460 1416.730 324.600 ;
        RECT 1415.965 324.415 1416.255 324.460 ;
        RECT 1416.410 324.400 1416.730 324.460 ;
        RECT 1415.965 275.980 1416.255 276.025 ;
        RECT 1416.870 275.980 1417.190 276.040 ;
        RECT 1415.965 275.840 1417.190 275.980 ;
        RECT 1415.965 275.795 1416.255 275.840 ;
        RECT 1416.870 275.780 1417.190 275.840 ;
        RECT 1415.950 228.380 1416.270 228.440 ;
        RECT 1415.755 228.240 1416.270 228.380 ;
        RECT 1415.950 228.180 1416.270 228.240 ;
        RECT 1415.950 227.700 1416.270 227.760 ;
        RECT 1415.755 227.560 1416.270 227.700 ;
        RECT 1415.950 227.500 1416.270 227.560 ;
        RECT 1415.950 179.760 1416.270 179.820 ;
        RECT 1415.755 179.620 1416.270 179.760 ;
        RECT 1415.950 179.560 1416.270 179.620 ;
        RECT 1416.410 137.740 1416.730 138.000 ;
        RECT 1416.500 137.320 1416.640 137.740 ;
        RECT 1416.410 137.060 1416.730 137.320 ;
        RECT 1007.010 49.540 1007.330 49.600 ;
        RECT 1416.410 49.540 1416.730 49.600 ;
        RECT 1007.010 49.400 1416.730 49.540 ;
        RECT 1007.010 49.340 1007.330 49.400 ;
        RECT 1416.410 49.340 1416.730 49.400 ;
=======
      LAYER met1 ;
        RECT 1007.010 1666.920 1007.330 1666.980 ;
        RECT 1421.470 1666.920 1421.790 1666.980 ;
        RECT 1007.010 1666.780 1421.790 1666.920 ;
        RECT 1007.010 1666.720 1007.330 1666.780 ;
        RECT 1421.470 1666.720 1421.790 1666.780 ;
>>>>>>> re-updated local openlane
        RECT 1001.950 2.960 1002.270 3.020 ;
        RECT 1007.010 2.960 1007.330 3.020 ;
        RECT 1001.950 2.820 1007.330 2.960 ;
        RECT 1001.950 2.760 1002.270 2.820 ;
        RECT 1007.010 2.760 1007.330 2.820 ;
      LAYER via ;
        RECT 1007.040 1666.720 1007.300 1666.980 ;
        RECT 1421.500 1666.720 1421.760 1666.980 ;
        RECT 1001.980 2.760 1002.240 3.020 ;
        RECT 1007.040 2.760 1007.300 3.020 ;
      LAYER met2 ;
        RECT 1421.490 1700.000 1421.770 1704.000 ;
        RECT 1421.560 1667.010 1421.700 1700.000 ;
        RECT 1007.040 1666.690 1007.300 1667.010 ;
        RECT 1421.500 1666.690 1421.760 1667.010 ;
        RECT 1007.100 3.050 1007.240 1666.690 ;
        RECT 1001.980 2.730 1002.240 3.050 ;
        RECT 1007.040 2.730 1007.300 3.050 ;
        RECT 1002.040 2.400 1002.180 2.730 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1416.430 1200.400 1416.710 1200.680 ;
        RECT 1416.430 1199.720 1416.710 1200.000 ;
        RECT 1416.430 1097.040 1416.710 1097.320 ;
        RECT 1417.350 1097.040 1417.630 1097.320 ;
        RECT 1416.430 1000.480 1416.710 1000.760 ;
        RECT 1417.810 1000.480 1418.090 1000.760 ;
        RECT 1415.970 724.400 1416.250 724.680 ;
        RECT 1416.890 724.400 1417.170 724.680 ;
        RECT 1416.430 573.440 1416.710 573.720 ;
        RECT 1415.970 572.760 1416.250 573.040 ;
      LAYER met3 ;
        RECT 1416.405 1200.690 1416.735 1200.705 ;
        RECT 1416.190 1200.375 1416.735 1200.690 ;
        RECT 1416.190 1200.025 1416.490 1200.375 ;
        RECT 1416.190 1199.710 1416.735 1200.025 ;
        RECT 1416.405 1199.695 1416.735 1199.710 ;
        RECT 1416.405 1097.330 1416.735 1097.345 ;
        RECT 1417.325 1097.330 1417.655 1097.345 ;
        RECT 1416.405 1097.030 1417.655 1097.330 ;
        RECT 1416.405 1097.015 1416.735 1097.030 ;
        RECT 1417.325 1097.015 1417.655 1097.030 ;
        RECT 1416.405 1000.770 1416.735 1000.785 ;
        RECT 1417.785 1000.770 1418.115 1000.785 ;
        RECT 1416.405 1000.470 1418.115 1000.770 ;
        RECT 1416.405 1000.455 1416.735 1000.470 ;
        RECT 1417.785 1000.455 1418.115 1000.470 ;
        RECT 1415.945 724.690 1416.275 724.705 ;
        RECT 1416.865 724.690 1417.195 724.705 ;
        RECT 1415.945 724.390 1417.195 724.690 ;
        RECT 1415.945 724.375 1416.275 724.390 ;
        RECT 1416.865 724.375 1417.195 724.390 ;
        RECT 1416.405 573.730 1416.735 573.745 ;
        RECT 1416.190 573.415 1416.735 573.730 ;
        RECT 1416.190 573.065 1416.490 573.415 ;
        RECT 1415.945 572.750 1416.490 573.065 ;
        RECT 1415.945 572.735 1416.275 572.750 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 0.300 ;
=======
      LAYER li1 ;
        RECT 1423.385 1635.485 1423.555 1683.595 ;
        RECT 1423.385 1442.025 1423.555 1490.475 ;
        RECT 1423.845 1352.605 1424.015 1400.715 ;
        RECT 1423.385 814.385 1423.555 862.495 ;
        RECT 1422.925 427.805 1423.095 475.915 ;
        RECT 1423.385 49.045 1423.555 113.815 ;
      LAYER mcon ;
        RECT 1423.385 1683.425 1423.555 1683.595 ;
        RECT 1423.385 1490.305 1423.555 1490.475 ;
        RECT 1423.845 1400.545 1424.015 1400.715 ;
        RECT 1423.385 862.325 1423.555 862.495 ;
        RECT 1422.925 475.745 1423.095 475.915 ;
        RECT 1423.385 113.645 1423.555 113.815 ;
      LAYER met1 ;
        RECT 1423.325 1683.580 1423.615 1683.625 ;
        RECT 1424.230 1683.580 1424.550 1683.640 ;
        RECT 1423.325 1683.440 1424.550 1683.580 ;
        RECT 1423.325 1683.395 1423.615 1683.440 ;
        RECT 1424.230 1683.380 1424.550 1683.440 ;
        RECT 1423.310 1635.640 1423.630 1635.700 ;
        RECT 1423.115 1635.500 1423.630 1635.640 ;
        RECT 1423.310 1635.440 1423.630 1635.500 ;
        RECT 1423.310 1545.880 1423.630 1545.940 ;
        RECT 1423.770 1545.880 1424.090 1545.940 ;
        RECT 1423.310 1545.740 1424.090 1545.880 ;
        RECT 1423.310 1545.680 1423.630 1545.740 ;
        RECT 1423.770 1545.680 1424.090 1545.740 ;
        RECT 1423.325 1490.460 1423.615 1490.505 ;
        RECT 1423.770 1490.460 1424.090 1490.520 ;
        RECT 1423.325 1490.320 1424.090 1490.460 ;
        RECT 1423.325 1490.275 1423.615 1490.320 ;
        RECT 1423.770 1490.260 1424.090 1490.320 ;
        RECT 1423.310 1442.180 1423.630 1442.240 ;
        RECT 1423.115 1442.040 1423.630 1442.180 ;
        RECT 1423.310 1441.980 1423.630 1442.040 ;
        RECT 1423.770 1400.700 1424.090 1400.760 ;
        RECT 1423.575 1400.560 1424.090 1400.700 ;
        RECT 1423.770 1400.500 1424.090 1400.560 ;
        RECT 1423.770 1352.760 1424.090 1352.820 ;
        RECT 1423.575 1352.620 1424.090 1352.760 ;
        RECT 1423.770 1352.560 1424.090 1352.620 ;
        RECT 1423.310 1303.940 1423.630 1304.200 ;
        RECT 1423.400 1303.800 1423.540 1303.940 ;
        RECT 1423.770 1303.800 1424.090 1303.860 ;
        RECT 1423.400 1303.660 1424.090 1303.800 ;
        RECT 1423.770 1303.600 1424.090 1303.660 ;
        RECT 1423.770 1159.640 1424.090 1159.700 ;
        RECT 1423.400 1159.500 1424.090 1159.640 ;
        RECT 1423.400 1159.360 1423.540 1159.500 ;
        RECT 1423.770 1159.440 1424.090 1159.500 ;
        RECT 1423.310 1159.100 1423.630 1159.360 ;
        RECT 1423.770 966.520 1424.090 966.580 ;
        RECT 1423.400 966.380 1424.090 966.520 ;
        RECT 1423.400 966.240 1423.540 966.380 ;
        RECT 1423.770 966.320 1424.090 966.380 ;
        RECT 1423.310 965.980 1423.630 966.240 ;
        RECT 1423.325 862.480 1423.615 862.525 ;
        RECT 1423.770 862.480 1424.090 862.540 ;
        RECT 1423.325 862.340 1424.090 862.480 ;
        RECT 1423.325 862.295 1423.615 862.340 ;
        RECT 1423.770 862.280 1424.090 862.340 ;
        RECT 1423.310 814.540 1423.630 814.600 ;
        RECT 1423.115 814.400 1423.630 814.540 ;
        RECT 1423.310 814.340 1423.630 814.400 ;
        RECT 1423.310 787.140 1423.630 787.400 ;
        RECT 1423.400 786.720 1423.540 787.140 ;
        RECT 1423.310 786.460 1423.630 786.720 ;
        RECT 1423.310 724.440 1423.630 724.500 ;
        RECT 1424.230 724.440 1424.550 724.500 ;
        RECT 1423.310 724.300 1424.550 724.440 ;
        RECT 1423.310 724.240 1423.630 724.300 ;
        RECT 1424.230 724.240 1424.550 724.300 ;
        RECT 1423.310 627.880 1423.630 627.940 ;
        RECT 1423.770 627.880 1424.090 627.940 ;
        RECT 1423.310 627.740 1424.090 627.880 ;
        RECT 1423.310 627.680 1423.630 627.740 ;
        RECT 1423.770 627.680 1424.090 627.740 ;
        RECT 1422.865 475.900 1423.155 475.945 ;
        RECT 1423.310 475.900 1423.630 475.960 ;
        RECT 1422.865 475.760 1423.630 475.900 ;
        RECT 1422.865 475.715 1423.155 475.760 ;
        RECT 1423.310 475.700 1423.630 475.760 ;
        RECT 1422.850 427.960 1423.170 428.020 ;
        RECT 1422.655 427.820 1423.170 427.960 ;
        RECT 1422.850 427.760 1423.170 427.820 ;
        RECT 1423.770 255.580 1424.090 255.640 ;
        RECT 1423.400 255.440 1424.090 255.580 ;
        RECT 1423.400 255.300 1423.540 255.440 ;
        RECT 1423.770 255.380 1424.090 255.440 ;
        RECT 1423.310 255.040 1423.630 255.300 ;
        RECT 1422.850 186.560 1423.170 186.620 ;
        RECT 1423.770 186.560 1424.090 186.620 ;
        RECT 1422.850 186.420 1424.090 186.560 ;
        RECT 1422.850 186.360 1423.170 186.420 ;
        RECT 1423.770 186.360 1424.090 186.420 ;
        RECT 1423.325 113.800 1423.615 113.845 ;
        RECT 1424.230 113.800 1424.550 113.860 ;
        RECT 1423.325 113.660 1424.550 113.800 ;
        RECT 1423.325 113.615 1423.615 113.660 ;
        RECT 1424.230 113.600 1424.550 113.660 ;
        RECT 1020.810 49.200 1021.130 49.260 ;
        RECT 1423.325 49.200 1423.615 49.245 ;
        RECT 1020.810 49.060 1423.615 49.200 ;
        RECT 1020.810 49.000 1021.130 49.060 ;
        RECT 1423.325 49.015 1423.615 49.060 ;
      LAYER via ;
        RECT 1424.260 1683.380 1424.520 1683.640 ;
        RECT 1423.340 1635.440 1423.600 1635.700 ;
        RECT 1423.340 1545.680 1423.600 1545.940 ;
        RECT 1423.800 1545.680 1424.060 1545.940 ;
        RECT 1423.800 1490.260 1424.060 1490.520 ;
        RECT 1423.340 1441.980 1423.600 1442.240 ;
        RECT 1423.800 1400.500 1424.060 1400.760 ;
        RECT 1423.800 1352.560 1424.060 1352.820 ;
        RECT 1423.340 1303.940 1423.600 1304.200 ;
        RECT 1423.800 1303.600 1424.060 1303.860 ;
        RECT 1423.800 1159.440 1424.060 1159.700 ;
        RECT 1423.340 1159.100 1423.600 1159.360 ;
        RECT 1423.800 966.320 1424.060 966.580 ;
        RECT 1423.340 965.980 1423.600 966.240 ;
        RECT 1423.800 862.280 1424.060 862.540 ;
        RECT 1423.340 814.340 1423.600 814.600 ;
        RECT 1423.340 787.140 1423.600 787.400 ;
        RECT 1423.340 786.460 1423.600 786.720 ;
        RECT 1423.340 724.240 1423.600 724.500 ;
        RECT 1424.260 724.240 1424.520 724.500 ;
        RECT 1423.340 627.680 1423.600 627.940 ;
        RECT 1423.800 627.680 1424.060 627.940 ;
        RECT 1423.340 475.700 1423.600 475.960 ;
        RECT 1422.880 427.760 1423.140 428.020 ;
        RECT 1423.800 255.380 1424.060 255.640 ;
        RECT 1423.340 255.040 1423.600 255.300 ;
        RECT 1422.880 186.360 1423.140 186.620 ;
        RECT 1423.800 186.360 1424.060 186.620 ;
        RECT 1424.260 113.600 1424.520 113.860 ;
        RECT 1020.840 49.000 1021.100 49.260 ;
      LAYER met2 ;
        RECT 1425.170 1700.410 1425.450 1704.000 ;
        RECT 1424.780 1700.270 1425.450 1700.410 ;
        RECT 1424.780 1686.640 1424.920 1700.270 ;
        RECT 1425.170 1700.000 1425.450 1700.270 ;
        RECT 1424.320 1686.500 1424.920 1686.640 ;
        RECT 1424.320 1683.670 1424.460 1686.500 ;
        RECT 1424.260 1683.350 1424.520 1683.670 ;
        RECT 1423.340 1635.410 1423.600 1635.730 ;
        RECT 1423.400 1545.970 1423.540 1635.410 ;
        RECT 1423.340 1545.650 1423.600 1545.970 ;
        RECT 1423.800 1545.650 1424.060 1545.970 ;
        RECT 1423.860 1490.550 1424.000 1545.650 ;
        RECT 1423.800 1490.230 1424.060 1490.550 ;
        RECT 1423.340 1441.950 1423.600 1442.270 ;
        RECT 1423.400 1425.010 1423.540 1441.950 ;
        RECT 1423.400 1424.870 1424.000 1425.010 ;
        RECT 1423.860 1400.790 1424.000 1424.870 ;
        RECT 1423.800 1400.470 1424.060 1400.790 ;
        RECT 1423.800 1352.530 1424.060 1352.850 ;
        RECT 1423.860 1316.890 1424.000 1352.530 ;
        RECT 1423.400 1316.750 1424.000 1316.890 ;
        RECT 1423.400 1304.230 1423.540 1316.750 ;
        RECT 1423.340 1303.910 1423.600 1304.230 ;
        RECT 1423.800 1303.570 1424.060 1303.890 ;
        RECT 1423.860 1159.730 1424.000 1303.570 ;
        RECT 1423.800 1159.410 1424.060 1159.730 ;
        RECT 1423.340 1159.070 1423.600 1159.390 ;
        RECT 1423.400 1136.010 1423.540 1159.070 ;
        RECT 1423.400 1135.870 1424.460 1136.010 ;
        RECT 1424.320 1124.450 1424.460 1135.870 ;
        RECT 1423.860 1124.310 1424.460 1124.450 ;
        RECT 1423.860 966.610 1424.000 1124.310 ;
        RECT 1423.800 966.290 1424.060 966.610 ;
        RECT 1423.340 965.950 1423.600 966.270 ;
        RECT 1423.400 917.900 1423.540 965.950 ;
        RECT 1423.400 917.760 1424.000 917.900 ;
        RECT 1423.860 862.570 1424.000 917.760 ;
        RECT 1423.800 862.250 1424.060 862.570 ;
        RECT 1423.340 814.310 1423.600 814.630 ;
        RECT 1423.400 787.430 1423.540 814.310 ;
        RECT 1423.340 787.110 1423.600 787.430 ;
        RECT 1423.340 786.430 1423.600 786.750 ;
        RECT 1423.400 724.530 1423.540 786.430 ;
        RECT 1423.340 724.210 1423.600 724.530 ;
        RECT 1424.260 724.210 1424.520 724.530 ;
        RECT 1424.320 699.450 1424.460 724.210 ;
        RECT 1423.860 699.310 1424.460 699.450 ;
        RECT 1423.860 651.850 1424.000 699.310 ;
        RECT 1423.400 651.710 1424.000 651.850 ;
        RECT 1423.400 627.970 1423.540 651.710 ;
        RECT 1423.340 627.650 1423.600 627.970 ;
        RECT 1423.800 627.650 1424.060 627.970 ;
        RECT 1423.860 531.320 1424.000 627.650 ;
        RECT 1423.860 531.180 1424.460 531.320 ;
        RECT 1424.320 483.325 1424.460 531.180 ;
        RECT 1423.330 482.955 1423.610 483.325 ;
        RECT 1424.250 482.955 1424.530 483.325 ;
        RECT 1423.400 475.990 1423.540 482.955 ;
        RECT 1423.340 475.670 1423.600 475.990 ;
        RECT 1422.880 427.730 1423.140 428.050 ;
        RECT 1422.940 404.330 1423.080 427.730 ;
        RECT 1422.940 404.190 1424.000 404.330 ;
        RECT 1423.860 255.670 1424.000 404.190 ;
        RECT 1423.800 255.350 1424.060 255.670 ;
        RECT 1423.340 255.010 1423.600 255.330 ;
        RECT 1423.400 234.330 1423.540 255.010 ;
        RECT 1422.940 234.190 1423.540 234.330 ;
        RECT 1422.940 186.650 1423.080 234.190 ;
        RECT 1422.880 186.330 1423.140 186.650 ;
        RECT 1423.800 186.330 1424.060 186.650 ;
        RECT 1423.860 186.050 1424.000 186.330 ;
        RECT 1423.860 185.910 1424.460 186.050 ;
        RECT 1424.320 113.890 1424.460 185.910 ;
        RECT 1424.260 113.570 1424.520 113.890 ;
        RECT 1020.840 48.970 1021.100 49.290 ;
        RECT 1020.900 3.130 1021.040 48.970 ;
        RECT 1019.520 2.990 1021.040 3.130 ;
        RECT 1019.520 2.400 1019.660 2.990 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
      LAYER via2 ;
        RECT 1423.330 483.000 1423.610 483.280 ;
        RECT 1424.250 483.000 1424.530 483.280 ;
      LAYER met3 ;
        RECT 1423.305 483.290 1423.635 483.305 ;
        RECT 1424.225 483.290 1424.555 483.305 ;
        RECT 1423.305 482.990 1424.555 483.290 ;
        RECT 1423.305 482.975 1423.635 482.990 ;
        RECT 1424.225 482.975 1424.555 482.990 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1020.810 1556.080 1021.130 1556.140 ;
        RECT 1424.690 1556.080 1425.010 1556.140 ;
        RECT 1020.810 1555.940 1425.010 1556.080 ;
        RECT 1020.810 1555.880 1021.130 1555.940 ;
        RECT 1424.690 1555.880 1425.010 1555.940 ;
      LAYER via ;
        RECT 1020.840 1555.880 1021.100 1556.140 ;
        RECT 1424.720 1555.880 1424.980 1556.140 ;
      LAYER met2 ;
        RECT 1426.090 1700.410 1426.370 1704.000 ;
        RECT 1425.240 1700.270 1426.370 1700.410 ;
        RECT 1425.240 1656.210 1425.380 1700.270 ;
        RECT 1426.090 1700.000 1426.370 1700.270 ;
        RECT 1424.780 1656.070 1425.380 1656.210 ;
        RECT 1424.780 1556.170 1424.920 1656.070 ;
        RECT 1020.840 1555.850 1021.100 1556.170 ;
        RECT 1424.720 1555.850 1424.980 1556.170 ;
        RECT 1020.900 3.130 1021.040 1555.850 ;
        RECT 1019.520 2.990 1021.040 3.130 ;
        RECT 1019.520 2.400 1019.660 2.990 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 0.300 ;
=======
      LAYER met1 ;
        RECT 1041.510 1660.120 1041.830 1660.180 ;
        RECT 1431.130 1660.120 1431.450 1660.180 ;
        RECT 1041.510 1659.980 1431.450 1660.120 ;
        RECT 1041.510 1659.920 1041.830 1659.980 ;
        RECT 1431.130 1659.920 1431.450 1659.980 ;
        RECT 1037.370 2.960 1037.690 3.020 ;
        RECT 1041.510 2.960 1041.830 3.020 ;
        RECT 1037.370 2.820 1041.830 2.960 ;
        RECT 1037.370 2.760 1037.690 2.820 ;
        RECT 1041.510 2.760 1041.830 2.820 ;
      LAYER via ;
        RECT 1041.540 1659.920 1041.800 1660.180 ;
        RECT 1431.160 1659.920 1431.420 1660.180 ;
        RECT 1037.400 2.760 1037.660 3.020 ;
        RECT 1041.540 2.760 1041.800 3.020 ;
      LAYER met2 ;
        RECT 1431.150 1700.000 1431.430 1704.000 ;
        RECT 1431.220 1660.210 1431.360 1700.000 ;
        RECT 1041.540 1659.890 1041.800 1660.210 ;
        RECT 1431.160 1659.890 1431.420 1660.210 ;
        RECT 1041.600 3.050 1041.740 1659.890 ;
        RECT 1037.400 2.730 1037.660 3.050 ;
        RECT 1041.540 2.730 1041.800 3.050 ;
        RECT 1037.460 2.400 1037.600 2.730 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1055.310 1646.180 1055.630 1646.240 ;
        RECT 1436.190 1646.180 1436.510 1646.240 ;
        RECT 1055.310 1646.040 1436.510 1646.180 ;
        RECT 1055.310 1645.980 1055.630 1646.040 ;
        RECT 1436.190 1645.980 1436.510 1646.040 ;
      LAYER via ;
        RECT 1055.340 1645.980 1055.600 1646.240 ;
        RECT 1436.220 1645.980 1436.480 1646.240 ;
      LAYER met2 ;
        RECT 1435.750 1700.410 1436.030 1704.000 ;
        RECT 1435.750 1700.270 1436.420 1700.410 ;
        RECT 1435.750 1700.000 1436.030 1700.270 ;
        RECT 1436.280 1646.270 1436.420 1700.270 ;
        RECT 1055.340 1645.950 1055.600 1646.270 ;
        RECT 1436.220 1645.950 1436.480 1646.270 ;
        RECT 1055.400 2.400 1055.540 1645.950 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1435.270 1678.140 1435.590 1678.200 ;
        RECT 1439.410 1678.140 1439.730 1678.200 ;
        RECT 1435.270 1678.000 1439.730 1678.140 ;
        RECT 1435.270 1677.940 1435.590 1678.000 ;
        RECT 1439.410 1677.940 1439.730 1678.000 ;
        RECT 1076.010 1653.320 1076.330 1653.380 ;
        RECT 1435.270 1653.320 1435.590 1653.380 ;
        RECT 1076.010 1653.180 1435.590 1653.320 ;
        RECT 1076.010 1653.120 1076.330 1653.180 ;
        RECT 1435.270 1653.120 1435.590 1653.180 ;
        RECT 1073.250 2.960 1073.570 3.020 ;
        RECT 1076.010 2.960 1076.330 3.020 ;
        RECT 1073.250 2.820 1076.330 2.960 ;
        RECT 1073.250 2.760 1073.570 2.820 ;
        RECT 1076.010 2.760 1076.330 2.820 ;
      LAYER via ;
        RECT 1435.300 1677.940 1435.560 1678.200 ;
        RECT 1439.440 1677.940 1439.700 1678.200 ;
        RECT 1076.040 1653.120 1076.300 1653.380 ;
        RECT 1435.300 1653.120 1435.560 1653.380 ;
        RECT 1073.280 2.760 1073.540 3.020 ;
        RECT 1076.040 2.760 1076.300 3.020 ;
      LAYER met2 ;
        RECT 1440.810 1700.410 1441.090 1704.000 ;
        RECT 1439.500 1700.270 1441.090 1700.410 ;
        RECT 1439.500 1678.230 1439.640 1700.270 ;
        RECT 1440.810 1700.000 1441.090 1700.270 ;
        RECT 1435.300 1677.910 1435.560 1678.230 ;
        RECT 1439.440 1677.910 1439.700 1678.230 ;
        RECT 1435.360 1653.410 1435.500 1677.910 ;
        RECT 1076.040 1653.090 1076.300 1653.410 ;
        RECT 1435.300 1653.090 1435.560 1653.410 ;
        RECT 1076.100 3.050 1076.240 1653.090 ;
        RECT 1073.280 2.730 1073.540 3.050 ;
        RECT 1076.040 2.730 1076.300 3.050 ;
        RECT 1073.340 2.400 1073.480 2.730 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1096.250 1673.720 1096.570 1673.780 ;
        RECT 1445.390 1673.720 1445.710 1673.780 ;
        RECT 1096.250 1673.580 1445.710 1673.720 ;
        RECT 1096.250 1673.520 1096.570 1673.580 ;
        RECT 1445.390 1673.520 1445.710 1673.580 ;
        RECT 1090.730 2.960 1091.050 3.020 ;
        RECT 1096.250 2.960 1096.570 3.020 ;
        RECT 1090.730 2.820 1096.570 2.960 ;
        RECT 1090.730 2.760 1091.050 2.820 ;
        RECT 1096.250 2.760 1096.570 2.820 ;
      LAYER via ;
        RECT 1096.280 1673.520 1096.540 1673.780 ;
        RECT 1445.420 1673.520 1445.680 1673.780 ;
        RECT 1090.760 2.760 1091.020 3.020 ;
        RECT 1096.280 2.760 1096.540 3.020 ;
      LAYER met2 ;
        RECT 1445.410 1700.000 1445.690 1704.000 ;
        RECT 1445.480 1673.810 1445.620 1700.000 ;
        RECT 1096.280 1673.490 1096.540 1673.810 ;
        RECT 1445.420 1673.490 1445.680 1673.810 ;
        RECT 1096.340 3.050 1096.480 1673.490 ;
        RECT 1090.760 2.730 1091.020 3.050 ;
        RECT 1096.280 2.730 1096.540 3.050 ;
        RECT 1090.820 2.400 1090.960 2.730 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 0.300 ;
=======
      LAYER li1 ;
        RECT 1450.065 1607.605 1450.235 1635.315 ;
        RECT 1450.065 1400.885 1450.235 1562.895 ;
        RECT 1450.065 1158.805 1450.235 1200.115 ;
        RECT 1450.065 1062.585 1450.235 1128.375 ;
        RECT 1450.525 869.805 1450.695 917.575 ;
        RECT 1450.065 662.405 1450.235 676.855 ;
        RECT 1450.065 403.665 1450.235 434.435 ;
        RECT 1450.065 96.645 1450.235 144.755 ;
        RECT 1450.065 42.245 1450.235 48.195 ;
      LAYER mcon ;
        RECT 1450.065 1635.145 1450.235 1635.315 ;
        RECT 1450.065 1562.725 1450.235 1562.895 ;
        RECT 1450.065 1199.945 1450.235 1200.115 ;
        RECT 1450.065 1128.205 1450.235 1128.375 ;
        RECT 1450.525 917.405 1450.695 917.575 ;
        RECT 1450.065 676.685 1450.235 676.855 ;
        RECT 1450.065 434.265 1450.235 434.435 ;
        RECT 1450.065 144.585 1450.235 144.755 ;
        RECT 1450.065 48.025 1450.235 48.195 ;
      LAYER met1 ;
        RECT 1449.070 1656.380 1449.390 1656.440 ;
        RECT 1449.990 1656.380 1450.310 1656.440 ;
        RECT 1449.070 1656.240 1450.310 1656.380 ;
        RECT 1449.070 1656.180 1449.390 1656.240 ;
        RECT 1449.990 1656.180 1450.310 1656.240 ;
        RECT 1449.990 1635.300 1450.310 1635.360 ;
        RECT 1449.795 1635.160 1450.310 1635.300 ;
        RECT 1449.990 1635.100 1450.310 1635.160 ;
        RECT 1450.005 1607.760 1450.295 1607.805 ;
        RECT 1451.830 1607.760 1452.150 1607.820 ;
        RECT 1450.005 1607.620 1452.150 1607.760 ;
        RECT 1450.005 1607.575 1450.295 1607.620 ;
        RECT 1451.830 1607.560 1452.150 1607.620 ;
        RECT 1450.005 1562.880 1450.295 1562.925 ;
        RECT 1451.830 1562.880 1452.150 1562.940 ;
        RECT 1450.005 1562.740 1452.150 1562.880 ;
        RECT 1450.005 1562.695 1450.295 1562.740 ;
        RECT 1451.830 1562.680 1452.150 1562.740 ;
        RECT 1449.990 1401.040 1450.310 1401.100 ;
        RECT 1449.795 1400.900 1450.310 1401.040 ;
        RECT 1449.990 1400.840 1450.310 1400.900 ;
        RECT 1449.070 1297.340 1449.390 1297.400 ;
        RECT 1449.990 1297.340 1450.310 1297.400 ;
        RECT 1449.070 1297.200 1450.310 1297.340 ;
        RECT 1449.070 1297.140 1449.390 1297.200 ;
        RECT 1449.990 1297.140 1450.310 1297.200 ;
        RECT 1449.990 1249.060 1450.310 1249.120 ;
        RECT 1450.450 1249.060 1450.770 1249.120 ;
        RECT 1449.990 1248.920 1450.770 1249.060 ;
        RECT 1449.990 1248.860 1450.310 1248.920 ;
        RECT 1450.450 1248.860 1450.770 1248.920 ;
        RECT 1449.990 1200.100 1450.310 1200.160 ;
        RECT 1449.795 1199.960 1450.310 1200.100 ;
        RECT 1449.990 1199.900 1450.310 1199.960 ;
        RECT 1449.990 1158.960 1450.310 1159.020 ;
        RECT 1449.795 1158.820 1450.310 1158.960 ;
        RECT 1449.990 1158.760 1450.310 1158.820 ;
        RECT 1449.990 1128.360 1450.310 1128.420 ;
        RECT 1449.795 1128.220 1450.310 1128.360 ;
        RECT 1449.990 1128.160 1450.310 1128.220 ;
        RECT 1450.005 1062.740 1450.295 1062.785 ;
        RECT 1450.450 1062.740 1450.770 1062.800 ;
        RECT 1450.005 1062.600 1450.770 1062.740 ;
        RECT 1450.005 1062.555 1450.295 1062.600 ;
        RECT 1450.450 1062.540 1450.770 1062.600 ;
        RECT 1449.070 1014.460 1449.390 1014.520 ;
        RECT 1449.990 1014.460 1450.310 1014.520 ;
        RECT 1449.070 1014.320 1450.310 1014.460 ;
        RECT 1449.070 1014.260 1449.390 1014.320 ;
        RECT 1449.990 1014.260 1450.310 1014.320 ;
        RECT 1449.070 917.900 1449.390 917.960 ;
        RECT 1449.990 917.900 1450.310 917.960 ;
        RECT 1449.070 917.760 1450.310 917.900 ;
        RECT 1449.070 917.700 1449.390 917.760 ;
        RECT 1449.990 917.700 1450.310 917.760 ;
        RECT 1450.450 917.560 1450.770 917.620 ;
        RECT 1450.255 917.420 1450.770 917.560 ;
        RECT 1450.450 917.360 1450.770 917.420 ;
        RECT 1450.450 869.960 1450.770 870.020 ;
        RECT 1450.255 869.820 1450.770 869.960 ;
        RECT 1450.450 869.760 1450.770 869.820 ;
        RECT 1449.070 772.720 1449.390 772.780 ;
        RECT 1450.450 772.720 1450.770 772.780 ;
        RECT 1449.070 772.580 1450.770 772.720 ;
        RECT 1449.070 772.520 1449.390 772.580 ;
        RECT 1450.450 772.520 1450.770 772.580 ;
        RECT 1449.990 676.840 1450.310 676.900 ;
        RECT 1449.795 676.700 1450.310 676.840 ;
        RECT 1449.990 676.640 1450.310 676.700 ;
        RECT 1449.990 662.560 1450.310 662.620 ;
        RECT 1449.795 662.420 1450.310 662.560 ;
        RECT 1449.990 662.360 1450.310 662.420 ;
        RECT 1449.990 651.140 1450.310 651.400 ;
        RECT 1450.080 650.720 1450.220 651.140 ;
        RECT 1449.990 650.460 1450.310 650.720 ;
        RECT 1449.990 593.680 1450.310 593.940 ;
        RECT 1450.080 593.260 1450.220 593.680 ;
        RECT 1449.990 593.000 1450.310 593.260 ;
        RECT 1449.990 531.320 1450.310 531.380 ;
        RECT 1450.450 531.320 1450.770 531.380 ;
        RECT 1449.990 531.180 1450.770 531.320 ;
        RECT 1449.990 531.120 1450.310 531.180 ;
        RECT 1450.450 531.120 1450.770 531.180 ;
        RECT 1449.070 524.180 1449.390 524.240 ;
        RECT 1450.450 524.180 1450.770 524.240 ;
        RECT 1449.070 524.040 1450.770 524.180 ;
        RECT 1449.070 523.980 1449.390 524.040 ;
        RECT 1450.450 523.980 1450.770 524.040 ;
        RECT 1449.990 434.420 1450.310 434.480 ;
        RECT 1449.795 434.280 1450.310 434.420 ;
        RECT 1449.990 434.220 1450.310 434.280 ;
        RECT 1450.005 403.820 1450.295 403.865 ;
        RECT 1450.450 403.820 1450.770 403.880 ;
        RECT 1450.005 403.680 1450.770 403.820 ;
        RECT 1450.005 403.635 1450.295 403.680 ;
        RECT 1450.450 403.620 1450.770 403.680 ;
        RECT 1449.070 310.660 1449.390 310.720 ;
        RECT 1449.990 310.660 1450.310 310.720 ;
        RECT 1449.070 310.520 1450.310 310.660 ;
        RECT 1449.070 310.460 1449.390 310.520 ;
        RECT 1449.990 310.460 1450.310 310.520 ;
        RECT 1449.070 295.020 1449.390 295.080 ;
        RECT 1449.990 295.020 1450.310 295.080 ;
        RECT 1449.070 294.880 1450.310 295.020 ;
        RECT 1449.070 294.820 1449.390 294.880 ;
        RECT 1449.990 294.820 1450.310 294.880 ;
        RECT 1449.070 241.640 1449.390 241.700 ;
        RECT 1449.990 241.640 1450.310 241.700 ;
        RECT 1449.070 241.500 1450.310 241.640 ;
        RECT 1449.070 241.440 1449.390 241.500 ;
        RECT 1449.990 241.440 1450.310 241.500 ;
        RECT 1449.990 144.740 1450.310 144.800 ;
        RECT 1449.795 144.600 1450.310 144.740 ;
        RECT 1449.990 144.540 1450.310 144.600 ;
        RECT 1450.005 96.800 1450.295 96.845 ;
        RECT 1450.450 96.800 1450.770 96.860 ;
        RECT 1450.005 96.660 1450.770 96.800 ;
        RECT 1450.005 96.615 1450.295 96.660 ;
        RECT 1450.450 96.600 1450.770 96.660 ;
        RECT 1450.450 62.460 1450.770 62.520 ;
        RECT 1450.080 62.320 1450.770 62.460 ;
        RECT 1450.080 62.180 1450.220 62.320 ;
        RECT 1450.450 62.260 1450.770 62.320 ;
        RECT 1449.990 61.920 1450.310 62.180 ;
        RECT 1449.990 48.180 1450.310 48.240 ;
        RECT 1449.795 48.040 1450.310 48.180 ;
        RECT 1449.990 47.980 1450.310 48.040 ;
        RECT 1108.670 42.400 1108.990 42.460 ;
        RECT 1450.005 42.400 1450.295 42.445 ;
        RECT 1108.670 42.260 1450.295 42.400 ;
        RECT 1108.670 42.200 1108.990 42.260 ;
        RECT 1450.005 42.215 1450.295 42.260 ;
      LAYER via ;
        RECT 1449.100 1656.180 1449.360 1656.440 ;
        RECT 1450.020 1656.180 1450.280 1656.440 ;
        RECT 1450.020 1635.100 1450.280 1635.360 ;
        RECT 1451.860 1607.560 1452.120 1607.820 ;
        RECT 1451.860 1562.680 1452.120 1562.940 ;
        RECT 1450.020 1400.840 1450.280 1401.100 ;
        RECT 1449.100 1297.140 1449.360 1297.400 ;
        RECT 1450.020 1297.140 1450.280 1297.400 ;
        RECT 1450.020 1248.860 1450.280 1249.120 ;
        RECT 1450.480 1248.860 1450.740 1249.120 ;
        RECT 1450.020 1199.900 1450.280 1200.160 ;
        RECT 1450.020 1158.760 1450.280 1159.020 ;
        RECT 1450.020 1128.160 1450.280 1128.420 ;
        RECT 1450.480 1062.540 1450.740 1062.800 ;
        RECT 1449.100 1014.260 1449.360 1014.520 ;
        RECT 1450.020 1014.260 1450.280 1014.520 ;
        RECT 1449.100 917.700 1449.360 917.960 ;
        RECT 1450.020 917.700 1450.280 917.960 ;
        RECT 1450.480 917.360 1450.740 917.620 ;
        RECT 1450.480 869.760 1450.740 870.020 ;
        RECT 1449.100 772.520 1449.360 772.780 ;
        RECT 1450.480 772.520 1450.740 772.780 ;
        RECT 1450.020 676.640 1450.280 676.900 ;
        RECT 1450.020 662.360 1450.280 662.620 ;
        RECT 1450.020 651.140 1450.280 651.400 ;
        RECT 1450.020 650.460 1450.280 650.720 ;
        RECT 1450.020 593.680 1450.280 593.940 ;
        RECT 1450.020 593.000 1450.280 593.260 ;
        RECT 1450.020 531.120 1450.280 531.380 ;
        RECT 1450.480 531.120 1450.740 531.380 ;
        RECT 1449.100 523.980 1449.360 524.240 ;
        RECT 1450.480 523.980 1450.740 524.240 ;
        RECT 1450.020 434.220 1450.280 434.480 ;
        RECT 1450.480 403.620 1450.740 403.880 ;
        RECT 1449.100 310.460 1449.360 310.720 ;
        RECT 1450.020 310.460 1450.280 310.720 ;
        RECT 1449.100 294.820 1449.360 295.080 ;
        RECT 1450.020 294.820 1450.280 295.080 ;
        RECT 1449.100 241.440 1449.360 241.700 ;
        RECT 1450.020 241.440 1450.280 241.700 ;
        RECT 1450.020 144.540 1450.280 144.800 ;
        RECT 1450.480 96.600 1450.740 96.860 ;
        RECT 1450.480 62.260 1450.740 62.520 ;
        RECT 1450.020 61.920 1450.280 62.180 ;
        RECT 1450.020 47.980 1450.280 48.240 ;
        RECT 1108.700 42.200 1108.960 42.460 ;
      LAYER met2 ;
        RECT 1449.090 1700.000 1449.370 1704.000 ;
        RECT 1449.160 1656.470 1449.300 1700.000 ;
        RECT 1449.100 1656.150 1449.360 1656.470 ;
        RECT 1450.020 1656.150 1450.280 1656.470 ;
        RECT 1450.080 1635.390 1450.220 1656.150 ;
        RECT 1450.020 1635.070 1450.280 1635.390 ;
        RECT 1451.860 1607.530 1452.120 1607.850 ;
        RECT 1451.920 1562.970 1452.060 1607.530 ;
        RECT 1451.860 1562.650 1452.120 1562.970 ;
        RECT 1450.020 1400.810 1450.280 1401.130 ;
        RECT 1450.080 1393.845 1450.220 1400.810 ;
        RECT 1450.010 1393.475 1450.290 1393.845 ;
        RECT 1449.090 1345.195 1449.370 1345.565 ;
        RECT 1449.160 1297.430 1449.300 1345.195 ;
        RECT 1449.100 1297.110 1449.360 1297.430 ;
        RECT 1450.020 1297.285 1450.280 1297.430 ;
        RECT 1450.010 1296.915 1450.290 1297.285 ;
        RECT 1450.470 1296.235 1450.750 1296.605 ;
        RECT 1450.540 1249.150 1450.680 1296.235 ;
        RECT 1450.020 1248.830 1450.280 1249.150 ;
        RECT 1450.480 1248.830 1450.740 1249.150 ;
        RECT 1450.080 1200.190 1450.220 1248.830 ;
        RECT 1450.020 1199.870 1450.280 1200.190 ;
        RECT 1450.020 1158.730 1450.280 1159.050 ;
        RECT 1450.080 1128.450 1450.220 1158.730 ;
        RECT 1450.020 1128.130 1450.280 1128.450 ;
        RECT 1450.480 1062.685 1450.740 1062.830 ;
        RECT 1449.090 1062.315 1449.370 1062.685 ;
        RECT 1450.470 1062.315 1450.750 1062.685 ;
        RECT 1449.160 1014.550 1449.300 1062.315 ;
        RECT 1449.100 1014.230 1449.360 1014.550 ;
        RECT 1450.020 1014.405 1450.280 1014.550 ;
        RECT 1450.010 1014.035 1450.290 1014.405 ;
        RECT 1449.090 965.755 1449.370 966.125 ;
        RECT 1449.160 917.990 1449.300 965.755 ;
        RECT 1450.080 917.990 1450.220 918.145 ;
        RECT 1449.100 917.670 1449.360 917.990 ;
        RECT 1450.020 917.730 1450.280 917.990 ;
        RECT 1450.020 917.670 1450.680 917.730 ;
        RECT 1450.080 917.650 1450.680 917.670 ;
        RECT 1450.080 917.590 1450.740 917.650 ;
        RECT 1450.480 917.330 1450.740 917.590 ;
        RECT 1450.480 869.730 1450.740 870.050 ;
        RECT 1450.540 869.565 1450.680 869.730 ;
        RECT 1449.090 869.195 1449.370 869.565 ;
        RECT 1450.470 869.195 1450.750 869.565 ;
        RECT 1449.160 821.285 1449.300 869.195 ;
        RECT 1449.090 820.915 1449.370 821.285 ;
        RECT 1450.010 820.915 1450.290 821.285 ;
        RECT 1450.080 772.890 1450.220 820.915 ;
        RECT 1450.080 772.810 1450.680 772.890 ;
        RECT 1449.100 772.490 1449.360 772.810 ;
        RECT 1450.080 772.750 1450.740 772.810 ;
        RECT 1450.480 772.490 1450.740 772.750 ;
        RECT 1449.160 724.725 1449.300 772.490 ;
        RECT 1450.540 772.335 1450.680 772.490 ;
        RECT 1449.090 724.355 1449.370 724.725 ;
        RECT 1450.010 724.355 1450.290 724.725 ;
        RECT 1450.080 676.930 1450.220 724.355 ;
        RECT 1450.020 676.610 1450.280 676.930 ;
        RECT 1450.020 662.330 1450.280 662.650 ;
        RECT 1450.080 651.430 1450.220 662.330 ;
        RECT 1450.020 651.110 1450.280 651.430 ;
        RECT 1450.020 650.430 1450.280 650.750 ;
        RECT 1450.080 593.970 1450.220 650.430 ;
        RECT 1450.020 593.650 1450.280 593.970 ;
        RECT 1450.020 592.970 1450.280 593.290 ;
        RECT 1450.080 531.410 1450.220 592.970 ;
        RECT 1450.020 531.090 1450.280 531.410 ;
        RECT 1450.480 531.090 1450.740 531.410 ;
        RECT 1450.540 524.270 1450.680 531.090 ;
        RECT 1449.100 523.950 1449.360 524.270 ;
        RECT 1450.480 523.950 1450.740 524.270 ;
        RECT 1449.160 435.045 1449.300 523.950 ;
        RECT 1449.090 434.675 1449.370 435.045 ;
        RECT 1450.010 434.675 1450.290 435.045 ;
        RECT 1450.080 434.510 1450.220 434.675 ;
        RECT 1450.020 434.190 1450.280 434.510 ;
        RECT 1450.480 403.590 1450.740 403.910 ;
        RECT 1450.540 358.885 1450.680 403.590 ;
        RECT 1449.090 358.515 1449.370 358.885 ;
        RECT 1450.470 358.515 1450.750 358.885 ;
        RECT 1449.160 310.750 1449.300 358.515 ;
        RECT 1449.100 310.430 1449.360 310.750 ;
        RECT 1450.020 310.430 1450.280 310.750 ;
        RECT 1450.080 295.110 1450.220 310.430 ;
        RECT 1449.100 294.790 1449.360 295.110 ;
        RECT 1450.020 294.790 1450.280 295.110 ;
        RECT 1449.160 241.730 1449.300 294.790 ;
        RECT 1449.100 241.410 1449.360 241.730 ;
        RECT 1450.020 241.410 1450.280 241.730 ;
        RECT 1450.080 217.330 1450.220 241.410 ;
        RECT 1450.080 217.190 1450.680 217.330 ;
        RECT 1450.540 145.250 1450.680 217.190 ;
        RECT 1450.080 145.110 1450.680 145.250 ;
        RECT 1450.080 144.830 1450.220 145.110 ;
        RECT 1450.020 144.510 1450.280 144.830 ;
        RECT 1450.480 96.570 1450.740 96.890 ;
        RECT 1450.540 62.550 1450.680 96.570 ;
        RECT 1450.480 62.230 1450.740 62.550 ;
        RECT 1450.020 61.890 1450.280 62.210 ;
        RECT 1450.080 48.270 1450.220 61.890 ;
        RECT 1450.020 47.950 1450.280 48.270 ;
        RECT 1108.700 42.170 1108.960 42.490 ;
        RECT 1108.760 2.400 1108.900 42.170 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
      LAYER via2 ;
        RECT 1450.010 1393.520 1450.290 1393.800 ;
        RECT 1449.090 1345.240 1449.370 1345.520 ;
        RECT 1450.010 1296.960 1450.290 1297.240 ;
        RECT 1450.470 1296.280 1450.750 1296.560 ;
        RECT 1449.090 1062.360 1449.370 1062.640 ;
        RECT 1450.470 1062.360 1450.750 1062.640 ;
        RECT 1450.010 1014.080 1450.290 1014.360 ;
        RECT 1449.090 965.800 1449.370 966.080 ;
        RECT 1449.090 869.240 1449.370 869.520 ;
        RECT 1450.470 869.240 1450.750 869.520 ;
        RECT 1449.090 820.960 1449.370 821.240 ;
        RECT 1450.010 820.960 1450.290 821.240 ;
        RECT 1449.090 724.400 1449.370 724.680 ;
        RECT 1450.010 724.400 1450.290 724.680 ;
        RECT 1449.090 434.720 1449.370 435.000 ;
        RECT 1450.010 434.720 1450.290 435.000 ;
        RECT 1449.090 358.560 1449.370 358.840 ;
        RECT 1450.470 358.560 1450.750 358.840 ;
      LAYER met3 ;
        RECT 1449.985 1393.810 1450.315 1393.825 ;
        RECT 1451.110 1393.810 1451.490 1393.820 ;
        RECT 1449.985 1393.510 1451.490 1393.810 ;
        RECT 1449.985 1393.495 1450.315 1393.510 ;
        RECT 1451.110 1393.500 1451.490 1393.510 ;
        RECT 1451.110 1345.900 1451.490 1346.220 ;
        RECT 1449.065 1345.530 1449.395 1345.545 ;
        RECT 1451.150 1345.530 1451.450 1345.900 ;
        RECT 1449.065 1345.230 1451.450 1345.530 ;
        RECT 1449.065 1345.215 1449.395 1345.230 ;
        RECT 1449.985 1297.250 1450.315 1297.265 ;
        RECT 1449.985 1296.935 1450.530 1297.250 ;
        RECT 1450.230 1296.585 1450.530 1296.935 ;
        RECT 1450.230 1296.270 1450.775 1296.585 ;
        RECT 1450.445 1296.255 1450.775 1296.270 ;
        RECT 1449.065 1062.650 1449.395 1062.665 ;
        RECT 1450.445 1062.650 1450.775 1062.665 ;
        RECT 1449.065 1062.350 1450.775 1062.650 ;
        RECT 1449.065 1062.335 1449.395 1062.350 ;
        RECT 1450.445 1062.335 1450.775 1062.350 ;
        RECT 1449.985 1014.380 1450.315 1014.385 ;
        RECT 1449.985 1014.370 1450.570 1014.380 ;
        RECT 1449.760 1014.070 1450.570 1014.370 ;
        RECT 1449.985 1014.060 1450.570 1014.070 ;
        RECT 1449.985 1014.055 1450.315 1014.060 ;
        RECT 1450.190 967.450 1450.570 967.460 ;
        RECT 1450.190 967.150 1451.450 967.450 ;
        RECT 1450.190 967.140 1450.570 967.150 ;
        RECT 1449.065 966.090 1449.395 966.105 ;
        RECT 1451.150 966.090 1451.450 967.150 ;
        RECT 1449.065 965.790 1451.450 966.090 ;
        RECT 1449.065 965.775 1449.395 965.790 ;
        RECT 1449.065 869.530 1449.395 869.545 ;
        RECT 1450.445 869.530 1450.775 869.545 ;
        RECT 1449.065 869.230 1450.775 869.530 ;
        RECT 1449.065 869.215 1449.395 869.230 ;
        RECT 1450.445 869.215 1450.775 869.230 ;
        RECT 1449.065 821.250 1449.395 821.265 ;
        RECT 1449.985 821.250 1450.315 821.265 ;
        RECT 1449.065 820.950 1450.315 821.250 ;
        RECT 1449.065 820.935 1449.395 820.950 ;
        RECT 1449.985 820.935 1450.315 820.950 ;
        RECT 1449.065 724.690 1449.395 724.705 ;
        RECT 1449.985 724.690 1450.315 724.705 ;
        RECT 1449.065 724.390 1450.315 724.690 ;
        RECT 1449.065 724.375 1449.395 724.390 ;
        RECT 1449.985 724.375 1450.315 724.390 ;
        RECT 1449.065 435.010 1449.395 435.025 ;
        RECT 1449.985 435.010 1450.315 435.025 ;
        RECT 1449.065 434.710 1450.315 435.010 ;
        RECT 1449.065 434.695 1449.395 434.710 ;
        RECT 1449.985 434.695 1450.315 434.710 ;
        RECT 1449.065 358.850 1449.395 358.865 ;
        RECT 1450.445 358.850 1450.775 358.865 ;
        RECT 1449.065 358.550 1450.775 358.850 ;
        RECT 1449.065 358.535 1449.395 358.550 ;
        RECT 1450.445 358.535 1450.775 358.550 ;
      LAYER via3 ;
        RECT 1451.140 1393.500 1451.460 1393.820 ;
        RECT 1451.140 1345.900 1451.460 1346.220 ;
        RECT 1450.220 1014.060 1450.540 1014.380 ;
        RECT 1450.220 967.140 1450.540 967.460 ;
      LAYER met4 ;
        RECT 1451.135 1393.495 1451.465 1393.825 ;
        RECT 1451.150 1346.225 1451.450 1393.495 ;
        RECT 1451.135 1345.895 1451.465 1346.225 ;
        RECT 1450.215 1014.055 1450.545 1014.385 ;
        RECT 1450.230 967.465 1450.530 1014.055 ;
        RECT 1450.215 967.135 1450.545 967.465 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1108.670 42.740 1108.990 42.800 ;
        RECT 1449.530 42.740 1449.850 42.800 ;
        RECT 1108.670 42.600 1449.850 42.740 ;
        RECT 1108.670 42.540 1108.990 42.600 ;
        RECT 1449.530 42.540 1449.850 42.600 ;
      LAYER via ;
        RECT 1108.700 42.540 1108.960 42.800 ;
        RECT 1449.560 42.540 1449.820 42.800 ;
      LAYER met2 ;
        RECT 1450.470 1700.410 1450.750 1704.000 ;
        RECT 1449.620 1700.270 1450.750 1700.410 ;
        RECT 1449.620 42.830 1449.760 1700.270 ;
        RECT 1450.470 1700.000 1450.750 1700.270 ;
        RECT 1108.700 42.510 1108.960 42.830 ;
        RECT 1449.560 42.510 1449.820 42.830 ;
        RECT 1108.760 2.400 1108.900 42.510 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 0.300 ;
=======
      LAYER li1 ;
        RECT 1452.365 1545.045 1452.535 1635.315 ;
        RECT 1451.905 965.005 1452.075 1007.335 ;
        RECT 1451.905 917.745 1452.075 931.855 ;
        RECT 1451.905 379.525 1452.075 434.435 ;
        RECT 1451.905 41.905 1452.075 48.195 ;
      LAYER mcon ;
        RECT 1452.365 1635.145 1452.535 1635.315 ;
        RECT 1451.905 1007.165 1452.075 1007.335 ;
        RECT 1451.905 931.685 1452.075 931.855 ;
        RECT 1451.905 434.265 1452.075 434.435 ;
        RECT 1451.905 48.025 1452.075 48.195 ;
      LAYER met1 ;
        RECT 1451.830 1635.300 1452.150 1635.360 ;
        RECT 1452.305 1635.300 1452.595 1635.345 ;
        RECT 1451.830 1635.160 1452.595 1635.300 ;
        RECT 1451.830 1635.100 1452.150 1635.160 ;
        RECT 1452.305 1635.115 1452.595 1635.160 ;
        RECT 1452.305 1545.200 1452.595 1545.245 ;
        RECT 1452.750 1545.200 1453.070 1545.260 ;
        RECT 1452.305 1545.060 1453.070 1545.200 ;
        RECT 1452.305 1545.015 1452.595 1545.060 ;
        RECT 1452.750 1545.000 1453.070 1545.060 ;
        RECT 1452.750 1490.260 1453.070 1490.520 ;
        RECT 1452.840 1489.840 1452.980 1490.260 ;
        RECT 1452.750 1489.580 1453.070 1489.840 ;
        RECT 1451.830 1393.900 1452.150 1393.960 ;
        RECT 1452.750 1393.900 1453.070 1393.960 ;
        RECT 1451.830 1393.760 1453.070 1393.900 ;
        RECT 1451.830 1393.700 1452.150 1393.760 ;
        RECT 1452.750 1393.700 1453.070 1393.760 ;
        RECT 1451.830 1345.620 1452.150 1345.680 ;
        RECT 1453.210 1345.620 1453.530 1345.680 ;
        RECT 1451.830 1345.480 1453.530 1345.620 ;
        RECT 1451.830 1345.420 1452.150 1345.480 ;
        RECT 1453.210 1345.420 1453.530 1345.480 ;
        RECT 1451.830 1297.340 1452.150 1297.400 ;
        RECT 1452.750 1297.340 1453.070 1297.400 ;
        RECT 1451.830 1297.200 1453.070 1297.340 ;
        RECT 1451.830 1297.140 1452.150 1297.200 ;
        RECT 1452.750 1297.140 1453.070 1297.200 ;
        RECT 1451.830 1269.600 1452.150 1269.860 ;
        RECT 1451.920 1269.460 1452.060 1269.600 ;
        RECT 1452.290 1269.460 1452.610 1269.520 ;
        RECT 1451.920 1269.320 1452.610 1269.460 ;
        RECT 1452.290 1269.260 1452.610 1269.320 ;
        RECT 1451.830 1152.500 1452.150 1152.560 ;
        RECT 1452.750 1152.500 1453.070 1152.560 ;
        RECT 1451.830 1152.360 1453.070 1152.500 ;
        RECT 1451.830 1152.300 1452.150 1152.360 ;
        RECT 1452.750 1152.300 1453.070 1152.360 ;
        RECT 1451.830 1007.320 1452.150 1007.380 ;
        RECT 1451.635 1007.180 1452.150 1007.320 ;
        RECT 1451.830 1007.120 1452.150 1007.180 ;
        RECT 1451.830 965.160 1452.150 965.220 ;
        RECT 1451.635 965.020 1452.150 965.160 ;
        RECT 1451.830 964.960 1452.150 965.020 ;
        RECT 1451.830 931.840 1452.150 931.900 ;
        RECT 1451.635 931.700 1452.150 931.840 ;
        RECT 1451.830 931.640 1452.150 931.700 ;
        RECT 1451.830 917.900 1452.150 917.960 ;
        RECT 1451.635 917.760 1452.150 917.900 ;
        RECT 1451.830 917.700 1452.150 917.760 ;
        RECT 1451.830 910.760 1452.150 910.820 ;
        RECT 1453.210 910.760 1453.530 910.820 ;
        RECT 1451.830 910.620 1453.530 910.760 ;
        RECT 1451.830 910.560 1452.150 910.620 ;
        RECT 1453.210 910.560 1453.530 910.620 ;
        RECT 1452.290 820.800 1452.610 821.060 ;
        RECT 1452.380 820.380 1452.520 820.800 ;
        RECT 1452.290 820.120 1452.610 820.380 ;
        RECT 1452.290 765.920 1452.610 765.980 ;
        RECT 1453.210 765.920 1453.530 765.980 ;
        RECT 1452.290 765.780 1453.530 765.920 ;
        RECT 1452.290 765.720 1452.610 765.780 ;
        RECT 1453.210 765.720 1453.530 765.780 ;
        RECT 1451.830 593.340 1452.150 593.600 ;
        RECT 1451.920 593.200 1452.060 593.340 ;
        RECT 1452.290 593.200 1452.610 593.260 ;
        RECT 1451.920 593.060 1452.610 593.200 ;
        RECT 1452.290 593.000 1452.610 593.060 ;
        RECT 1452.290 449.040 1452.610 449.100 ;
        RECT 1451.920 448.900 1452.610 449.040 ;
        RECT 1451.920 448.420 1452.060 448.900 ;
        RECT 1452.290 448.840 1452.610 448.900 ;
        RECT 1451.830 448.160 1452.150 448.420 ;
        RECT 1451.830 434.420 1452.150 434.480 ;
        RECT 1451.635 434.280 1452.150 434.420 ;
        RECT 1451.830 434.220 1452.150 434.280 ;
        RECT 1451.845 379.680 1452.135 379.725 ;
        RECT 1452.290 379.680 1452.610 379.740 ;
        RECT 1451.845 379.540 1452.610 379.680 ;
        RECT 1451.845 379.495 1452.135 379.540 ;
        RECT 1452.290 379.480 1452.610 379.540 ;
        RECT 1451.830 303.520 1452.150 303.580 ;
        RECT 1453.210 303.520 1453.530 303.580 ;
        RECT 1451.830 303.380 1453.530 303.520 ;
        RECT 1451.830 303.320 1452.150 303.380 ;
        RECT 1453.210 303.320 1453.530 303.380 ;
        RECT 1451.830 214.100 1452.150 214.160 ;
        RECT 1452.290 214.100 1452.610 214.160 ;
        RECT 1451.830 213.960 1452.610 214.100 ;
        RECT 1451.830 213.900 1452.150 213.960 ;
        RECT 1452.290 213.900 1452.610 213.960 ;
        RECT 1451.830 193.360 1452.150 193.420 ;
        RECT 1452.290 193.360 1452.610 193.420 ;
        RECT 1451.830 193.220 1452.610 193.360 ;
        RECT 1451.830 193.160 1452.150 193.220 ;
        RECT 1452.290 193.160 1452.610 193.220 ;
        RECT 1452.290 96.800 1452.610 96.860 ;
        RECT 1452.750 96.800 1453.070 96.860 ;
        RECT 1452.290 96.660 1453.070 96.800 ;
        RECT 1452.290 96.600 1452.610 96.660 ;
        RECT 1452.750 96.600 1453.070 96.660 ;
        RECT 1451.830 48.180 1452.150 48.240 ;
        RECT 1451.635 48.040 1452.150 48.180 ;
        RECT 1451.830 47.980 1452.150 48.040 ;
        RECT 1126.610 42.060 1126.930 42.120 ;
        RECT 1451.845 42.060 1452.135 42.105 ;
        RECT 1126.610 41.920 1452.135 42.060 ;
        RECT 1126.610 41.860 1126.930 41.920 ;
        RECT 1451.845 41.875 1452.135 41.920 ;
      LAYER via ;
        RECT 1451.860 1635.100 1452.120 1635.360 ;
        RECT 1452.780 1545.000 1453.040 1545.260 ;
        RECT 1452.780 1490.260 1453.040 1490.520 ;
        RECT 1452.780 1489.580 1453.040 1489.840 ;
        RECT 1451.860 1393.700 1452.120 1393.960 ;
        RECT 1452.780 1393.700 1453.040 1393.960 ;
        RECT 1451.860 1345.420 1452.120 1345.680 ;
        RECT 1453.240 1345.420 1453.500 1345.680 ;
        RECT 1451.860 1297.140 1452.120 1297.400 ;
        RECT 1452.780 1297.140 1453.040 1297.400 ;
        RECT 1451.860 1269.600 1452.120 1269.860 ;
        RECT 1452.320 1269.260 1452.580 1269.520 ;
        RECT 1451.860 1152.300 1452.120 1152.560 ;
        RECT 1452.780 1152.300 1453.040 1152.560 ;
        RECT 1451.860 1007.120 1452.120 1007.380 ;
        RECT 1451.860 964.960 1452.120 965.220 ;
        RECT 1451.860 931.640 1452.120 931.900 ;
        RECT 1451.860 917.700 1452.120 917.960 ;
        RECT 1451.860 910.560 1452.120 910.820 ;
        RECT 1453.240 910.560 1453.500 910.820 ;
        RECT 1452.320 820.800 1452.580 821.060 ;
        RECT 1452.320 820.120 1452.580 820.380 ;
        RECT 1452.320 765.720 1452.580 765.980 ;
        RECT 1453.240 765.720 1453.500 765.980 ;
        RECT 1451.860 593.340 1452.120 593.600 ;
        RECT 1452.320 593.000 1452.580 593.260 ;
        RECT 1452.320 448.840 1452.580 449.100 ;
        RECT 1451.860 448.160 1452.120 448.420 ;
        RECT 1451.860 434.220 1452.120 434.480 ;
        RECT 1452.320 379.480 1452.580 379.740 ;
        RECT 1451.860 303.320 1452.120 303.580 ;
        RECT 1453.240 303.320 1453.500 303.580 ;
        RECT 1451.860 213.900 1452.120 214.160 ;
        RECT 1452.320 213.900 1452.580 214.160 ;
        RECT 1451.860 193.160 1452.120 193.420 ;
        RECT 1452.320 193.160 1452.580 193.420 ;
        RECT 1452.320 96.600 1452.580 96.860 ;
        RECT 1452.780 96.600 1453.040 96.860 ;
        RECT 1451.860 47.980 1452.120 48.240 ;
        RECT 1126.640 41.860 1126.900 42.120 ;
      LAYER met2 ;
        RECT 1453.690 1700.410 1453.970 1704.000 ;
        RECT 1453.300 1700.270 1453.970 1700.410 ;
        RECT 1453.300 1656.210 1453.440 1700.270 ;
        RECT 1453.690 1700.000 1453.970 1700.270 ;
        RECT 1451.920 1656.070 1453.440 1656.210 ;
        RECT 1451.920 1635.390 1452.060 1656.070 ;
        RECT 1451.860 1635.070 1452.120 1635.390 ;
        RECT 1452.780 1544.970 1453.040 1545.290 ;
        RECT 1452.840 1490.550 1452.980 1544.970 ;
        RECT 1452.780 1490.230 1453.040 1490.550 ;
        RECT 1452.780 1489.550 1453.040 1489.870 ;
        RECT 1452.840 1393.990 1452.980 1489.550 ;
        RECT 1451.860 1393.845 1452.120 1393.990 ;
        RECT 1451.850 1393.475 1452.130 1393.845 ;
        RECT 1452.780 1393.670 1453.040 1393.990 ;
        RECT 1453.230 1393.475 1453.510 1393.845 ;
        RECT 1453.300 1345.710 1453.440 1393.475 ;
        RECT 1451.860 1345.565 1452.120 1345.710 ;
        RECT 1451.850 1345.195 1452.130 1345.565 ;
        RECT 1452.770 1345.195 1453.050 1345.565 ;
        RECT 1453.240 1345.390 1453.500 1345.710 ;
        RECT 1452.840 1297.430 1452.980 1345.195 ;
        RECT 1451.860 1297.110 1452.120 1297.430 ;
        RECT 1452.780 1297.110 1453.040 1297.430 ;
        RECT 1451.920 1269.890 1452.060 1297.110 ;
        RECT 1451.860 1269.570 1452.120 1269.890 ;
        RECT 1452.320 1269.230 1452.580 1269.550 ;
        RECT 1452.380 1231.890 1452.520 1269.230 ;
        RECT 1452.380 1231.750 1452.980 1231.890 ;
        RECT 1452.840 1152.590 1452.980 1231.750 ;
        RECT 1451.860 1152.270 1452.120 1152.590 ;
        RECT 1452.780 1152.270 1453.040 1152.590 ;
        RECT 1451.920 1110.965 1452.060 1152.270 ;
        RECT 1451.850 1110.595 1452.130 1110.965 ;
        RECT 1453.230 1110.595 1453.510 1110.965 ;
        RECT 1453.300 1049.650 1453.440 1110.595 ;
        RECT 1452.840 1049.510 1453.440 1049.650 ;
        RECT 1452.840 1049.085 1452.980 1049.510 ;
        RECT 1451.850 1048.715 1452.130 1049.085 ;
        RECT 1452.770 1048.715 1453.050 1049.085 ;
        RECT 1451.920 1007.410 1452.060 1048.715 ;
        RECT 1451.860 1007.090 1452.120 1007.410 ;
        RECT 1451.860 964.930 1452.120 965.250 ;
        RECT 1451.920 931.930 1452.060 964.930 ;
        RECT 1451.860 931.610 1452.120 931.930 ;
        RECT 1451.860 917.670 1452.120 917.990 ;
        RECT 1451.920 910.850 1452.060 917.670 ;
        RECT 1451.860 910.530 1452.120 910.850 ;
        RECT 1453.240 910.530 1453.500 910.850 ;
        RECT 1453.300 862.765 1453.440 910.530 ;
        RECT 1452.310 862.395 1452.590 862.765 ;
        RECT 1453.230 862.395 1453.510 862.765 ;
        RECT 1452.380 821.090 1452.520 862.395 ;
        RECT 1452.320 820.770 1452.580 821.090 ;
        RECT 1452.320 820.090 1452.580 820.410 ;
        RECT 1452.380 766.010 1452.520 820.090 ;
        RECT 1452.320 765.690 1452.580 766.010 ;
        RECT 1453.240 765.690 1453.500 766.010 ;
        RECT 1453.300 717.925 1453.440 765.690 ;
        RECT 1451.850 717.555 1452.130 717.925 ;
        RECT 1453.230 717.555 1453.510 717.925 ;
        RECT 1451.920 593.630 1452.060 717.555 ;
        RECT 1451.860 593.310 1452.120 593.630 ;
        RECT 1452.320 592.970 1452.580 593.290 ;
        RECT 1452.380 548.490 1452.520 592.970 ;
        RECT 1452.380 548.350 1453.440 548.490 ;
        RECT 1453.300 494.090 1453.440 548.350 ;
        RECT 1452.840 493.950 1453.440 494.090 ;
        RECT 1452.840 483.210 1452.980 493.950 ;
        RECT 1452.380 483.070 1452.980 483.210 ;
        RECT 1452.380 449.130 1452.520 483.070 ;
        RECT 1452.320 448.810 1452.580 449.130 ;
        RECT 1451.860 448.130 1452.120 448.450 ;
        RECT 1451.920 434.510 1452.060 448.130 ;
        RECT 1451.860 434.190 1452.120 434.510 ;
        RECT 1452.320 379.450 1452.580 379.770 ;
        RECT 1452.380 311.170 1452.520 379.450 ;
        RECT 1451.920 311.030 1452.520 311.170 ;
        RECT 1451.920 303.610 1452.060 311.030 ;
        RECT 1451.860 303.290 1452.120 303.610 ;
        RECT 1453.240 303.290 1453.500 303.610 ;
        RECT 1453.300 255.525 1453.440 303.290 ;
        RECT 1452.310 255.155 1452.590 255.525 ;
        RECT 1453.230 255.155 1453.510 255.525 ;
        RECT 1452.380 214.190 1452.520 255.155 ;
        RECT 1451.860 213.870 1452.120 214.190 ;
        RECT 1452.320 213.870 1452.580 214.190 ;
        RECT 1451.920 193.450 1452.060 213.870 ;
        RECT 1451.860 193.130 1452.120 193.450 ;
        RECT 1452.320 193.130 1452.580 193.450 ;
        RECT 1452.380 145.365 1452.520 193.130 ;
        RECT 1452.310 144.995 1452.590 145.365 ;
        RECT 1452.770 143.635 1453.050 144.005 ;
        RECT 1452.840 96.890 1452.980 143.635 ;
        RECT 1452.320 96.570 1452.580 96.890 ;
        RECT 1452.780 96.570 1453.040 96.890 ;
        RECT 1452.380 62.970 1452.520 96.570 ;
        RECT 1452.380 62.830 1452.980 62.970 ;
        RECT 1452.840 48.690 1452.980 62.830 ;
        RECT 1451.920 48.550 1452.980 48.690 ;
        RECT 1451.920 48.270 1452.060 48.550 ;
        RECT 1451.860 47.950 1452.120 48.270 ;
        RECT 1126.640 41.830 1126.900 42.150 ;
        RECT 1126.700 2.400 1126.840 41.830 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
      LAYER via2 ;
        RECT 1451.850 1393.520 1452.130 1393.800 ;
        RECT 1453.230 1393.520 1453.510 1393.800 ;
        RECT 1451.850 1345.240 1452.130 1345.520 ;
        RECT 1452.770 1345.240 1453.050 1345.520 ;
        RECT 1451.850 1110.640 1452.130 1110.920 ;
        RECT 1453.230 1110.640 1453.510 1110.920 ;
        RECT 1451.850 1048.760 1452.130 1049.040 ;
        RECT 1452.770 1048.760 1453.050 1049.040 ;
        RECT 1452.310 862.440 1452.590 862.720 ;
        RECT 1453.230 862.440 1453.510 862.720 ;
        RECT 1451.850 717.600 1452.130 717.880 ;
        RECT 1453.230 717.600 1453.510 717.880 ;
        RECT 1452.310 255.200 1452.590 255.480 ;
        RECT 1453.230 255.200 1453.510 255.480 ;
        RECT 1452.310 145.040 1452.590 145.320 ;
        RECT 1452.770 143.680 1453.050 143.960 ;
      LAYER met3 ;
        RECT 1451.825 1393.810 1452.155 1393.825 ;
        RECT 1453.205 1393.810 1453.535 1393.825 ;
        RECT 1451.825 1393.510 1453.535 1393.810 ;
        RECT 1451.825 1393.495 1452.155 1393.510 ;
        RECT 1453.205 1393.495 1453.535 1393.510 ;
        RECT 1451.825 1345.530 1452.155 1345.545 ;
        RECT 1452.745 1345.530 1453.075 1345.545 ;
        RECT 1451.825 1345.230 1453.075 1345.530 ;
        RECT 1451.825 1345.215 1452.155 1345.230 ;
        RECT 1452.745 1345.215 1453.075 1345.230 ;
        RECT 1451.825 1110.930 1452.155 1110.945 ;
        RECT 1453.205 1110.930 1453.535 1110.945 ;
        RECT 1451.825 1110.630 1453.535 1110.930 ;
        RECT 1451.825 1110.615 1452.155 1110.630 ;
        RECT 1453.205 1110.615 1453.535 1110.630 ;
        RECT 1451.825 1049.050 1452.155 1049.065 ;
        RECT 1452.745 1049.050 1453.075 1049.065 ;
        RECT 1451.825 1048.750 1453.075 1049.050 ;
        RECT 1451.825 1048.735 1452.155 1048.750 ;
        RECT 1452.745 1048.735 1453.075 1048.750 ;
        RECT 1452.285 862.730 1452.615 862.745 ;
        RECT 1453.205 862.730 1453.535 862.745 ;
        RECT 1452.285 862.430 1453.535 862.730 ;
        RECT 1452.285 862.415 1452.615 862.430 ;
        RECT 1453.205 862.415 1453.535 862.430 ;
        RECT 1451.825 717.890 1452.155 717.905 ;
        RECT 1453.205 717.890 1453.535 717.905 ;
        RECT 1451.825 717.590 1453.535 717.890 ;
        RECT 1451.825 717.575 1452.155 717.590 ;
        RECT 1453.205 717.575 1453.535 717.590 ;
        RECT 1452.285 255.490 1452.615 255.505 ;
        RECT 1453.205 255.490 1453.535 255.505 ;
        RECT 1452.285 255.190 1453.535 255.490 ;
        RECT 1452.285 255.175 1452.615 255.190 ;
        RECT 1453.205 255.175 1453.535 255.190 ;
        RECT 1452.285 145.330 1452.615 145.345 ;
        RECT 1451.150 145.030 1452.615 145.330 ;
        RECT 1451.150 143.970 1451.450 145.030 ;
        RECT 1452.285 145.015 1452.615 145.030 ;
        RECT 1452.745 143.970 1453.075 143.985 ;
        RECT 1451.150 143.670 1453.075 143.970 ;
        RECT 1452.745 143.655 1453.075 143.670 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1449.990 1678.480 1450.310 1678.540 ;
        RECT 1454.130 1678.480 1454.450 1678.540 ;
        RECT 1449.990 1678.340 1454.450 1678.480 ;
        RECT 1449.990 1678.280 1450.310 1678.340 ;
        RECT 1454.130 1678.280 1454.450 1678.340 ;
        RECT 1126.610 42.400 1126.930 42.460 ;
        RECT 1449.990 42.400 1450.310 42.460 ;
        RECT 1126.610 42.260 1450.310 42.400 ;
        RECT 1126.610 42.200 1126.930 42.260 ;
        RECT 1449.990 42.200 1450.310 42.260 ;
      LAYER via ;
        RECT 1450.020 1678.280 1450.280 1678.540 ;
        RECT 1454.160 1678.280 1454.420 1678.540 ;
        RECT 1126.640 42.200 1126.900 42.460 ;
        RECT 1450.020 42.200 1450.280 42.460 ;
      LAYER met2 ;
        RECT 1455.070 1700.410 1455.350 1704.000 ;
        RECT 1454.220 1700.270 1455.350 1700.410 ;
        RECT 1454.220 1678.570 1454.360 1700.270 ;
        RECT 1455.070 1700.000 1455.350 1700.270 ;
        RECT 1450.020 1678.250 1450.280 1678.570 ;
        RECT 1454.160 1678.250 1454.420 1678.570 ;
        RECT 1450.080 42.490 1450.220 1678.250 ;
        RECT 1126.640 42.170 1126.900 42.490 ;
        RECT 1450.020 42.170 1450.280 42.490 ;
        RECT 1126.700 2.400 1126.840 42.170 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1144.550 41.720 1144.870 41.780 ;
        RECT 1457.810 41.720 1458.130 41.780 ;
        RECT 1144.550 41.580 1458.130 41.720 ;
        RECT 1144.550 41.520 1144.870 41.580 ;
        RECT 1457.810 41.520 1458.130 41.580 ;
      LAYER via ;
        RECT 1144.580 41.520 1144.840 41.780 ;
        RECT 1457.840 41.520 1458.100 41.780 ;
=======
      LAYER li1 ;
        RECT 1457.885 1442.025 1458.055 1490.475 ;
      LAYER mcon ;
        RECT 1457.885 1490.305 1458.055 1490.475 ;
      LAYER met1 ;
        RECT 1457.810 1539.080 1458.130 1539.140 ;
        RECT 1458.730 1539.080 1459.050 1539.140 ;
        RECT 1457.810 1538.940 1459.050 1539.080 ;
        RECT 1457.810 1538.880 1458.130 1538.940 ;
        RECT 1458.730 1538.880 1459.050 1538.940 ;
        RECT 1457.810 1497.600 1458.130 1497.660 ;
        RECT 1458.270 1497.600 1458.590 1497.660 ;
        RECT 1457.810 1497.460 1458.590 1497.600 ;
        RECT 1457.810 1497.400 1458.130 1497.460 ;
        RECT 1458.270 1497.400 1458.590 1497.460 ;
        RECT 1457.825 1490.460 1458.115 1490.505 ;
        RECT 1458.270 1490.460 1458.590 1490.520 ;
        RECT 1457.825 1490.320 1458.590 1490.460 ;
        RECT 1457.825 1490.275 1458.115 1490.320 ;
        RECT 1458.270 1490.260 1458.590 1490.320 ;
        RECT 1457.810 1442.180 1458.130 1442.240 ;
        RECT 1457.615 1442.040 1458.130 1442.180 ;
        RECT 1457.810 1441.980 1458.130 1442.040 ;
        RECT 1456.890 821.000 1457.210 821.060 ;
        RECT 1457.810 821.000 1458.130 821.060 ;
        RECT 1456.890 820.860 1458.130 821.000 ;
        RECT 1456.890 820.800 1457.210 820.860 ;
        RECT 1457.810 820.800 1458.130 820.860 ;
        RECT 1458.270 145.080 1458.590 145.140 ;
        RECT 1458.730 145.080 1459.050 145.140 ;
        RECT 1458.270 144.940 1459.050 145.080 ;
        RECT 1458.270 144.880 1458.590 144.940 ;
        RECT 1458.730 144.880 1459.050 144.940 ;
        RECT 1457.810 96.800 1458.130 96.860 ;
        RECT 1458.730 96.800 1459.050 96.860 ;
        RECT 1457.810 96.660 1459.050 96.800 ;
        RECT 1457.810 96.600 1458.130 96.660 ;
        RECT 1458.730 96.600 1459.050 96.660 ;
        RECT 1144.550 42.060 1144.870 42.120 ;
        RECT 1457.350 42.060 1457.670 42.120 ;
        RECT 1144.550 41.920 1457.670 42.060 ;
        RECT 1144.550 41.860 1144.870 41.920 ;
        RECT 1457.350 41.860 1457.670 41.920 ;
      LAYER via ;
        RECT 1457.840 1538.880 1458.100 1539.140 ;
        RECT 1458.760 1538.880 1459.020 1539.140 ;
        RECT 1457.840 1497.400 1458.100 1497.660 ;
        RECT 1458.300 1497.400 1458.560 1497.660 ;
        RECT 1458.300 1490.260 1458.560 1490.520 ;
        RECT 1457.840 1441.980 1458.100 1442.240 ;
        RECT 1456.920 820.800 1457.180 821.060 ;
        RECT 1457.840 820.800 1458.100 821.060 ;
        RECT 1458.300 144.880 1458.560 145.140 ;
        RECT 1458.760 144.880 1459.020 145.140 ;
        RECT 1457.840 96.600 1458.100 96.860 ;
        RECT 1458.760 96.600 1459.020 96.860 ;
        RECT 1144.580 41.860 1144.840 42.120 ;
        RECT 1457.380 41.860 1457.640 42.120 ;
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1460.130 1700.410 1460.410 1704.000 ;
        RECT 1458.820 1700.270 1460.410 1700.410 ;
        RECT 1458.820 1539.170 1458.960 1700.270 ;
        RECT 1460.130 1700.000 1460.410 1700.270 ;
        RECT 1457.840 1538.850 1458.100 1539.170 ;
        RECT 1458.760 1538.850 1459.020 1539.170 ;
        RECT 1457.900 1497.690 1458.040 1538.850 ;
        RECT 1457.840 1497.370 1458.100 1497.690 ;
        RECT 1458.300 1497.370 1458.560 1497.690 ;
        RECT 1458.360 1490.550 1458.500 1497.370 ;
        RECT 1458.300 1490.230 1458.560 1490.550 ;
        RECT 1457.840 1441.950 1458.100 1442.270 ;
        RECT 1457.900 1414.810 1458.040 1441.950 ;
        RECT 1457.440 1414.670 1458.040 1414.810 ;
        RECT 1457.440 1414.130 1457.580 1414.670 ;
        RECT 1457.440 1413.990 1458.040 1414.130 ;
        RECT 1457.900 1318.250 1458.040 1413.990 ;
        RECT 1457.440 1318.110 1458.040 1318.250 ;
        RECT 1457.440 1317.570 1457.580 1318.110 ;
        RECT 1457.440 1317.430 1458.040 1317.570 ;
        RECT 1457.900 1221.690 1458.040 1317.430 ;
        RECT 1457.440 1221.550 1458.040 1221.690 ;
        RECT 1457.440 1221.010 1457.580 1221.550 ;
        RECT 1457.440 1220.870 1458.040 1221.010 ;
        RECT 1457.900 1125.130 1458.040 1220.870 ;
        RECT 1457.440 1124.990 1458.040 1125.130 ;
        RECT 1457.440 1124.450 1457.580 1124.990 ;
        RECT 1457.440 1124.310 1458.040 1124.450 ;
        RECT 1457.900 1028.570 1458.040 1124.310 ;
        RECT 1457.440 1028.430 1458.040 1028.570 ;
        RECT 1457.440 1027.890 1457.580 1028.430 ;
        RECT 1457.440 1027.750 1458.040 1027.890 ;
        RECT 1457.900 932.010 1458.040 1027.750 ;
        RECT 1457.440 931.870 1458.040 932.010 ;
        RECT 1457.440 931.330 1457.580 931.870 ;
        RECT 1457.440 931.190 1458.040 931.330 ;
        RECT 1457.900 835.450 1458.040 931.190 ;
        RECT 1457.440 835.310 1458.040 835.450 ;
        RECT 1457.440 834.770 1457.580 835.310 ;
        RECT 1457.440 834.630 1458.040 834.770 ;
        RECT 1457.900 821.090 1458.040 834.630 ;
        RECT 1456.920 820.770 1457.180 821.090 ;
        RECT 1457.840 820.770 1458.100 821.090 ;
        RECT 1456.980 773.005 1457.120 820.770 ;
        RECT 1456.910 772.635 1457.190 773.005 ;
        RECT 1457.830 772.635 1458.110 773.005 ;
        RECT 1457.900 642.330 1458.040 772.635 ;
        RECT 1457.440 642.190 1458.040 642.330 ;
        RECT 1457.440 641.650 1457.580 642.190 ;
        RECT 1457.440 641.510 1458.040 641.650 ;
        RECT 1457.900 545.770 1458.040 641.510 ;
        RECT 1457.440 545.630 1458.040 545.770 ;
        RECT 1457.440 545.090 1457.580 545.630 ;
        RECT 1457.440 544.950 1458.040 545.090 ;
        RECT 1457.900 449.210 1458.040 544.950 ;
        RECT 1457.440 449.070 1458.040 449.210 ;
        RECT 1457.440 448.530 1457.580 449.070 ;
        RECT 1457.440 448.390 1458.040 448.530 ;
        RECT 1457.900 351.970 1458.040 448.390 ;
        RECT 1457.440 351.830 1458.040 351.970 ;
        RECT 1457.440 351.290 1457.580 351.830 ;
        RECT 1457.440 351.150 1458.040 351.290 ;
        RECT 1457.900 255.410 1458.040 351.150 ;
        RECT 1457.440 255.270 1458.040 255.410 ;
        RECT 1457.440 254.730 1457.580 255.270 ;
        RECT 1457.440 254.590 1458.040 254.730 ;
        RECT 1457.900 169.050 1458.040 254.590 ;
        RECT 1457.900 168.910 1458.500 169.050 ;
        RECT 1458.360 145.170 1458.500 168.910 ;
        RECT 1458.300 144.850 1458.560 145.170 ;
        RECT 1458.760 144.850 1459.020 145.170 ;
        RECT 1458.820 96.890 1458.960 144.850 ;
        RECT 1457.840 96.570 1458.100 96.890 ;
        RECT 1458.760 96.570 1459.020 96.890 ;
        RECT 1457.900 72.490 1458.040 96.570 ;
        RECT 1457.440 72.350 1458.040 72.490 ;
        RECT 1457.440 42.150 1457.580 72.350 ;
        RECT 1144.580 41.830 1144.840 42.150 ;
        RECT 1457.380 41.830 1457.640 42.150 ;
        RECT 1144.640 2.400 1144.780 41.830 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 1456.910 772.680 1457.190 772.960 ;
        RECT 1457.830 772.680 1458.110 772.960 ;
      LAYER met3 ;
        RECT 1456.885 772.970 1457.215 772.985 ;
        RECT 1457.805 772.970 1458.135 772.985 ;
        RECT 1456.885 772.670 1458.135 772.970 ;
        RECT 1456.885 772.655 1457.215 772.670 ;
        RECT 1457.805 772.655 1458.135 772.670 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1162.490 44.780 1162.810 44.840 ;
        RECT 1464.710 44.780 1465.030 44.840 ;
        RECT 1162.490 44.640 1465.030 44.780 ;
        RECT 1162.490 44.580 1162.810 44.640 ;
        RECT 1464.710 44.580 1465.030 44.640 ;
      LAYER via ;
        RECT 1162.520 44.580 1162.780 44.840 ;
        RECT 1464.740 44.580 1465.000 44.840 ;
      LAYER met2 ;
        RECT 1464.730 1700.000 1465.010 1704.000 ;
        RECT 1464.800 44.870 1464.940 1700.000 ;
        RECT 1162.520 44.550 1162.780 44.870 ;
        RECT 1464.740 44.550 1465.000 44.870 ;
        RECT 1162.580 2.400 1162.720 44.550 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1331.770 1678.140 1332.090 1678.200 ;
        RECT 1333.150 1678.140 1333.470 1678.200 ;
        RECT 1331.770 1678.000 1333.470 1678.140 ;
        RECT 1331.770 1677.940 1332.090 1678.000 ;
        RECT 1333.150 1677.940 1333.470 1678.000 ;
        RECT 680.410 47.500 680.730 47.560 ;
        RECT 1331.770 47.500 1332.090 47.560 ;
        RECT 680.410 47.360 1332.090 47.500 ;
        RECT 680.410 47.300 680.730 47.360 ;
        RECT 1331.770 47.300 1332.090 47.360 ;
      LAYER via ;
        RECT 1331.800 1677.940 1332.060 1678.200 ;
        RECT 1333.180 1677.940 1333.440 1678.200 ;
        RECT 680.440 47.300 680.700 47.560 ;
        RECT 1331.800 47.300 1332.060 47.560 ;
      LAYER met2 ;
        RECT 1334.090 1700.410 1334.370 1704.000 ;
        RECT 1333.240 1700.270 1334.370 1700.410 ;
        RECT 1333.240 1678.230 1333.380 1700.270 ;
        RECT 1334.090 1700.000 1334.370 1700.270 ;
        RECT 1331.800 1677.910 1332.060 1678.230 ;
        RECT 1333.180 1677.910 1333.440 1678.230 ;
        RECT 1331.860 47.590 1332.000 1677.910 ;
        RECT 680.440 47.270 680.700 47.590 ;
        RECT 1331.800 47.270 1332.060 47.590 ;
        RECT 680.500 2.400 680.640 47.270 ;
        RECT 680.290 -4.800 680.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 0.300 ;
=======
      LAYER li1 ;
        RECT 1465.245 386.325 1465.415 410.635 ;
      LAYER mcon ;
        RECT 1465.245 410.465 1465.415 410.635 ;
      LAYER met1 ;
        RECT 1464.710 1607.900 1465.030 1608.160 ;
        RECT 1464.800 1607.480 1464.940 1607.900 ;
        RECT 1464.710 1607.220 1465.030 1607.480 ;
        RECT 1464.710 1497.060 1465.030 1497.320 ;
        RECT 1464.800 1496.920 1464.940 1497.060 ;
        RECT 1465.630 1496.920 1465.950 1496.980 ;
        RECT 1464.800 1496.780 1465.950 1496.920 ;
        RECT 1465.630 1496.720 1465.950 1496.780 ;
        RECT 1465.170 1111.020 1465.490 1111.080 ;
        RECT 1466.090 1111.020 1466.410 1111.080 ;
        RECT 1465.170 1110.880 1466.410 1111.020 ;
        RECT 1465.170 1110.820 1465.490 1110.880 ;
        RECT 1466.090 1110.820 1466.410 1110.880 ;
        RECT 1465.170 869.620 1465.490 869.680 ;
        RECT 1465.630 869.620 1465.950 869.680 ;
        RECT 1465.170 869.480 1465.950 869.620 ;
        RECT 1465.170 869.420 1465.490 869.480 ;
        RECT 1465.630 869.420 1465.950 869.480 ;
        RECT 1465.185 410.620 1465.475 410.665 ;
        RECT 1465.630 410.620 1465.950 410.680 ;
        RECT 1465.185 410.480 1465.950 410.620 ;
        RECT 1465.185 410.435 1465.475 410.480 ;
        RECT 1465.630 410.420 1465.950 410.480 ;
        RECT 1465.170 386.480 1465.490 386.540 ;
        RECT 1464.975 386.340 1465.490 386.480 ;
        RECT 1465.170 386.280 1465.490 386.340 ;
        RECT 1179.970 17.240 1180.290 17.300 ;
        RECT 1465.170 17.240 1465.490 17.300 ;
        RECT 1179.970 17.100 1465.490 17.240 ;
        RECT 1179.970 17.040 1180.290 17.100 ;
        RECT 1465.170 17.040 1465.490 17.100 ;
      LAYER via ;
        RECT 1464.740 1607.900 1465.000 1608.160 ;
        RECT 1464.740 1607.220 1465.000 1607.480 ;
        RECT 1464.740 1497.060 1465.000 1497.320 ;
        RECT 1465.660 1496.720 1465.920 1496.980 ;
        RECT 1465.200 1110.820 1465.460 1111.080 ;
        RECT 1466.120 1110.820 1466.380 1111.080 ;
        RECT 1465.200 869.420 1465.460 869.680 ;
        RECT 1465.660 869.420 1465.920 869.680 ;
        RECT 1465.660 410.420 1465.920 410.680 ;
        RECT 1465.200 386.280 1465.460 386.540 ;
        RECT 1180.000 17.040 1180.260 17.300 ;
        RECT 1465.200 17.040 1465.460 17.300 ;
      LAYER met2 ;
        RECT 1468.410 1700.410 1468.690 1704.000 ;
        RECT 1467.560 1700.270 1468.690 1700.410 ;
        RECT 1467.560 1677.290 1467.700 1700.270 ;
        RECT 1468.410 1700.000 1468.690 1700.270 ;
        RECT 1464.800 1677.150 1467.700 1677.290 ;
        RECT 1464.800 1608.190 1464.940 1677.150 ;
        RECT 1464.740 1607.870 1465.000 1608.190 ;
        RECT 1464.740 1607.190 1465.000 1607.510 ;
        RECT 1464.800 1497.350 1464.940 1607.190 ;
        RECT 1464.740 1497.030 1465.000 1497.350 ;
        RECT 1465.660 1496.690 1465.920 1497.010 ;
        RECT 1465.720 1366.530 1465.860 1496.690 ;
        RECT 1464.800 1366.390 1465.860 1366.530 ;
        RECT 1464.800 1365.850 1464.940 1366.390 ;
        RECT 1464.800 1365.710 1465.400 1365.850 ;
        RECT 1465.260 1297.170 1465.400 1365.710 ;
        RECT 1465.260 1297.030 1465.860 1297.170 ;
        RECT 1465.720 1207.410 1465.860 1297.030 ;
        RECT 1465.720 1207.270 1466.320 1207.410 ;
        RECT 1466.180 1200.725 1466.320 1207.270 ;
        RECT 1465.190 1200.355 1465.470 1200.725 ;
        RECT 1466.110 1200.355 1466.390 1200.725 ;
        RECT 1465.260 1157.770 1465.400 1200.355 ;
        RECT 1465.260 1157.630 1466.320 1157.770 ;
        RECT 1466.180 1111.110 1466.320 1157.630 ;
        RECT 1465.200 1110.790 1465.460 1111.110 ;
        RECT 1466.120 1110.790 1466.380 1111.110 ;
        RECT 1465.260 1014.290 1465.400 1110.790 ;
        RECT 1465.260 1014.150 1465.860 1014.290 ;
        RECT 1465.720 869.710 1465.860 1014.150 ;
        RECT 1465.200 869.390 1465.460 869.710 ;
        RECT 1465.660 869.390 1465.920 869.710 ;
        RECT 1465.260 786.490 1465.400 869.390 ;
        RECT 1464.800 786.350 1465.400 786.490 ;
        RECT 1464.800 785.130 1464.940 786.350 ;
        RECT 1464.800 784.990 1465.400 785.130 ;
        RECT 1465.260 594.050 1465.400 784.990 ;
        RECT 1464.800 593.910 1465.400 594.050 ;
        RECT 1464.800 593.370 1464.940 593.910 ;
        RECT 1464.800 593.230 1465.400 593.370 ;
        RECT 1465.260 483.210 1465.400 593.230 ;
        RECT 1465.260 483.070 1465.860 483.210 ;
        RECT 1465.720 410.710 1465.860 483.070 ;
        RECT 1465.660 410.390 1465.920 410.710 ;
        RECT 1465.200 386.250 1465.460 386.570 ;
        RECT 1465.260 207.130 1465.400 386.250 ;
        RECT 1464.800 206.990 1465.400 207.130 ;
        RECT 1464.800 206.450 1464.940 206.990 ;
        RECT 1464.800 206.310 1465.400 206.450 ;
        RECT 1465.260 110.570 1465.400 206.310 ;
        RECT 1464.800 110.430 1465.400 110.570 ;
        RECT 1464.800 109.890 1464.940 110.430 ;
        RECT 1464.800 109.750 1465.400 109.890 ;
        RECT 1465.260 17.330 1465.400 109.750 ;
        RECT 1180.000 17.010 1180.260 17.330 ;
        RECT 1465.200 17.010 1465.460 17.330 ;
        RECT 1180.060 2.400 1180.200 17.010 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
      LAYER via2 ;
        RECT 1465.190 1200.400 1465.470 1200.680 ;
        RECT 1466.110 1200.400 1466.390 1200.680 ;
      LAYER met3 ;
        RECT 1465.165 1200.690 1465.495 1200.705 ;
        RECT 1466.085 1200.690 1466.415 1200.705 ;
        RECT 1465.165 1200.390 1466.415 1200.690 ;
        RECT 1465.165 1200.375 1465.495 1200.390 ;
        RECT 1466.085 1200.375 1466.415 1200.390 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1179.970 41.720 1180.290 41.780 ;
        RECT 1470.690 41.720 1471.010 41.780 ;
        RECT 1179.970 41.580 1471.010 41.720 ;
        RECT 1179.970 41.520 1180.290 41.580 ;
        RECT 1470.690 41.520 1471.010 41.580 ;
      LAYER via ;
        RECT 1180.000 41.520 1180.260 41.780 ;
        RECT 1470.720 41.520 1470.980 41.780 ;
      LAYER met2 ;
        RECT 1469.790 1700.410 1470.070 1704.000 ;
        RECT 1469.790 1700.270 1470.920 1700.410 ;
        RECT 1469.790 1700.000 1470.070 1700.270 ;
        RECT 1470.780 41.810 1470.920 1700.270 ;
        RECT 1180.000 41.490 1180.260 41.810 ;
        RECT 1470.720 41.490 1470.980 41.810 ;
        RECT 1180.060 2.400 1180.200 41.490 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1197.790 -4.800 1198.350 0.300 ;
=======
        RECT 1473.010 1700.410 1473.290 1704.000 ;
        RECT 1472.160 1700.270 1473.290 1700.410 ;
        RECT 1472.160 18.885 1472.300 1700.270 ;
        RECT 1473.010 1700.000 1473.290 1700.270 ;
        RECT 1197.930 18.515 1198.210 18.885 ;
        RECT 1472.090 18.515 1472.370 18.885 ;
        RECT 1198.000 2.400 1198.140 18.515 ;
=======
      LAYER li1 ;
        RECT 1473.525 1607.605 1473.695 1635.315 ;
        RECT 1473.985 1490.645 1474.155 1538.755 ;
        RECT 1473.065 1317.245 1473.235 1352.435 ;
        RECT 1473.525 1207.425 1473.695 1297.015 ;
        RECT 1473.525 386.325 1473.695 434.775 ;
        RECT 1473.525 186.405 1473.695 234.515 ;
        RECT 1473.065 89.845 1473.235 121.635 ;
      LAYER mcon ;
        RECT 1473.525 1635.145 1473.695 1635.315 ;
        RECT 1473.985 1538.585 1474.155 1538.755 ;
        RECT 1473.065 1352.265 1473.235 1352.435 ;
        RECT 1473.525 1296.845 1473.695 1297.015 ;
        RECT 1473.525 434.605 1473.695 434.775 ;
        RECT 1473.525 234.345 1473.695 234.515 ;
        RECT 1473.065 121.465 1473.235 121.635 ;
      LAYER met1 ;
        RECT 1473.450 1683.920 1473.770 1683.980 ;
        RECT 1473.910 1683.920 1474.230 1683.980 ;
        RECT 1473.450 1683.780 1474.230 1683.920 ;
        RECT 1473.450 1683.720 1473.770 1683.780 ;
        RECT 1473.910 1683.720 1474.230 1683.780 ;
        RECT 1473.910 1635.980 1474.230 1636.040 ;
        RECT 1474.370 1635.980 1474.690 1636.040 ;
        RECT 1473.910 1635.840 1474.690 1635.980 ;
        RECT 1473.910 1635.780 1474.230 1635.840 ;
        RECT 1474.370 1635.780 1474.690 1635.840 ;
        RECT 1473.465 1635.300 1473.755 1635.345 ;
        RECT 1473.910 1635.300 1474.230 1635.360 ;
        RECT 1473.465 1635.160 1474.230 1635.300 ;
        RECT 1473.465 1635.115 1473.755 1635.160 ;
        RECT 1473.910 1635.100 1474.230 1635.160 ;
        RECT 1473.450 1607.760 1473.770 1607.820 ;
        RECT 1473.255 1607.620 1473.770 1607.760 ;
        RECT 1473.450 1607.560 1473.770 1607.620 ;
        RECT 1473.450 1545.340 1473.770 1545.600 ;
        RECT 1472.530 1544.860 1472.850 1544.920 ;
        RECT 1473.540 1544.860 1473.680 1545.340 ;
        RECT 1472.530 1544.720 1473.680 1544.860 ;
        RECT 1472.530 1544.660 1472.850 1544.720 ;
        RECT 1473.910 1538.740 1474.230 1538.800 ;
        RECT 1473.715 1538.600 1474.230 1538.740 ;
        RECT 1473.910 1538.540 1474.230 1538.600 ;
        RECT 1473.910 1490.800 1474.230 1490.860 ;
        RECT 1473.715 1490.660 1474.230 1490.800 ;
        RECT 1473.910 1490.600 1474.230 1490.660 ;
        RECT 1473.450 1442.520 1473.770 1442.580 ;
        RECT 1474.370 1442.520 1474.690 1442.580 ;
        RECT 1473.450 1442.380 1474.690 1442.520 ;
        RECT 1473.450 1442.320 1473.770 1442.380 ;
        RECT 1474.370 1442.320 1474.690 1442.380 ;
        RECT 1473.910 1414.640 1474.230 1414.700 ;
        RECT 1473.080 1414.500 1474.230 1414.640 ;
        RECT 1473.080 1414.020 1473.220 1414.500 ;
        RECT 1473.910 1414.440 1474.230 1414.500 ;
        RECT 1472.990 1413.760 1473.310 1414.020 ;
        RECT 1472.990 1352.420 1473.310 1352.480 ;
        RECT 1472.795 1352.280 1473.310 1352.420 ;
        RECT 1472.990 1352.220 1473.310 1352.280 ;
        RECT 1473.005 1317.400 1473.295 1317.445 ;
        RECT 1473.450 1317.400 1473.770 1317.460 ;
        RECT 1473.005 1317.260 1473.770 1317.400 ;
        RECT 1473.005 1317.215 1473.295 1317.260 ;
        RECT 1473.450 1317.200 1473.770 1317.260 ;
        RECT 1473.450 1297.000 1473.770 1297.060 ;
        RECT 1473.255 1296.860 1473.770 1297.000 ;
        RECT 1473.450 1296.800 1473.770 1296.860 ;
        RECT 1473.465 1207.580 1473.755 1207.625 ;
        RECT 1473.910 1207.580 1474.230 1207.640 ;
        RECT 1473.465 1207.440 1474.230 1207.580 ;
        RECT 1473.465 1207.395 1473.755 1207.440 ;
        RECT 1473.910 1207.380 1474.230 1207.440 ;
        RECT 1472.530 1062.740 1472.850 1062.800 ;
        RECT 1473.450 1062.740 1473.770 1062.800 ;
        RECT 1472.530 1062.600 1473.770 1062.740 ;
        RECT 1472.530 1062.540 1472.850 1062.600 ;
        RECT 1473.450 1062.540 1473.770 1062.600 ;
        RECT 1472.990 931.640 1473.310 931.900 ;
        RECT 1473.080 931.160 1473.220 931.640 ;
        RECT 1473.450 931.160 1473.770 931.220 ;
        RECT 1473.080 931.020 1473.770 931.160 ;
        RECT 1473.450 930.960 1473.770 931.020 ;
        RECT 1473.450 910.760 1473.770 910.820 ;
        RECT 1474.370 910.760 1474.690 910.820 ;
        RECT 1473.450 910.620 1474.690 910.760 ;
        RECT 1473.450 910.560 1473.770 910.620 ;
        RECT 1474.370 910.560 1474.690 910.620 ;
        RECT 1472.990 834.940 1473.310 835.000 ;
        RECT 1473.910 834.940 1474.230 835.000 ;
        RECT 1472.990 834.800 1474.230 834.940 ;
        RECT 1472.990 834.740 1473.310 834.800 ;
        RECT 1473.910 834.740 1474.230 834.800 ;
        RECT 1473.910 787.140 1474.230 787.400 ;
        RECT 1473.450 786.320 1473.770 786.380 ;
        RECT 1474.000 786.320 1474.140 787.140 ;
        RECT 1473.450 786.180 1474.140 786.320 ;
        RECT 1473.450 786.120 1473.770 786.180 ;
        RECT 1473.910 627.880 1474.230 627.940 ;
        RECT 1474.830 627.880 1475.150 627.940 ;
        RECT 1473.910 627.740 1475.150 627.880 ;
        RECT 1473.910 627.680 1474.230 627.740 ;
        RECT 1474.830 627.680 1475.150 627.740 ;
        RECT 1472.990 483.040 1473.310 483.100 ;
        RECT 1473.910 483.040 1474.230 483.100 ;
        RECT 1472.990 482.900 1474.230 483.040 ;
        RECT 1472.990 482.840 1473.310 482.900 ;
        RECT 1473.910 482.840 1474.230 482.900 ;
        RECT 1473.465 434.760 1473.755 434.805 ;
        RECT 1473.910 434.760 1474.230 434.820 ;
        RECT 1473.465 434.620 1474.230 434.760 ;
        RECT 1473.465 434.575 1473.755 434.620 ;
        RECT 1473.910 434.560 1474.230 434.620 ;
        RECT 1473.450 386.480 1473.770 386.540 ;
        RECT 1473.255 386.340 1473.770 386.480 ;
        RECT 1473.450 386.280 1473.770 386.340 ;
        RECT 1473.450 255.380 1473.770 255.640 ;
        RECT 1473.540 254.900 1473.680 255.380 ;
        RECT 1473.910 254.900 1474.230 254.960 ;
        RECT 1473.540 254.760 1474.230 254.900 ;
        RECT 1473.910 254.700 1474.230 254.760 ;
        RECT 1473.465 234.500 1473.755 234.545 ;
        RECT 1473.910 234.500 1474.230 234.560 ;
        RECT 1473.465 234.360 1474.230 234.500 ;
        RECT 1473.465 234.315 1473.755 234.360 ;
        RECT 1473.910 234.300 1474.230 234.360 ;
        RECT 1473.450 186.560 1473.770 186.620 ;
        RECT 1473.255 186.420 1473.770 186.560 ;
        RECT 1473.450 186.360 1473.770 186.420 ;
        RECT 1473.005 121.620 1473.295 121.665 ;
        RECT 1473.450 121.620 1473.770 121.680 ;
        RECT 1473.005 121.480 1473.770 121.620 ;
        RECT 1473.005 121.435 1473.295 121.480 ;
        RECT 1473.450 121.420 1473.770 121.480 ;
        RECT 1472.990 90.000 1473.310 90.060 ;
        RECT 1472.795 89.860 1473.310 90.000 ;
        RECT 1472.990 89.800 1473.310 89.860 ;
        RECT 1197.910 45.120 1198.230 45.180 ;
        RECT 1472.990 45.120 1473.310 45.180 ;
        RECT 1197.910 44.980 1473.310 45.120 ;
        RECT 1197.910 44.920 1198.230 44.980 ;
        RECT 1472.990 44.920 1473.310 44.980 ;
      LAYER via ;
        RECT 1473.480 1683.720 1473.740 1683.980 ;
        RECT 1473.940 1683.720 1474.200 1683.980 ;
        RECT 1473.940 1635.780 1474.200 1636.040 ;
        RECT 1474.400 1635.780 1474.660 1636.040 ;
        RECT 1473.940 1635.100 1474.200 1635.360 ;
        RECT 1473.480 1607.560 1473.740 1607.820 ;
        RECT 1473.480 1545.340 1473.740 1545.600 ;
        RECT 1472.560 1544.660 1472.820 1544.920 ;
        RECT 1473.940 1538.540 1474.200 1538.800 ;
        RECT 1473.940 1490.600 1474.200 1490.860 ;
        RECT 1473.480 1442.320 1473.740 1442.580 ;
        RECT 1474.400 1442.320 1474.660 1442.580 ;
        RECT 1473.940 1414.440 1474.200 1414.700 ;
        RECT 1473.020 1413.760 1473.280 1414.020 ;
        RECT 1473.020 1352.220 1473.280 1352.480 ;
        RECT 1473.480 1317.200 1473.740 1317.460 ;
        RECT 1473.480 1296.800 1473.740 1297.060 ;
        RECT 1473.940 1207.380 1474.200 1207.640 ;
        RECT 1472.560 1062.540 1472.820 1062.800 ;
        RECT 1473.480 1062.540 1473.740 1062.800 ;
        RECT 1473.020 931.640 1473.280 931.900 ;
        RECT 1473.480 930.960 1473.740 931.220 ;
        RECT 1473.480 910.560 1473.740 910.820 ;
        RECT 1474.400 910.560 1474.660 910.820 ;
        RECT 1473.020 834.740 1473.280 835.000 ;
        RECT 1473.940 834.740 1474.200 835.000 ;
        RECT 1473.940 787.140 1474.200 787.400 ;
        RECT 1473.480 786.120 1473.740 786.380 ;
        RECT 1473.940 627.680 1474.200 627.940 ;
        RECT 1474.860 627.680 1475.120 627.940 ;
        RECT 1473.020 482.840 1473.280 483.100 ;
        RECT 1473.940 482.840 1474.200 483.100 ;
        RECT 1473.940 434.560 1474.200 434.820 ;
        RECT 1473.480 386.280 1473.740 386.540 ;
        RECT 1473.480 255.380 1473.740 255.640 ;
        RECT 1473.940 254.700 1474.200 254.960 ;
        RECT 1473.940 234.300 1474.200 234.560 ;
        RECT 1473.480 186.360 1473.740 186.620 ;
        RECT 1473.480 121.420 1473.740 121.680 ;
        RECT 1473.020 89.800 1473.280 90.060 ;
        RECT 1197.940 44.920 1198.200 45.180 ;
        RECT 1473.020 44.920 1473.280 45.180 ;
      LAYER met2 ;
        RECT 1474.390 1700.410 1474.670 1704.000 ;
        RECT 1473.540 1700.270 1474.670 1700.410 ;
        RECT 1473.540 1684.010 1473.680 1700.270 ;
        RECT 1474.390 1700.000 1474.670 1700.270 ;
        RECT 1473.480 1683.690 1473.740 1684.010 ;
        RECT 1473.940 1683.690 1474.200 1684.010 ;
        RECT 1474.000 1683.525 1474.140 1683.690 ;
        RECT 1473.930 1683.155 1474.210 1683.525 ;
        RECT 1474.390 1682.475 1474.670 1682.845 ;
        RECT 1474.460 1636.070 1474.600 1682.475 ;
        RECT 1473.940 1635.750 1474.200 1636.070 ;
        RECT 1474.400 1635.750 1474.660 1636.070 ;
        RECT 1474.000 1635.390 1474.140 1635.750 ;
        RECT 1473.940 1635.070 1474.200 1635.390 ;
        RECT 1473.480 1607.530 1473.740 1607.850 ;
        RECT 1473.540 1545.630 1473.680 1607.530 ;
        RECT 1473.480 1545.310 1473.740 1545.630 ;
        RECT 1472.560 1544.630 1472.820 1544.950 ;
        RECT 1472.620 1539.365 1472.760 1544.630 ;
        RECT 1472.550 1538.995 1472.830 1539.365 ;
        RECT 1473.930 1538.995 1474.210 1539.365 ;
        RECT 1474.000 1538.830 1474.140 1538.995 ;
        RECT 1473.940 1538.510 1474.200 1538.830 ;
        RECT 1473.940 1490.570 1474.200 1490.890 ;
        RECT 1474.000 1463.090 1474.140 1490.570 ;
        RECT 1474.000 1462.950 1474.600 1463.090 ;
        RECT 1474.460 1442.610 1474.600 1462.950 ;
        RECT 1473.480 1442.290 1473.740 1442.610 ;
        RECT 1474.400 1442.290 1474.660 1442.610 ;
        RECT 1473.540 1442.010 1473.680 1442.290 ;
        RECT 1473.540 1441.870 1474.140 1442.010 ;
        RECT 1474.000 1414.730 1474.140 1441.870 ;
        RECT 1473.940 1414.410 1474.200 1414.730 ;
        RECT 1473.020 1413.730 1473.280 1414.050 ;
        RECT 1473.080 1352.510 1473.220 1413.730 ;
        RECT 1473.020 1352.190 1473.280 1352.510 ;
        RECT 1473.480 1317.170 1473.740 1317.490 ;
        RECT 1473.540 1297.090 1473.680 1317.170 ;
        RECT 1473.480 1296.770 1473.740 1297.090 ;
        RECT 1473.940 1207.350 1474.200 1207.670 ;
        RECT 1474.000 1173.410 1474.140 1207.350 ;
        RECT 1473.080 1173.270 1474.140 1173.410 ;
        RECT 1473.080 1124.450 1473.220 1173.270 ;
        RECT 1473.080 1124.310 1474.140 1124.450 ;
        RECT 1474.000 1110.965 1474.140 1124.310 ;
        RECT 1472.550 1110.595 1472.830 1110.965 ;
        RECT 1473.930 1110.595 1474.210 1110.965 ;
        RECT 1472.620 1062.830 1472.760 1110.595 ;
        RECT 1472.560 1062.510 1472.820 1062.830 ;
        RECT 1473.480 1062.510 1473.740 1062.830 ;
        RECT 1473.540 980.290 1473.680 1062.510 ;
        RECT 1473.080 980.150 1473.680 980.290 ;
        RECT 1473.080 931.930 1473.220 980.150 ;
        RECT 1473.020 931.610 1473.280 931.930 ;
        RECT 1473.480 930.930 1473.740 931.250 ;
        RECT 1473.540 910.850 1473.680 930.930 ;
        RECT 1473.480 910.530 1473.740 910.850 ;
        RECT 1474.400 910.530 1474.660 910.850 ;
        RECT 1474.460 862.765 1474.600 910.530 ;
        RECT 1473.010 862.395 1473.290 862.765 ;
        RECT 1474.390 862.395 1474.670 862.765 ;
        RECT 1473.080 835.030 1473.220 862.395 ;
        RECT 1473.020 834.710 1473.280 835.030 ;
        RECT 1473.940 834.710 1474.200 835.030 ;
        RECT 1474.000 787.430 1474.140 834.710 ;
        RECT 1473.940 787.110 1474.200 787.430 ;
        RECT 1473.480 786.090 1473.740 786.410 ;
        RECT 1473.540 690.610 1473.680 786.090 ;
        RECT 1473.080 690.470 1473.680 690.610 ;
        RECT 1473.080 641.650 1473.220 690.470 ;
        RECT 1473.080 641.510 1474.140 641.650 ;
        RECT 1474.000 627.970 1474.140 641.510 ;
        RECT 1473.940 627.650 1474.200 627.970 ;
        RECT 1474.860 627.650 1475.120 627.970 ;
        RECT 1474.920 579.885 1475.060 627.650 ;
        RECT 1473.470 579.515 1473.750 579.885 ;
        RECT 1474.850 579.515 1475.130 579.885 ;
        RECT 1473.540 497.490 1473.680 579.515 ;
        RECT 1473.080 497.350 1473.680 497.490 ;
        RECT 1473.080 483.130 1473.220 497.350 ;
        RECT 1473.020 482.810 1473.280 483.130 ;
        RECT 1473.940 482.810 1474.200 483.130 ;
        RECT 1474.000 434.850 1474.140 482.810 ;
        RECT 1473.940 434.530 1474.200 434.850 ;
        RECT 1473.480 386.250 1473.740 386.570 ;
        RECT 1473.540 352.085 1473.680 386.250 ;
        RECT 1472.550 351.715 1472.830 352.085 ;
        RECT 1473.470 351.715 1473.750 352.085 ;
        RECT 1472.620 328.170 1472.760 351.715 ;
        RECT 1472.620 328.030 1473.680 328.170 ;
        RECT 1473.540 255.670 1473.680 328.030 ;
        RECT 1473.480 255.350 1473.740 255.670 ;
        RECT 1473.940 254.670 1474.200 254.990 ;
        RECT 1474.000 234.590 1474.140 254.670 ;
        RECT 1473.940 234.270 1474.200 234.590 ;
        RECT 1473.480 186.330 1473.740 186.650 ;
        RECT 1473.540 121.710 1473.680 186.330 ;
        RECT 1473.480 121.390 1473.740 121.710 ;
        RECT 1473.020 89.770 1473.280 90.090 ;
        RECT 1473.080 45.210 1473.220 89.770 ;
        RECT 1197.940 44.890 1198.200 45.210 ;
        RECT 1473.020 44.890 1473.280 45.210 ;
        RECT 1198.000 2.400 1198.140 44.890 ;
>>>>>>> re-updated local openlane
        RECT 1197.790 -4.800 1198.350 2.400 ;
      LAYER via2 ;
        RECT 1473.930 1683.200 1474.210 1683.480 ;
        RECT 1474.390 1682.520 1474.670 1682.800 ;
        RECT 1472.550 1539.040 1472.830 1539.320 ;
        RECT 1473.930 1539.040 1474.210 1539.320 ;
        RECT 1472.550 1110.640 1472.830 1110.920 ;
        RECT 1473.930 1110.640 1474.210 1110.920 ;
        RECT 1473.010 862.440 1473.290 862.720 ;
        RECT 1474.390 862.440 1474.670 862.720 ;
        RECT 1473.470 579.560 1473.750 579.840 ;
        RECT 1474.850 579.560 1475.130 579.840 ;
        RECT 1472.550 351.760 1472.830 352.040 ;
        RECT 1473.470 351.760 1473.750 352.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1197.905 18.850 1198.235 18.865 ;
        RECT 1472.065 18.850 1472.395 18.865 ;
        RECT 1197.905 18.550 1472.395 18.850 ;
        RECT 1197.905 18.535 1198.235 18.550 ;
        RECT 1472.065 18.535 1472.395 18.550 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1473.905 1683.490 1474.235 1683.505 ;
        RECT 1473.230 1683.190 1474.235 1683.490 ;
        RECT 1473.230 1682.810 1473.530 1683.190 ;
        RECT 1473.905 1683.175 1474.235 1683.190 ;
        RECT 1474.365 1682.810 1474.695 1682.825 ;
        RECT 1473.230 1682.510 1474.695 1682.810 ;
        RECT 1474.365 1682.495 1474.695 1682.510 ;
        RECT 1472.525 1539.330 1472.855 1539.345 ;
        RECT 1473.905 1539.330 1474.235 1539.345 ;
        RECT 1472.525 1539.030 1474.235 1539.330 ;
        RECT 1472.525 1539.015 1472.855 1539.030 ;
        RECT 1473.905 1539.015 1474.235 1539.030 ;
        RECT 1472.525 1110.930 1472.855 1110.945 ;
        RECT 1473.905 1110.930 1474.235 1110.945 ;
        RECT 1472.525 1110.630 1474.235 1110.930 ;
        RECT 1472.525 1110.615 1472.855 1110.630 ;
        RECT 1473.905 1110.615 1474.235 1110.630 ;
        RECT 1472.985 862.730 1473.315 862.745 ;
        RECT 1474.365 862.730 1474.695 862.745 ;
        RECT 1472.985 862.430 1474.695 862.730 ;
        RECT 1472.985 862.415 1473.315 862.430 ;
        RECT 1474.365 862.415 1474.695 862.430 ;
        RECT 1473.445 579.850 1473.775 579.865 ;
        RECT 1474.825 579.850 1475.155 579.865 ;
        RECT 1473.445 579.550 1475.155 579.850 ;
        RECT 1473.445 579.535 1473.775 579.550 ;
        RECT 1474.825 579.535 1475.155 579.550 ;
        RECT 1472.525 352.050 1472.855 352.065 ;
        RECT 1473.445 352.050 1473.775 352.065 ;
        RECT 1472.525 351.750 1473.775 352.050 ;
        RECT 1472.525 351.735 1472.855 351.750 ;
        RECT 1473.445 351.735 1473.775 351.750 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1215.850 45.460 1216.170 45.520 ;
        RECT 1477.130 45.460 1477.450 45.520 ;
        RECT 1215.850 45.320 1477.450 45.460 ;
        RECT 1215.850 45.260 1216.170 45.320 ;
        RECT 1477.130 45.260 1477.450 45.320 ;
      LAYER via ;
        RECT 1215.880 45.260 1216.140 45.520 ;
        RECT 1477.160 45.260 1477.420 45.520 ;
      LAYER met2 ;
        RECT 1479.450 1700.410 1479.730 1704.000 ;
        RECT 1478.140 1700.270 1479.730 1700.410 ;
        RECT 1478.140 1678.140 1478.280 1700.270 ;
        RECT 1479.450 1700.000 1479.730 1700.270 ;
        RECT 1477.220 1678.000 1478.280 1678.140 ;
        RECT 1477.220 45.550 1477.360 1678.000 ;
        RECT 1215.880 45.230 1216.140 45.550 ;
        RECT 1477.160 45.230 1477.420 45.550 ;
        RECT 1215.940 2.400 1216.080 45.230 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1215.870 19.920 1216.150 20.200 ;
        RECT 1476.690 19.920 1476.970 20.200 ;
      LAYER met3 ;
        RECT 1215.845 20.210 1216.175 20.225 ;
        RECT 1476.665 20.210 1476.995 20.225 ;
        RECT 1215.845 19.910 1476.995 20.210 ;
        RECT 1215.845 19.895 1216.175 19.910 ;
        RECT 1476.665 19.895 1476.995 19.910 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 0.300 ;
=======
      LAYER li1 ;
        RECT 1438.105 1684.445 1438.275 1687.335 ;
      LAYER mcon ;
        RECT 1438.105 1687.165 1438.275 1687.335 ;
      LAYER met1 ;
        RECT 1259.550 1687.320 1259.870 1687.380 ;
        RECT 1438.045 1687.320 1438.335 1687.365 ;
        RECT 1259.550 1687.180 1438.335 1687.320 ;
        RECT 1259.550 1687.120 1259.870 1687.180 ;
        RECT 1438.045 1687.135 1438.335 1687.180 ;
        RECT 1438.045 1684.600 1438.335 1684.645 ;
        RECT 1438.045 1684.460 1472.760 1684.600 ;
        RECT 1438.045 1684.415 1438.335 1684.460 ;
        RECT 1472.620 1684.260 1472.760 1684.460 ;
        RECT 1482.650 1684.260 1482.970 1684.320 ;
        RECT 1472.620 1684.120 1482.970 1684.260 ;
        RECT 1482.650 1684.060 1482.970 1684.120 ;
        RECT 1233.790 20.300 1234.110 20.360 ;
        RECT 1259.550 20.300 1259.870 20.360 ;
        RECT 1233.790 20.160 1259.870 20.300 ;
        RECT 1233.790 20.100 1234.110 20.160 ;
        RECT 1259.550 20.100 1259.870 20.160 ;
      LAYER via ;
        RECT 1259.580 1687.120 1259.840 1687.380 ;
        RECT 1482.680 1684.060 1482.940 1684.320 ;
        RECT 1233.820 20.100 1234.080 20.360 ;
        RECT 1259.580 20.100 1259.840 20.360 ;
      LAYER met2 ;
        RECT 1482.670 1700.000 1482.950 1704.000 ;
        RECT 1259.580 1687.090 1259.840 1687.410 ;
        RECT 1259.640 20.390 1259.780 1687.090 ;
        RECT 1482.740 1684.350 1482.880 1700.000 ;
        RECT 1482.680 1684.030 1482.940 1684.350 ;
        RECT 1233.820 20.070 1234.080 20.390 ;
        RECT 1259.580 20.070 1259.840 20.390 ;
        RECT 1233.880 2.400 1234.020 20.070 ;
=======
      LAYER met1 ;
        RECT 1233.790 59.060 1234.110 59.120 ;
        RECT 1484.950 59.060 1485.270 59.120 ;
        RECT 1233.790 58.920 1485.270 59.060 ;
        RECT 1233.790 58.860 1234.110 58.920 ;
        RECT 1484.950 58.860 1485.270 58.920 ;
      LAYER via ;
        RECT 1233.820 58.860 1234.080 59.120 ;
        RECT 1484.980 58.860 1485.240 59.120 ;
      LAYER met2 ;
        RECT 1484.050 1700.410 1484.330 1704.000 ;
        RECT 1484.050 1700.270 1485.180 1700.410 ;
        RECT 1484.050 1700.000 1484.330 1700.270 ;
        RECT 1485.040 59.150 1485.180 1700.270 ;
        RECT 1233.820 58.830 1234.080 59.150 ;
        RECT 1484.980 58.830 1485.240 59.150 ;
        RECT 1233.880 2.400 1234.020 58.830 ;
>>>>>>> re-updated local openlane
        RECT 1233.670 -4.800 1234.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1483.570 1678.480 1483.890 1678.540 ;
        RECT 1487.710 1678.480 1488.030 1678.540 ;
        RECT 1483.570 1678.340 1488.030 1678.480 ;
        RECT 1483.570 1678.280 1483.890 1678.340 ;
        RECT 1487.710 1678.280 1488.030 1678.340 ;
        RECT 1251.730 17.240 1252.050 17.300 ;
        RECT 1483.570 17.240 1483.890 17.300 ;
        RECT 1251.730 17.100 1483.890 17.240 ;
        RECT 1251.730 17.040 1252.050 17.100 ;
        RECT 1483.570 17.040 1483.890 17.100 ;
      LAYER via ;
        RECT 1483.600 1678.280 1483.860 1678.540 ;
        RECT 1487.740 1678.280 1488.000 1678.540 ;
        RECT 1251.760 17.040 1252.020 17.300 ;
        RECT 1483.600 17.040 1483.860 17.300 ;
      LAYER met2 ;
        RECT 1489.110 1700.410 1489.390 1704.000 ;
        RECT 1487.800 1700.270 1489.390 1700.410 ;
        RECT 1487.800 1678.570 1487.940 1700.270 ;
        RECT 1489.110 1700.000 1489.390 1700.270 ;
        RECT 1483.600 1678.250 1483.860 1678.570 ;
        RECT 1487.740 1678.250 1488.000 1678.570 ;
        RECT 1483.660 17.330 1483.800 1678.250 ;
        RECT 1251.760 17.010 1252.020 17.330 ;
        RECT 1483.600 17.010 1483.860 17.330 ;
        RECT 1251.820 2.400 1251.960 17.010 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 0.300 ;
=======
      LAYER li1 ;
        RECT 1341.965 1642.965 1342.135 1689.035 ;
        RECT 1308.385 1580.065 1308.555 1594.175 ;
        RECT 1308.385 1145.885 1308.555 1193.655 ;
        RECT 1309.305 807.245 1309.475 821.355 ;
        RECT 1309.305 421.345 1309.475 469.115 ;
        RECT 1309.765 379.185 1309.935 420.835 ;
        RECT 1307.925 34.425 1308.095 82.875 ;
      LAYER mcon ;
        RECT 1341.965 1688.865 1342.135 1689.035 ;
        RECT 1308.385 1594.005 1308.555 1594.175 ;
        RECT 1308.385 1193.485 1308.555 1193.655 ;
        RECT 1309.305 821.185 1309.475 821.355 ;
        RECT 1309.305 468.945 1309.475 469.115 ;
        RECT 1309.765 420.665 1309.935 420.835 ;
        RECT 1307.925 82.705 1308.095 82.875 ;
      LAYER met1 ;
        RECT 1341.905 1689.020 1342.195 1689.065 ;
        RECT 1492.310 1689.020 1492.630 1689.080 ;
        RECT 1341.905 1688.880 1492.630 1689.020 ;
        RECT 1341.905 1688.835 1342.195 1688.880 ;
        RECT 1492.310 1688.820 1492.630 1688.880 ;
        RECT 1308.770 1643.120 1309.090 1643.180 ;
        RECT 1341.905 1643.120 1342.195 1643.165 ;
        RECT 1308.770 1642.980 1342.195 1643.120 ;
        RECT 1308.770 1642.920 1309.090 1642.980 ;
        RECT 1341.905 1642.935 1342.195 1642.980 ;
        RECT 1308.325 1594.160 1308.615 1594.205 ;
        RECT 1308.770 1594.160 1309.090 1594.220 ;
        RECT 1308.325 1594.020 1309.090 1594.160 ;
        RECT 1308.325 1593.975 1308.615 1594.020 ;
        RECT 1308.770 1593.960 1309.090 1594.020 ;
        RECT 1308.310 1580.220 1308.630 1580.280 ;
        RECT 1308.115 1580.080 1308.630 1580.220 ;
        RECT 1308.310 1580.020 1308.630 1580.080 ;
        RECT 1307.850 1490.460 1308.170 1490.520 ;
        RECT 1308.770 1490.460 1309.090 1490.520 ;
        RECT 1307.850 1490.320 1309.090 1490.460 ;
        RECT 1307.850 1490.260 1308.170 1490.320 ;
        RECT 1308.770 1490.260 1309.090 1490.320 ;
        RECT 1308.310 1249.060 1308.630 1249.120 ;
        RECT 1308.770 1249.060 1309.090 1249.120 ;
        RECT 1308.310 1248.920 1309.090 1249.060 ;
        RECT 1308.310 1248.860 1308.630 1248.920 ;
        RECT 1308.770 1248.860 1309.090 1248.920 ;
        RECT 1308.325 1193.640 1308.615 1193.685 ;
        RECT 1308.770 1193.640 1309.090 1193.700 ;
        RECT 1308.325 1193.500 1309.090 1193.640 ;
        RECT 1308.325 1193.455 1308.615 1193.500 ;
        RECT 1308.770 1193.440 1309.090 1193.500 ;
        RECT 1308.310 1146.040 1308.630 1146.100 ;
        RECT 1308.115 1145.900 1308.630 1146.040 ;
        RECT 1308.310 1145.840 1308.630 1145.900 ;
        RECT 1307.850 1145.360 1308.170 1145.420 ;
        RECT 1308.310 1145.360 1308.630 1145.420 ;
        RECT 1307.850 1145.220 1308.630 1145.360 ;
        RECT 1307.850 1145.160 1308.170 1145.220 ;
        RECT 1308.310 1145.160 1308.630 1145.220 ;
        RECT 1308.310 1072.940 1308.630 1073.000 ;
        RECT 1309.230 1072.940 1309.550 1073.000 ;
        RECT 1308.310 1072.800 1309.550 1072.940 ;
        RECT 1308.310 1072.740 1308.630 1072.800 ;
        RECT 1309.230 1072.740 1309.550 1072.800 ;
        RECT 1308.310 917.900 1308.630 917.960 ;
        RECT 1308.770 917.900 1309.090 917.960 ;
        RECT 1308.310 917.760 1309.090 917.900 ;
        RECT 1308.310 917.700 1308.630 917.760 ;
        RECT 1308.770 917.700 1309.090 917.760 ;
        RECT 1308.770 910.760 1309.090 910.820 ;
        RECT 1309.230 910.760 1309.550 910.820 ;
        RECT 1308.770 910.620 1309.550 910.760 ;
        RECT 1308.770 910.560 1309.090 910.620 ;
        RECT 1309.230 910.560 1309.550 910.620 ;
        RECT 1309.230 821.340 1309.550 821.400 ;
        RECT 1309.035 821.200 1309.550 821.340 ;
        RECT 1309.230 821.140 1309.550 821.200 ;
        RECT 1309.230 807.400 1309.550 807.460 ;
        RECT 1309.035 807.260 1309.550 807.400 ;
        RECT 1309.230 807.200 1309.550 807.260 ;
        RECT 1308.770 613.940 1309.090 614.000 ;
        RECT 1309.230 613.940 1309.550 614.000 ;
        RECT 1308.770 613.800 1309.550 613.940 ;
        RECT 1308.770 613.740 1309.090 613.800 ;
        RECT 1309.230 613.740 1309.550 613.800 ;
        RECT 1308.770 524.520 1309.090 524.580 ;
        RECT 1309.230 524.520 1309.550 524.580 ;
        RECT 1308.770 524.380 1309.550 524.520 ;
        RECT 1308.770 524.320 1309.090 524.380 ;
        RECT 1309.230 524.320 1309.550 524.380 ;
        RECT 1308.770 517.380 1309.090 517.440 ;
        RECT 1309.230 517.380 1309.550 517.440 ;
        RECT 1308.770 517.240 1309.550 517.380 ;
        RECT 1308.770 517.180 1309.090 517.240 ;
        RECT 1309.230 517.180 1309.550 517.240 ;
        RECT 1309.230 469.100 1309.550 469.160 ;
        RECT 1309.035 468.960 1309.550 469.100 ;
        RECT 1309.230 468.900 1309.550 468.960 ;
        RECT 1309.245 421.500 1309.535 421.545 ;
        RECT 1309.690 421.500 1310.010 421.560 ;
        RECT 1309.245 421.360 1310.010 421.500 ;
        RECT 1309.245 421.315 1309.535 421.360 ;
        RECT 1309.690 421.300 1310.010 421.360 ;
        RECT 1309.690 420.820 1310.010 420.880 ;
        RECT 1309.495 420.680 1310.010 420.820 ;
        RECT 1309.690 420.620 1310.010 420.680 ;
        RECT 1309.690 379.340 1310.010 379.400 ;
        RECT 1309.495 379.200 1310.010 379.340 ;
        RECT 1309.690 379.140 1310.010 379.200 ;
        RECT 1308.770 324.600 1309.090 324.660 ;
        RECT 1309.690 324.600 1310.010 324.660 ;
        RECT 1308.770 324.460 1310.010 324.600 ;
        RECT 1308.770 324.400 1309.090 324.460 ;
        RECT 1309.690 324.400 1310.010 324.460 ;
        RECT 1308.310 282.780 1308.630 282.840 ;
        RECT 1308.770 282.780 1309.090 282.840 ;
        RECT 1308.310 282.640 1309.090 282.780 ;
        RECT 1308.310 282.580 1308.630 282.640 ;
        RECT 1308.770 282.580 1309.090 282.640 ;
        RECT 1308.310 179.420 1308.630 179.480 ;
        RECT 1309.230 179.420 1309.550 179.480 ;
        RECT 1308.310 179.280 1309.550 179.420 ;
        RECT 1308.310 179.220 1308.630 179.280 ;
        RECT 1309.230 179.220 1309.550 179.280 ;
        RECT 1307.865 82.860 1308.155 82.905 ;
        RECT 1308.310 82.860 1308.630 82.920 ;
        RECT 1307.865 82.720 1308.630 82.860 ;
        RECT 1307.865 82.675 1308.155 82.720 ;
        RECT 1308.310 82.660 1308.630 82.720 ;
        RECT 1307.850 34.580 1308.170 34.640 ;
        RECT 1307.655 34.440 1308.170 34.580 ;
        RECT 1307.850 34.380 1308.170 34.440 ;
        RECT 1269.210 19.620 1269.530 19.680 ;
        RECT 1307.850 19.620 1308.170 19.680 ;
        RECT 1269.210 19.480 1308.170 19.620 ;
        RECT 1269.210 19.420 1269.530 19.480 ;
        RECT 1307.850 19.420 1308.170 19.480 ;
      LAYER via ;
        RECT 1492.340 1688.820 1492.600 1689.080 ;
        RECT 1308.800 1642.920 1309.060 1643.180 ;
        RECT 1308.800 1593.960 1309.060 1594.220 ;
        RECT 1308.340 1580.020 1308.600 1580.280 ;
        RECT 1307.880 1490.260 1308.140 1490.520 ;
        RECT 1308.800 1490.260 1309.060 1490.520 ;
        RECT 1308.340 1248.860 1308.600 1249.120 ;
        RECT 1308.800 1248.860 1309.060 1249.120 ;
        RECT 1308.800 1193.440 1309.060 1193.700 ;
        RECT 1308.340 1145.840 1308.600 1146.100 ;
        RECT 1307.880 1145.160 1308.140 1145.420 ;
        RECT 1308.340 1145.160 1308.600 1145.420 ;
        RECT 1308.340 1072.740 1308.600 1073.000 ;
        RECT 1309.260 1072.740 1309.520 1073.000 ;
        RECT 1308.340 917.700 1308.600 917.960 ;
        RECT 1308.800 917.700 1309.060 917.960 ;
        RECT 1308.800 910.560 1309.060 910.820 ;
        RECT 1309.260 910.560 1309.520 910.820 ;
        RECT 1309.260 821.140 1309.520 821.400 ;
        RECT 1309.260 807.200 1309.520 807.460 ;
        RECT 1308.800 613.740 1309.060 614.000 ;
        RECT 1309.260 613.740 1309.520 614.000 ;
        RECT 1308.800 524.320 1309.060 524.580 ;
        RECT 1309.260 524.320 1309.520 524.580 ;
        RECT 1308.800 517.180 1309.060 517.440 ;
        RECT 1309.260 517.180 1309.520 517.440 ;
        RECT 1309.260 468.900 1309.520 469.160 ;
        RECT 1309.720 421.300 1309.980 421.560 ;
        RECT 1309.720 420.620 1309.980 420.880 ;
        RECT 1309.720 379.140 1309.980 379.400 ;
        RECT 1308.800 324.400 1309.060 324.660 ;
        RECT 1309.720 324.400 1309.980 324.660 ;
        RECT 1308.340 282.580 1308.600 282.840 ;
        RECT 1308.800 282.580 1309.060 282.840 ;
        RECT 1308.340 179.220 1308.600 179.480 ;
        RECT 1309.260 179.220 1309.520 179.480 ;
        RECT 1308.340 82.660 1308.600 82.920 ;
        RECT 1307.880 34.380 1308.140 34.640 ;
        RECT 1269.240 19.420 1269.500 19.680 ;
        RECT 1307.880 19.420 1308.140 19.680 ;
      LAYER met2 ;
        RECT 1492.330 1700.000 1492.610 1704.000 ;
        RECT 1492.400 1689.110 1492.540 1700.000 ;
        RECT 1492.340 1688.790 1492.600 1689.110 ;
        RECT 1308.800 1642.890 1309.060 1643.210 ;
        RECT 1308.860 1594.250 1309.000 1642.890 ;
        RECT 1308.800 1593.930 1309.060 1594.250 ;
        RECT 1308.340 1579.990 1308.600 1580.310 ;
        RECT 1308.400 1514.770 1308.540 1579.990 ;
        RECT 1308.400 1514.630 1309.460 1514.770 ;
        RECT 1309.320 1510.690 1309.460 1514.630 ;
        RECT 1308.860 1510.550 1309.460 1510.690 ;
        RECT 1308.860 1490.550 1309.000 1510.550 ;
        RECT 1307.880 1490.230 1308.140 1490.550 ;
        RECT 1308.800 1490.230 1309.060 1490.550 ;
        RECT 1307.940 1435.325 1308.080 1490.230 ;
        RECT 1307.870 1434.955 1308.150 1435.325 ;
        RECT 1309.250 1434.955 1309.530 1435.325 ;
        RECT 1309.320 1387.725 1309.460 1434.955 ;
        RECT 1309.250 1387.355 1309.530 1387.725 ;
        RECT 1309.250 1386.675 1309.530 1387.045 ;
        RECT 1309.320 1363.130 1309.460 1386.675 ;
        RECT 1308.860 1362.990 1309.460 1363.130 ;
        RECT 1308.860 1249.150 1309.000 1362.990 ;
        RECT 1308.340 1249.005 1308.600 1249.150 ;
        RECT 1308.330 1248.635 1308.610 1249.005 ;
        RECT 1308.800 1248.830 1309.060 1249.150 ;
        RECT 1309.250 1248.635 1309.530 1249.005 ;
        RECT 1309.320 1221.010 1309.460 1248.635 ;
        RECT 1308.860 1220.870 1309.460 1221.010 ;
        RECT 1308.860 1193.730 1309.000 1220.870 ;
        RECT 1308.800 1193.410 1309.060 1193.730 ;
        RECT 1308.340 1145.810 1308.600 1146.130 ;
        RECT 1308.400 1145.450 1308.540 1145.810 ;
        RECT 1307.880 1145.130 1308.140 1145.450 ;
        RECT 1308.340 1145.130 1308.600 1145.450 ;
        RECT 1307.940 1097.365 1308.080 1145.130 ;
        RECT 1307.870 1096.995 1308.150 1097.365 ;
        RECT 1309.250 1096.995 1309.530 1097.365 ;
        RECT 1309.320 1073.030 1309.460 1096.995 ;
        RECT 1308.340 1072.710 1308.600 1073.030 ;
        RECT 1309.260 1072.710 1309.520 1073.030 ;
        RECT 1308.400 917.990 1308.540 1072.710 ;
        RECT 1308.340 917.670 1308.600 917.990 ;
        RECT 1308.800 917.670 1309.060 917.990 ;
        RECT 1308.860 910.850 1309.000 917.670 ;
        RECT 1308.800 910.530 1309.060 910.850 ;
        RECT 1309.260 910.530 1309.520 910.850 ;
        RECT 1309.320 821.430 1309.460 910.530 ;
        RECT 1309.260 821.110 1309.520 821.430 ;
        RECT 1309.260 807.170 1309.520 807.490 ;
        RECT 1309.320 782.410 1309.460 807.170 ;
        RECT 1308.400 782.270 1309.460 782.410 ;
        RECT 1308.400 741.610 1308.540 782.270 ;
        RECT 1308.400 741.470 1309.000 741.610 ;
        RECT 1308.860 669.530 1309.000 741.470 ;
        RECT 1308.400 669.390 1309.000 669.530 ;
        RECT 1308.400 644.370 1308.540 669.390 ;
        RECT 1308.400 644.230 1309.000 644.370 ;
        RECT 1308.860 614.030 1309.000 644.230 ;
        RECT 1308.800 613.710 1309.060 614.030 ;
        RECT 1309.260 613.710 1309.520 614.030 ;
        RECT 1309.320 524.610 1309.460 613.710 ;
        RECT 1308.800 524.290 1309.060 524.610 ;
        RECT 1309.260 524.290 1309.520 524.610 ;
        RECT 1308.860 517.470 1309.000 524.290 ;
        RECT 1308.800 517.150 1309.060 517.470 ;
        RECT 1309.260 517.150 1309.520 517.470 ;
        RECT 1309.320 469.190 1309.460 517.150 ;
        RECT 1309.260 468.870 1309.520 469.190 ;
        RECT 1309.720 421.270 1309.980 421.590 ;
        RECT 1309.780 420.910 1309.920 421.270 ;
        RECT 1309.720 420.590 1309.980 420.910 ;
        RECT 1309.720 379.110 1309.980 379.430 ;
        RECT 1309.780 324.690 1309.920 379.110 ;
        RECT 1308.800 324.370 1309.060 324.690 ;
        RECT 1309.720 324.370 1309.980 324.690 ;
        RECT 1308.860 282.870 1309.000 324.370 ;
        RECT 1308.340 282.550 1308.600 282.870 ;
        RECT 1308.800 282.550 1309.060 282.870 ;
        RECT 1308.400 258.130 1308.540 282.550 ;
        RECT 1308.400 257.990 1309.000 258.130 ;
        RECT 1308.860 186.730 1309.000 257.990 ;
        RECT 1308.400 186.590 1309.000 186.730 ;
        RECT 1308.400 179.510 1308.540 186.590 ;
        RECT 1308.340 179.190 1308.600 179.510 ;
        RECT 1309.260 179.190 1309.520 179.510 ;
        RECT 1309.320 107.170 1309.460 179.190 ;
        RECT 1308.400 107.030 1309.460 107.170 ;
        RECT 1308.400 82.950 1308.540 107.030 ;
        RECT 1308.340 82.630 1308.600 82.950 ;
        RECT 1307.880 34.350 1308.140 34.670 ;
        RECT 1307.940 19.710 1308.080 34.350 ;
        RECT 1269.240 19.390 1269.500 19.710 ;
        RECT 1307.880 19.390 1308.140 19.710 ;
        RECT 1269.300 2.400 1269.440 19.390 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
      LAYER via2 ;
        RECT 1307.870 1435.000 1308.150 1435.280 ;
        RECT 1309.250 1435.000 1309.530 1435.280 ;
        RECT 1309.250 1387.400 1309.530 1387.680 ;
        RECT 1309.250 1386.720 1309.530 1387.000 ;
        RECT 1308.330 1248.680 1308.610 1248.960 ;
        RECT 1309.250 1248.680 1309.530 1248.960 ;
        RECT 1307.870 1097.040 1308.150 1097.320 ;
        RECT 1309.250 1097.040 1309.530 1097.320 ;
      LAYER met3 ;
        RECT 1307.845 1435.290 1308.175 1435.305 ;
        RECT 1309.225 1435.290 1309.555 1435.305 ;
        RECT 1307.845 1434.990 1309.555 1435.290 ;
        RECT 1307.845 1434.975 1308.175 1434.990 ;
        RECT 1309.225 1434.975 1309.555 1434.990 ;
        RECT 1309.225 1387.690 1309.555 1387.705 ;
        RECT 1308.550 1387.390 1309.555 1387.690 ;
        RECT 1308.550 1387.010 1308.850 1387.390 ;
        RECT 1309.225 1387.375 1309.555 1387.390 ;
        RECT 1309.225 1387.010 1309.555 1387.025 ;
        RECT 1308.550 1386.710 1309.555 1387.010 ;
        RECT 1309.225 1386.695 1309.555 1386.710 ;
        RECT 1308.305 1248.970 1308.635 1248.985 ;
        RECT 1309.225 1248.970 1309.555 1248.985 ;
        RECT 1308.305 1248.670 1309.555 1248.970 ;
        RECT 1308.305 1248.655 1308.635 1248.670 ;
        RECT 1309.225 1248.655 1309.555 1248.670 ;
        RECT 1307.845 1097.330 1308.175 1097.345 ;
        RECT 1309.225 1097.330 1309.555 1097.345 ;
        RECT 1307.845 1097.030 1309.555 1097.330 ;
        RECT 1307.845 1097.015 1308.175 1097.030 ;
        RECT 1309.225 1097.015 1309.555 1097.030 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1269.210 17.580 1269.530 17.640 ;
        RECT 1269.210 17.440 1484.260 17.580 ;
        RECT 1269.210 17.380 1269.530 17.440 ;
        RECT 1484.120 17.240 1484.260 17.440 ;
        RECT 1492.770 17.240 1493.090 17.300 ;
        RECT 1484.120 17.100 1493.090 17.240 ;
        RECT 1492.770 17.040 1493.090 17.100 ;
      LAYER via ;
        RECT 1269.240 17.380 1269.500 17.640 ;
        RECT 1492.800 17.040 1493.060 17.300 ;
      LAYER met2 ;
        RECT 1493.710 1700.410 1493.990 1704.000 ;
        RECT 1492.860 1700.270 1493.990 1700.410 ;
        RECT 1269.240 17.350 1269.500 17.670 ;
        RECT 1269.300 2.400 1269.440 17.350 ;
        RECT 1492.860 17.330 1493.000 1700.270 ;
        RECT 1493.710 1700.000 1493.990 1700.270 ;
        RECT 1492.800 17.010 1493.060 17.330 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1289.910 1686.980 1290.230 1687.040 ;
        RECT 1498.750 1686.980 1499.070 1687.040 ;
        RECT 1289.910 1686.840 1499.070 1686.980 ;
        RECT 1289.910 1686.780 1290.230 1686.840 ;
        RECT 1498.750 1686.780 1499.070 1686.840 ;
        RECT 1287.150 20.640 1287.470 20.700 ;
        RECT 1289.910 20.640 1290.230 20.700 ;
        RECT 1287.150 20.500 1290.230 20.640 ;
        RECT 1287.150 20.440 1287.470 20.500 ;
        RECT 1289.910 20.440 1290.230 20.500 ;
      LAYER via ;
        RECT 1289.940 1686.780 1290.200 1687.040 ;
        RECT 1498.780 1686.780 1499.040 1687.040 ;
        RECT 1287.180 20.440 1287.440 20.700 ;
        RECT 1289.940 20.440 1290.200 20.700 ;
      LAYER met2 ;
        RECT 1498.770 1700.000 1499.050 1704.000 ;
        RECT 1498.840 1687.070 1498.980 1700.000 ;
        RECT 1289.940 1686.750 1290.200 1687.070 ;
        RECT 1498.780 1686.750 1499.040 1687.070 ;
        RECT 1290.000 20.730 1290.140 1686.750 ;
        RECT 1287.180 20.410 1287.440 20.730 ;
        RECT 1289.940 20.410 1290.200 20.730 ;
        RECT 1287.240 2.400 1287.380 20.410 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1310.610 1687.660 1310.930 1687.720 ;
        RECT 1503.350 1687.660 1503.670 1687.720 ;
        RECT 1310.610 1687.520 1503.670 1687.660 ;
        RECT 1310.610 1687.460 1310.930 1687.520 ;
        RECT 1503.350 1687.460 1503.670 1687.520 ;
        RECT 1305.090 18.260 1305.410 18.320 ;
        RECT 1310.610 18.260 1310.930 18.320 ;
        RECT 1305.090 18.120 1310.930 18.260 ;
        RECT 1305.090 18.060 1305.410 18.120 ;
        RECT 1310.610 18.060 1310.930 18.120 ;
      LAYER via ;
        RECT 1310.640 1687.460 1310.900 1687.720 ;
        RECT 1503.380 1687.460 1503.640 1687.720 ;
        RECT 1305.120 18.060 1305.380 18.320 ;
        RECT 1310.640 18.060 1310.900 18.320 ;
      LAYER met2 ;
        RECT 1503.370 1700.000 1503.650 1704.000 ;
        RECT 1503.440 1687.750 1503.580 1700.000 ;
        RECT 1310.640 1687.430 1310.900 1687.750 ;
        RECT 1503.380 1687.430 1503.640 1687.750 ;
        RECT 1310.700 18.350 1310.840 1687.430 ;
        RECT 1305.120 18.030 1305.380 18.350 ;
        RECT 1310.640 18.030 1310.900 18.350 ;
        RECT 1305.180 2.400 1305.320 18.030 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 0.300 ;
=======
      LAYER li1 ;
        RECT 1505.725 1400.885 1505.895 1448.995 ;
        RECT 1505.725 1304.325 1505.895 1352.435 ;
        RECT 1505.725 1207.765 1505.895 1255.875 ;
        RECT 1505.725 1159.485 1505.895 1207.255 ;
        RECT 1505.725 820.845 1505.895 862.495 ;
        RECT 1505.725 476.085 1505.895 524.195 ;
        RECT 1505.725 276.165 1505.895 324.275 ;
        RECT 1506.185 96.645 1506.355 144.755 ;
        RECT 1466.165 18.105 1466.335 20.995 ;
        RECT 1487.325 20.145 1487.495 20.995 ;
        RECT 1506.185 20.145 1506.355 48.195 ;
      LAYER mcon ;
        RECT 1505.725 1448.825 1505.895 1448.995 ;
        RECT 1505.725 1352.265 1505.895 1352.435 ;
        RECT 1505.725 1255.705 1505.895 1255.875 ;
        RECT 1505.725 1207.085 1505.895 1207.255 ;
        RECT 1505.725 862.325 1505.895 862.495 ;
        RECT 1505.725 524.025 1505.895 524.195 ;
        RECT 1505.725 324.105 1505.895 324.275 ;
        RECT 1506.185 144.585 1506.355 144.755 ;
        RECT 1506.185 48.025 1506.355 48.195 ;
        RECT 1466.165 20.825 1466.335 20.995 ;
        RECT 1487.325 20.825 1487.495 20.995 ;
      LAYER met1 ;
        RECT 1505.650 1546.360 1505.970 1546.620 ;
        RECT 1505.740 1545.940 1505.880 1546.360 ;
        RECT 1505.650 1545.680 1505.970 1545.940 ;
        RECT 1505.650 1448.980 1505.970 1449.040 ;
        RECT 1505.455 1448.840 1505.970 1448.980 ;
        RECT 1505.650 1448.780 1505.970 1448.840 ;
        RECT 1505.650 1401.040 1505.970 1401.100 ;
        RECT 1505.455 1400.900 1505.970 1401.040 ;
        RECT 1505.650 1400.840 1505.970 1400.900 ;
        RECT 1505.650 1352.420 1505.970 1352.480 ;
        RECT 1505.455 1352.280 1505.970 1352.420 ;
        RECT 1505.650 1352.220 1505.970 1352.280 ;
        RECT 1505.650 1304.480 1505.970 1304.540 ;
        RECT 1505.455 1304.340 1505.970 1304.480 ;
        RECT 1505.650 1304.280 1505.970 1304.340 ;
        RECT 1505.650 1255.860 1505.970 1255.920 ;
        RECT 1505.455 1255.720 1505.970 1255.860 ;
        RECT 1505.650 1255.660 1505.970 1255.720 ;
        RECT 1505.650 1207.920 1505.970 1207.980 ;
        RECT 1505.455 1207.780 1505.970 1207.920 ;
        RECT 1505.650 1207.720 1505.970 1207.780 ;
        RECT 1505.650 1207.240 1505.970 1207.300 ;
        RECT 1505.455 1207.100 1505.970 1207.240 ;
        RECT 1505.650 1207.040 1505.970 1207.100 ;
        RECT 1505.650 1159.640 1505.970 1159.700 ;
        RECT 1505.455 1159.500 1505.970 1159.640 ;
        RECT 1505.650 1159.440 1505.970 1159.500 ;
        RECT 1505.650 1062.540 1505.970 1062.800 ;
        RECT 1505.740 1062.400 1505.880 1062.540 ;
        RECT 1506.110 1062.400 1506.430 1062.460 ;
        RECT 1505.740 1062.260 1506.430 1062.400 ;
        RECT 1506.110 1062.200 1506.430 1062.260 ;
        RECT 1505.650 1007.660 1505.970 1007.720 ;
        RECT 1506.570 1007.660 1506.890 1007.720 ;
        RECT 1505.650 1007.520 1506.890 1007.660 ;
        RECT 1505.650 1007.460 1505.970 1007.520 ;
        RECT 1506.570 1007.460 1506.890 1007.520 ;
        RECT 1505.650 1000.520 1505.970 1000.580 ;
        RECT 1507.030 1000.520 1507.350 1000.580 ;
        RECT 1505.650 1000.380 1507.350 1000.520 ;
        RECT 1505.650 1000.320 1505.970 1000.380 ;
        RECT 1507.030 1000.320 1507.350 1000.380 ;
        RECT 1505.650 862.480 1505.970 862.540 ;
        RECT 1505.455 862.340 1505.970 862.480 ;
        RECT 1505.650 862.280 1505.970 862.340 ;
        RECT 1505.665 821.000 1505.955 821.045 ;
        RECT 1506.570 821.000 1506.890 821.060 ;
        RECT 1505.665 820.860 1506.890 821.000 ;
        RECT 1505.665 820.815 1505.955 820.860 ;
        RECT 1506.570 820.800 1506.890 820.860 ;
        RECT 1505.650 766.260 1505.970 766.320 ;
        RECT 1507.030 766.260 1507.350 766.320 ;
        RECT 1505.650 766.120 1507.350 766.260 ;
        RECT 1505.650 766.060 1505.970 766.120 ;
        RECT 1507.030 766.060 1507.350 766.120 ;
        RECT 1505.650 532.140 1505.970 532.400 ;
        RECT 1505.740 531.720 1505.880 532.140 ;
        RECT 1505.650 531.460 1505.970 531.720 ;
        RECT 1505.650 524.180 1505.970 524.240 ;
        RECT 1505.455 524.040 1505.970 524.180 ;
        RECT 1505.650 523.980 1505.970 524.040 ;
        RECT 1505.650 476.240 1505.970 476.300 ;
        RECT 1505.455 476.100 1505.970 476.240 ;
        RECT 1505.650 476.040 1505.970 476.100 ;
        RECT 1506.570 434.900 1506.890 435.160 ;
        RECT 1506.110 434.420 1506.430 434.480 ;
        RECT 1506.660 434.420 1506.800 434.900 ;
        RECT 1506.110 434.280 1506.800 434.420 ;
        RECT 1506.110 434.220 1506.430 434.280 ;
        RECT 1505.650 324.260 1505.970 324.320 ;
        RECT 1505.455 324.120 1505.970 324.260 ;
        RECT 1505.650 324.060 1505.970 324.120 ;
        RECT 1505.665 276.320 1505.955 276.365 ;
        RECT 1507.030 276.320 1507.350 276.380 ;
        RECT 1505.665 276.180 1507.350 276.320 ;
        RECT 1505.665 276.135 1505.955 276.180 ;
        RECT 1507.030 276.120 1507.350 276.180 ;
        RECT 1505.650 158.480 1505.970 158.740 ;
        RECT 1505.740 158.340 1505.880 158.480 ;
        RECT 1506.110 158.340 1506.430 158.400 ;
        RECT 1505.740 158.200 1506.430 158.340 ;
        RECT 1506.110 158.140 1506.430 158.200 ;
        RECT 1506.110 144.740 1506.430 144.800 ;
        RECT 1505.915 144.600 1506.430 144.740 ;
        RECT 1506.110 144.540 1506.430 144.600 ;
        RECT 1506.110 96.800 1506.430 96.860 ;
        RECT 1505.915 96.660 1506.430 96.800 ;
        RECT 1506.110 96.600 1506.430 96.660 ;
        RECT 1506.110 48.180 1506.430 48.240 ;
        RECT 1505.915 48.040 1506.430 48.180 ;
        RECT 1506.110 47.980 1506.430 48.040 ;
        RECT 1466.105 20.980 1466.395 21.025 ;
        RECT 1487.265 20.980 1487.555 21.025 ;
        RECT 1466.105 20.840 1487.555 20.980 ;
        RECT 1466.105 20.795 1466.395 20.840 ;
        RECT 1487.265 20.795 1487.555 20.840 ;
        RECT 1487.265 20.300 1487.555 20.345 ;
        RECT 1506.125 20.300 1506.415 20.345 ;
        RECT 1487.265 20.160 1506.415 20.300 ;
        RECT 1487.265 20.115 1487.555 20.160 ;
        RECT 1506.125 20.115 1506.415 20.160 ;
        RECT 1323.030 18.260 1323.350 18.320 ;
        RECT 1466.105 18.260 1466.395 18.305 ;
        RECT 1323.030 18.120 1466.395 18.260 ;
        RECT 1323.030 18.060 1323.350 18.120 ;
        RECT 1466.105 18.075 1466.395 18.120 ;
      LAYER via ;
        RECT 1505.680 1546.360 1505.940 1546.620 ;
        RECT 1505.680 1545.680 1505.940 1545.940 ;
        RECT 1505.680 1448.780 1505.940 1449.040 ;
        RECT 1505.680 1400.840 1505.940 1401.100 ;
        RECT 1505.680 1352.220 1505.940 1352.480 ;
        RECT 1505.680 1304.280 1505.940 1304.540 ;
        RECT 1505.680 1255.660 1505.940 1255.920 ;
        RECT 1505.680 1207.720 1505.940 1207.980 ;
        RECT 1505.680 1207.040 1505.940 1207.300 ;
        RECT 1505.680 1159.440 1505.940 1159.700 ;
        RECT 1505.680 1062.540 1505.940 1062.800 ;
        RECT 1506.140 1062.200 1506.400 1062.460 ;
        RECT 1505.680 1007.460 1505.940 1007.720 ;
        RECT 1506.600 1007.460 1506.860 1007.720 ;
        RECT 1505.680 1000.320 1505.940 1000.580 ;
        RECT 1507.060 1000.320 1507.320 1000.580 ;
        RECT 1505.680 862.280 1505.940 862.540 ;
        RECT 1506.600 820.800 1506.860 821.060 ;
        RECT 1505.680 766.060 1505.940 766.320 ;
        RECT 1507.060 766.060 1507.320 766.320 ;
        RECT 1505.680 532.140 1505.940 532.400 ;
        RECT 1505.680 531.460 1505.940 531.720 ;
        RECT 1505.680 523.980 1505.940 524.240 ;
        RECT 1505.680 476.040 1505.940 476.300 ;
        RECT 1506.600 434.900 1506.860 435.160 ;
        RECT 1506.140 434.220 1506.400 434.480 ;
        RECT 1505.680 324.060 1505.940 324.320 ;
        RECT 1507.060 276.120 1507.320 276.380 ;
        RECT 1505.680 158.480 1505.940 158.740 ;
        RECT 1506.140 158.140 1506.400 158.400 ;
        RECT 1506.140 144.540 1506.400 144.800 ;
        RECT 1506.140 96.600 1506.400 96.860 ;
        RECT 1506.140 47.980 1506.400 48.240 ;
        RECT 1323.060 18.060 1323.320 18.320 ;
      LAYER met2 ;
        RECT 1508.430 1700.410 1508.710 1704.000 ;
        RECT 1507.580 1700.270 1508.710 1700.410 ;
        RECT 1507.580 1678.140 1507.720 1700.270 ;
        RECT 1508.430 1700.000 1508.710 1700.270 ;
        RECT 1505.740 1678.000 1507.720 1678.140 ;
        RECT 1505.740 1546.650 1505.880 1678.000 ;
        RECT 1505.680 1546.330 1505.940 1546.650 ;
        RECT 1505.680 1545.650 1505.940 1545.970 ;
        RECT 1505.740 1449.070 1505.880 1545.650 ;
        RECT 1505.680 1448.750 1505.940 1449.070 ;
        RECT 1505.680 1400.810 1505.940 1401.130 ;
        RECT 1505.740 1352.510 1505.880 1400.810 ;
        RECT 1505.680 1352.190 1505.940 1352.510 ;
        RECT 1505.680 1304.250 1505.940 1304.570 ;
        RECT 1505.740 1255.950 1505.880 1304.250 ;
        RECT 1505.680 1255.630 1505.940 1255.950 ;
        RECT 1505.680 1207.690 1505.940 1208.010 ;
        RECT 1505.740 1207.330 1505.880 1207.690 ;
        RECT 1505.680 1207.010 1505.940 1207.330 ;
        RECT 1505.680 1159.410 1505.940 1159.730 ;
        RECT 1505.740 1062.830 1505.880 1159.410 ;
        RECT 1505.680 1062.510 1505.940 1062.830 ;
        RECT 1506.140 1062.170 1506.400 1062.490 ;
        RECT 1506.200 1014.970 1506.340 1062.170 ;
        RECT 1506.200 1014.830 1506.800 1014.970 ;
        RECT 1506.660 1007.750 1506.800 1014.830 ;
        RECT 1505.680 1007.430 1505.940 1007.750 ;
        RECT 1506.600 1007.430 1506.860 1007.750 ;
        RECT 1505.740 1000.610 1505.880 1007.430 ;
        RECT 1505.680 1000.290 1505.940 1000.610 ;
        RECT 1507.060 1000.290 1507.320 1000.610 ;
        RECT 1507.120 952.525 1507.260 1000.290 ;
        RECT 1506.130 952.155 1506.410 952.525 ;
        RECT 1507.050 952.155 1507.330 952.525 ;
        RECT 1506.200 931.330 1506.340 952.155 ;
        RECT 1506.200 931.190 1506.800 931.330 ;
        RECT 1506.660 884.525 1506.800 931.190 ;
        RECT 1506.590 884.155 1506.870 884.525 ;
        RECT 1505.670 862.395 1505.950 862.765 ;
        RECT 1505.680 862.250 1505.940 862.395 ;
        RECT 1506.600 820.770 1506.860 821.090 ;
        RECT 1506.660 814.370 1506.800 820.770 ;
        RECT 1506.660 814.230 1507.260 814.370 ;
        RECT 1507.120 766.350 1507.260 814.230 ;
        RECT 1505.680 766.030 1505.940 766.350 ;
        RECT 1507.060 766.030 1507.320 766.350 ;
        RECT 1505.740 532.430 1505.880 766.030 ;
        RECT 1505.680 532.110 1505.940 532.430 ;
        RECT 1505.680 531.430 1505.940 531.750 ;
        RECT 1505.740 524.270 1505.880 531.430 ;
        RECT 1505.680 523.950 1505.940 524.270 ;
        RECT 1505.680 476.010 1505.940 476.330 ;
        RECT 1505.740 475.845 1505.880 476.010 ;
        RECT 1505.670 475.475 1505.950 475.845 ;
        RECT 1506.590 475.475 1506.870 475.845 ;
        RECT 1506.660 435.190 1506.800 475.475 ;
        RECT 1506.600 434.870 1506.860 435.190 ;
        RECT 1506.140 434.190 1506.400 434.510 ;
        RECT 1506.200 427.565 1506.340 434.190 ;
        RECT 1506.130 427.195 1506.410 427.565 ;
        RECT 1505.670 379.595 1505.950 379.965 ;
        RECT 1505.740 324.350 1505.880 379.595 ;
        RECT 1505.680 324.030 1505.940 324.350 ;
        RECT 1507.060 276.090 1507.320 276.410 ;
        RECT 1507.120 254.730 1507.260 276.090 ;
        RECT 1506.200 254.590 1507.260 254.730 ;
        RECT 1506.200 206.960 1506.340 254.590 ;
        RECT 1505.740 206.820 1506.340 206.960 ;
        RECT 1505.740 158.770 1505.880 206.820 ;
        RECT 1505.680 158.450 1505.940 158.770 ;
        RECT 1506.140 158.110 1506.400 158.430 ;
        RECT 1506.200 144.830 1506.340 158.110 ;
        RECT 1506.140 144.510 1506.400 144.830 ;
        RECT 1506.140 96.570 1506.400 96.890 ;
        RECT 1506.200 48.270 1506.340 96.570 ;
        RECT 1506.140 47.950 1506.400 48.270 ;
        RECT 1323.060 18.030 1323.320 18.350 ;
        RECT 1323.120 2.400 1323.260 18.030 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 1506.130 952.200 1506.410 952.480 ;
        RECT 1507.050 952.200 1507.330 952.480 ;
        RECT 1506.590 884.200 1506.870 884.480 ;
        RECT 1505.670 862.440 1505.950 862.720 ;
        RECT 1505.670 475.520 1505.950 475.800 ;
        RECT 1506.590 475.520 1506.870 475.800 ;
        RECT 1506.130 427.240 1506.410 427.520 ;
        RECT 1505.670 379.640 1505.950 379.920 ;
      LAYER met3 ;
        RECT 1506.105 952.490 1506.435 952.505 ;
        RECT 1507.025 952.490 1507.355 952.505 ;
        RECT 1506.105 952.190 1507.355 952.490 ;
        RECT 1506.105 952.175 1506.435 952.190 ;
        RECT 1507.025 952.175 1507.355 952.190 ;
        RECT 1505.390 884.490 1505.770 884.500 ;
        RECT 1506.565 884.490 1506.895 884.505 ;
        RECT 1505.390 884.190 1506.895 884.490 ;
        RECT 1505.390 884.180 1505.770 884.190 ;
        RECT 1506.565 884.175 1506.895 884.190 ;
        RECT 1505.645 862.740 1505.975 862.745 ;
        RECT 1505.390 862.730 1505.975 862.740 ;
        RECT 1505.390 862.430 1506.200 862.730 ;
        RECT 1505.390 862.420 1505.975 862.430 ;
        RECT 1505.645 862.415 1505.975 862.420 ;
        RECT 1505.645 475.810 1505.975 475.825 ;
        RECT 1506.565 475.810 1506.895 475.825 ;
        RECT 1505.645 475.510 1506.895 475.810 ;
        RECT 1505.645 475.495 1505.975 475.510 ;
        RECT 1506.565 475.495 1506.895 475.510 ;
        RECT 1505.390 427.530 1505.770 427.540 ;
        RECT 1506.105 427.530 1506.435 427.545 ;
        RECT 1505.390 427.230 1506.435 427.530 ;
        RECT 1505.390 427.220 1505.770 427.230 ;
        RECT 1506.105 427.215 1506.435 427.230 ;
        RECT 1505.645 379.940 1505.975 379.945 ;
        RECT 1505.390 379.930 1505.975 379.940 ;
        RECT 1505.390 379.630 1506.200 379.930 ;
        RECT 1505.390 379.620 1505.975 379.630 ;
        RECT 1505.645 379.615 1505.975 379.620 ;
      LAYER via3 ;
        RECT 1505.420 884.180 1505.740 884.500 ;
        RECT 1505.420 862.420 1505.740 862.740 ;
        RECT 1505.420 427.220 1505.740 427.540 ;
        RECT 1505.420 379.620 1505.740 379.940 ;
      LAYER met4 ;
        RECT 1505.415 884.175 1505.745 884.505 ;
        RECT 1505.430 862.745 1505.730 884.175 ;
        RECT 1505.415 862.415 1505.745 862.745 ;
        RECT 1505.415 427.215 1505.745 427.545 ;
        RECT 1505.430 379.945 1505.730 427.215 ;
        RECT 1505.415 379.615 1505.745 379.945 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 0.300 ;
=======
      LAYER li1 ;
        RECT 1390.265 1686.485 1390.435 1688.695 ;
      LAYER mcon ;
        RECT 1390.265 1688.525 1390.435 1688.695 ;
      LAYER met1 ;
        RECT 1513.010 1689.020 1513.330 1689.080 ;
        RECT 1486.880 1688.880 1513.330 1689.020 ;
        RECT 1390.205 1688.680 1390.495 1688.725 ;
        RECT 1486.880 1688.680 1487.020 1688.880 ;
        RECT 1513.010 1688.820 1513.330 1688.880 ;
        RECT 1390.205 1688.540 1487.020 1688.680 ;
        RECT 1390.205 1688.495 1390.495 1688.540 ;
        RECT 1345.110 1686.640 1345.430 1686.700 ;
        RECT 1390.205 1686.640 1390.495 1686.685 ;
        RECT 1345.110 1686.500 1390.495 1686.640 ;
        RECT 1345.110 1686.440 1345.430 1686.500 ;
        RECT 1390.205 1686.455 1390.495 1686.500 ;
        RECT 1345.110 1139.720 1345.430 1139.980 ;
        RECT 1345.200 1138.960 1345.340 1139.720 ;
        RECT 1345.110 1138.700 1345.430 1138.960 ;
        RECT 1340.510 20.640 1340.830 20.700 ;
        RECT 1345.110 20.640 1345.430 20.700 ;
        RECT 1340.510 20.500 1345.430 20.640 ;
        RECT 1340.510 20.440 1340.830 20.500 ;
        RECT 1345.110 20.440 1345.430 20.500 ;
      LAYER via ;
        RECT 1513.040 1688.820 1513.300 1689.080 ;
        RECT 1345.140 1686.440 1345.400 1686.700 ;
        RECT 1345.140 1139.720 1345.400 1139.980 ;
        RECT 1345.140 1138.700 1345.400 1138.960 ;
        RECT 1340.540 20.440 1340.800 20.700 ;
        RECT 1345.140 20.440 1345.400 20.700 ;
      LAYER met2 ;
        RECT 1513.030 1700.000 1513.310 1704.000 ;
        RECT 1513.100 1689.110 1513.240 1700.000 ;
        RECT 1513.040 1688.790 1513.300 1689.110 ;
        RECT 1345.140 1686.410 1345.400 1686.730 ;
        RECT 1345.200 1140.010 1345.340 1686.410 ;
        RECT 1345.140 1139.690 1345.400 1140.010 ;
        RECT 1345.140 1138.670 1345.400 1138.990 ;
        RECT 1345.200 20.730 1345.340 1138.670 ;
        RECT 1340.540 20.410 1340.800 20.730 ;
        RECT 1345.140 20.410 1345.400 20.730 ;
        RECT 1340.600 2.400 1340.740 20.410 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 0.300 ;
=======
      LAYER met1 ;
        RECT 698.350 47.840 698.670 47.900 ;
        RECT 1339.130 47.840 1339.450 47.900 ;
        RECT 698.350 47.700 1339.450 47.840 ;
        RECT 698.350 47.640 698.670 47.700 ;
        RECT 1339.130 47.640 1339.450 47.700 ;
      LAYER via ;
        RECT 698.380 47.640 698.640 47.900 ;
        RECT 1339.160 47.640 1339.420 47.900 ;
      LAYER met2 ;
        RECT 1339.150 1700.000 1339.430 1704.000 ;
        RECT 1339.220 47.930 1339.360 1700.000 ;
        RECT 698.380 47.610 698.640 47.930 ;
        RECT 1339.160 47.610 1339.420 47.930 ;
        RECT 698.440 2.400 698.580 47.610 ;
        RECT 698.230 -4.800 698.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 0.300 ;
=======
      LAYER li1 ;
        RECT 1510.785 15.725 1510.955 19.635 ;
      LAYER mcon ;
        RECT 1510.785 19.465 1510.955 19.635 ;
      LAYER met1 ;
        RECT 1487.250 19.620 1487.570 19.680 ;
        RECT 1510.725 19.620 1511.015 19.665 ;
        RECT 1487.250 19.480 1511.015 19.620 ;
        RECT 1487.250 19.420 1487.570 19.480 ;
        RECT 1510.725 19.435 1511.015 19.480 ;
        RECT 1358.450 18.600 1358.770 18.660 ;
        RECT 1485.410 18.600 1485.730 18.660 ;
        RECT 1358.450 18.460 1485.730 18.600 ;
        RECT 1358.450 18.400 1358.770 18.460 ;
        RECT 1485.410 18.400 1485.730 18.460 ;
        RECT 1510.725 15.880 1511.015 15.925 ;
        RECT 1518.530 15.880 1518.850 15.940 ;
        RECT 1510.725 15.740 1518.850 15.880 ;
        RECT 1510.725 15.695 1511.015 15.740 ;
        RECT 1518.530 15.680 1518.850 15.740 ;
      LAYER via ;
        RECT 1487.280 19.420 1487.540 19.680 ;
        RECT 1358.480 18.400 1358.740 18.660 ;
        RECT 1485.440 18.400 1485.700 18.660 ;
        RECT 1518.560 15.680 1518.820 15.940 ;
      LAYER met2 ;
        RECT 1518.090 1700.410 1518.370 1704.000 ;
        RECT 1518.090 1700.270 1519.220 1700.410 ;
        RECT 1518.090 1700.000 1518.370 1700.270 ;
        RECT 1487.280 19.390 1487.540 19.710 ;
        RECT 1487.340 18.770 1487.480 19.390 ;
        RECT 1519.080 18.770 1519.220 1700.270 ;
        RECT 1485.500 18.690 1487.480 18.770 ;
        RECT 1358.480 18.370 1358.740 18.690 ;
        RECT 1485.440 18.630 1487.480 18.690 ;
        RECT 1518.620 18.630 1519.220 18.770 ;
        RECT 1485.440 18.370 1485.700 18.630 ;
        RECT 1358.540 2.400 1358.680 18.370 ;
        RECT 1518.620 15.970 1518.760 18.630 ;
        RECT 1518.560 15.650 1518.820 15.970 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1513.950 1593.440 1514.230 1593.720 ;
        RECT 1514.870 1593.440 1515.150 1593.720 ;
        RECT 1513.490 1338.440 1513.770 1338.720 ;
        RECT 1513.030 1289.480 1513.310 1289.760 ;
        RECT 1513.030 1241.880 1513.310 1242.160 ;
        RECT 1513.950 1241.880 1514.230 1242.160 ;
        RECT 1513.490 1048.760 1513.770 1049.040 ;
        RECT 1514.870 1048.760 1515.150 1049.040 ;
        RECT 1513.490 965.800 1513.770 966.080 ;
        RECT 1515.330 965.800 1515.610 966.080 ;
        RECT 1513.950 917.520 1514.230 917.800 ;
        RECT 1515.330 917.520 1515.610 917.800 ;
        RECT 1513.950 434.040 1514.230 434.320 ;
        RECT 1513.490 386.440 1513.770 386.720 ;
        RECT 1513.030 338.840 1513.310 339.120 ;
        RECT 1513.950 338.160 1514.230 338.440 ;
        RECT 1513.950 241.600 1514.230 241.880 ;
        RECT 1514.870 241.600 1515.150 241.880 ;
      LAYER met3 ;
        RECT 1513.925 1593.730 1514.255 1593.745 ;
        RECT 1514.845 1593.730 1515.175 1593.745 ;
        RECT 1513.925 1593.430 1515.175 1593.730 ;
        RECT 1513.925 1593.415 1514.255 1593.430 ;
        RECT 1514.845 1593.415 1515.175 1593.430 ;
        RECT 1513.465 1338.740 1513.795 1338.745 ;
        RECT 1513.465 1338.730 1514.050 1338.740 ;
        RECT 1513.465 1338.430 1514.250 1338.730 ;
        RECT 1513.465 1338.420 1514.050 1338.430 ;
        RECT 1513.465 1338.415 1513.795 1338.420 ;
        RECT 1513.670 1290.140 1514.050 1290.460 ;
        RECT 1513.005 1289.770 1513.335 1289.785 ;
        RECT 1513.710 1289.770 1514.010 1290.140 ;
        RECT 1513.005 1289.470 1514.010 1289.770 ;
        RECT 1513.005 1289.455 1513.335 1289.470 ;
        RECT 1513.005 1242.170 1513.335 1242.185 ;
        RECT 1513.925 1242.170 1514.255 1242.185 ;
        RECT 1513.005 1241.870 1514.255 1242.170 ;
        RECT 1513.005 1241.855 1513.335 1241.870 ;
        RECT 1513.925 1241.855 1514.255 1241.870 ;
        RECT 1513.465 1049.050 1513.795 1049.065 ;
        RECT 1514.845 1049.050 1515.175 1049.065 ;
        RECT 1513.465 1048.750 1515.175 1049.050 ;
        RECT 1513.465 1048.735 1513.795 1048.750 ;
        RECT 1514.845 1048.735 1515.175 1048.750 ;
        RECT 1513.465 966.090 1513.795 966.105 ;
        RECT 1515.305 966.090 1515.635 966.105 ;
        RECT 1513.465 965.790 1515.635 966.090 ;
        RECT 1513.465 965.775 1513.795 965.790 ;
        RECT 1515.305 965.775 1515.635 965.790 ;
        RECT 1513.925 917.810 1514.255 917.825 ;
        RECT 1515.305 917.810 1515.635 917.825 ;
        RECT 1513.925 917.510 1515.635 917.810 ;
        RECT 1513.925 917.495 1514.255 917.510 ;
        RECT 1515.305 917.495 1515.635 917.510 ;
        RECT 1513.925 434.340 1514.255 434.345 ;
        RECT 1513.670 434.330 1514.255 434.340 ;
        RECT 1513.470 434.030 1514.255 434.330 ;
        RECT 1513.670 434.020 1514.255 434.030 ;
        RECT 1513.925 434.015 1514.255 434.020 ;
        RECT 1513.465 386.740 1513.795 386.745 ;
        RECT 1513.465 386.730 1514.050 386.740 ;
        RECT 1513.240 386.430 1514.050 386.730 ;
        RECT 1513.465 386.420 1514.050 386.430 ;
        RECT 1513.465 386.415 1513.795 386.420 ;
        RECT 1513.005 339.130 1513.335 339.145 ;
        RECT 1513.005 338.830 1514.930 339.130 ;
        RECT 1513.005 338.815 1513.335 338.830 ;
        RECT 1513.925 338.450 1514.255 338.465 ;
        RECT 1514.630 338.450 1514.930 338.830 ;
        RECT 1513.925 338.150 1514.930 338.450 ;
        RECT 1513.925 338.135 1514.255 338.150 ;
        RECT 1513.925 241.890 1514.255 241.905 ;
        RECT 1514.845 241.890 1515.175 241.905 ;
        RECT 1513.925 241.590 1515.175 241.890 ;
        RECT 1513.925 241.575 1514.255 241.590 ;
        RECT 1514.845 241.575 1515.175 241.590 ;
      LAYER via3 ;
        RECT 1513.700 1338.420 1514.020 1338.740 ;
        RECT 1513.700 1290.140 1514.020 1290.460 ;
        RECT 1513.700 434.020 1514.020 434.340 ;
        RECT 1513.700 386.420 1514.020 386.740 ;
      LAYER met4 ;
        RECT 1513.695 1338.415 1514.025 1338.745 ;
        RECT 1513.710 1290.465 1514.010 1338.415 ;
        RECT 1513.695 1290.135 1514.025 1290.465 ;
        RECT 1513.695 434.015 1514.025 434.345 ;
        RECT 1513.710 386.745 1514.010 434.015 ;
        RECT 1513.695 386.415 1514.025 386.745 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 0.300 ;
=======
      LAYER met1 ;
        RECT 1518.530 1678.140 1518.850 1678.200 ;
        RECT 1521.750 1678.140 1522.070 1678.200 ;
        RECT 1518.530 1678.000 1522.070 1678.140 ;
        RECT 1518.530 1677.940 1518.850 1678.000 ;
        RECT 1521.750 1677.940 1522.070 1678.000 ;
        RECT 1518.530 20.300 1518.850 20.360 ;
        RECT 1506.660 20.160 1518.850 20.300 ;
        RECT 1506.660 19.960 1506.800 20.160 ;
        RECT 1518.530 20.100 1518.850 20.160 ;
        RECT 1486.880 19.820 1506.800 19.960 ;
        RECT 1376.390 19.620 1376.710 19.680 ;
        RECT 1486.880 19.620 1487.020 19.820 ;
        RECT 1376.390 19.480 1487.020 19.620 ;
        RECT 1376.390 19.420 1376.710 19.480 ;
      LAYER via ;
        RECT 1518.560 1677.940 1518.820 1678.200 ;
        RECT 1521.780 1677.940 1522.040 1678.200 ;
        RECT 1518.560 20.100 1518.820 20.360 ;
        RECT 1376.420 19.420 1376.680 19.680 ;
      LAYER met2 ;
        RECT 1522.690 1700.410 1522.970 1704.000 ;
        RECT 1521.840 1700.270 1522.970 1700.410 ;
        RECT 1521.840 1678.230 1521.980 1700.270 ;
        RECT 1522.690 1700.000 1522.970 1700.270 ;
        RECT 1518.560 1677.910 1518.820 1678.230 ;
        RECT 1521.780 1677.910 1522.040 1678.230 ;
        RECT 1518.620 20.390 1518.760 1677.910 ;
        RECT 1518.560 20.070 1518.820 20.390 ;
        RECT 1376.420 19.390 1376.680 19.710 ;
        RECT 1376.480 2.400 1376.620 19.390 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 0.300 ;
=======
      LAYER li1 ;
        RECT 1438.565 1686.485 1438.735 1689.035 ;
        RECT 1481.805 1688.865 1481.975 1690.395 ;
      LAYER mcon ;
        RECT 1481.805 1690.225 1481.975 1690.395 ;
        RECT 1438.565 1688.865 1438.735 1689.035 ;
      LAYER met1 ;
        RECT 1481.745 1690.380 1482.035 1690.425 ;
        RECT 1527.730 1690.380 1528.050 1690.440 ;
        RECT 1481.745 1690.240 1528.050 1690.380 ;
        RECT 1481.745 1690.195 1482.035 1690.240 ;
        RECT 1527.730 1690.180 1528.050 1690.240 ;
        RECT 1438.505 1689.020 1438.795 1689.065 ;
        RECT 1481.745 1689.020 1482.035 1689.065 ;
        RECT 1438.505 1688.880 1482.035 1689.020 ;
        RECT 1438.505 1688.835 1438.795 1688.880 ;
        RECT 1481.745 1688.835 1482.035 1688.880 ;
        RECT 1400.310 1686.640 1400.630 1686.700 ;
        RECT 1438.505 1686.640 1438.795 1686.685 ;
        RECT 1400.310 1686.500 1438.795 1686.640 ;
        RECT 1400.310 1686.440 1400.630 1686.500 ;
        RECT 1438.505 1686.455 1438.795 1686.500 ;
        RECT 1394.330 20.640 1394.650 20.700 ;
        RECT 1400.310 20.640 1400.630 20.700 ;
        RECT 1394.330 20.500 1400.630 20.640 ;
        RECT 1394.330 20.440 1394.650 20.500 ;
        RECT 1400.310 20.440 1400.630 20.500 ;
      LAYER via ;
        RECT 1527.760 1690.180 1528.020 1690.440 ;
        RECT 1400.340 1686.440 1400.600 1686.700 ;
        RECT 1394.360 20.440 1394.620 20.700 ;
        RECT 1400.340 20.440 1400.600 20.700 ;
      LAYER met2 ;
        RECT 1527.750 1700.000 1528.030 1704.000 ;
        RECT 1527.820 1690.470 1527.960 1700.000 ;
        RECT 1527.760 1690.150 1528.020 1690.470 ;
        RECT 1400.340 1686.410 1400.600 1686.730 ;
        RECT 1400.400 20.730 1400.540 1686.410 ;
        RECT 1394.360 20.410 1394.620 20.730 ;
        RECT 1400.340 20.410 1400.600 20.730 ;
        RECT 1394.420 2.400 1394.560 20.410 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 0.300 ;
=======
      LAYER li1 ;
        RECT 1486.405 18.785 1486.575 19.975 ;
      LAYER mcon ;
        RECT 1486.405 19.805 1486.575 19.975 ;
      LAYER met1 ;
        RECT 1412.270 19.960 1412.590 20.020 ;
        RECT 1486.345 19.960 1486.635 20.005 ;
        RECT 1412.270 19.820 1486.635 19.960 ;
        RECT 1412.270 19.760 1412.590 19.820 ;
        RECT 1486.345 19.775 1486.635 19.820 ;
        RECT 1486.345 18.940 1486.635 18.985 ;
        RECT 1532.330 18.940 1532.650 19.000 ;
        RECT 1486.345 18.800 1532.650 18.940 ;
        RECT 1486.345 18.755 1486.635 18.800 ;
        RECT 1532.330 18.740 1532.650 18.800 ;
      LAYER via ;
        RECT 1412.300 19.760 1412.560 20.020 ;
        RECT 1532.360 18.740 1532.620 19.000 ;
      LAYER met2 ;
        RECT 1532.350 1700.000 1532.630 1704.000 ;
        RECT 1412.300 19.730 1412.560 20.050 ;
        RECT 1412.360 2.400 1412.500 19.730 ;
        RECT 1532.420 19.030 1532.560 1700.000 ;
        RECT 1532.360 18.710 1532.620 19.030 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 0.300 ;
=======
      LAYER li1 ;
        RECT 1535.165 1497.445 1535.335 1545.555 ;
        RECT 1534.245 1400.885 1534.415 1466.335 ;
        RECT 1534.245 1304.325 1534.415 1352.435 ;
        RECT 1534.245 1207.425 1534.415 1255.875 ;
        RECT 1533.325 386.325 1533.495 434.775 ;
        RECT 1533.325 351.305 1533.495 372.555 ;
        RECT 1534.245 241.485 1534.415 289.595 ;
        RECT 1534.245 120.445 1534.415 186.235 ;
      LAYER mcon ;
        RECT 1535.165 1545.385 1535.335 1545.555 ;
        RECT 1534.245 1466.165 1534.415 1466.335 ;
        RECT 1534.245 1352.265 1534.415 1352.435 ;
        RECT 1534.245 1255.705 1534.415 1255.875 ;
        RECT 1533.325 434.605 1533.495 434.775 ;
        RECT 1533.325 372.385 1533.495 372.555 ;
        RECT 1534.245 289.425 1534.415 289.595 ;
        RECT 1534.245 186.065 1534.415 186.235 ;
      LAYER met1 ;
        RECT 1534.630 1663.180 1534.950 1663.240 ;
        RECT 1536.930 1663.180 1537.250 1663.240 ;
        RECT 1534.630 1663.040 1537.250 1663.180 ;
        RECT 1534.630 1662.980 1534.950 1663.040 ;
        RECT 1536.930 1662.980 1537.250 1663.040 ;
        RECT 1534.170 1594.160 1534.490 1594.220 ;
        RECT 1534.630 1594.160 1534.950 1594.220 ;
        RECT 1534.170 1594.020 1534.950 1594.160 ;
        RECT 1534.170 1593.960 1534.490 1594.020 ;
        RECT 1534.630 1593.960 1534.950 1594.020 ;
        RECT 1535.090 1545.540 1535.410 1545.600 ;
        RECT 1534.895 1545.400 1535.410 1545.540 ;
        RECT 1535.090 1545.340 1535.410 1545.400 ;
        RECT 1535.105 1497.600 1535.395 1497.645 ;
        RECT 1535.550 1497.600 1535.870 1497.660 ;
        RECT 1535.105 1497.460 1535.870 1497.600 ;
        RECT 1535.105 1497.415 1535.395 1497.460 ;
        RECT 1535.550 1497.400 1535.870 1497.460 ;
        RECT 1534.185 1466.320 1534.475 1466.365 ;
        RECT 1535.550 1466.320 1535.870 1466.380 ;
        RECT 1534.185 1466.180 1535.870 1466.320 ;
        RECT 1534.185 1466.135 1534.475 1466.180 ;
        RECT 1535.550 1466.120 1535.870 1466.180 ;
        RECT 1534.170 1401.040 1534.490 1401.100 ;
        RECT 1533.975 1400.900 1534.490 1401.040 ;
        RECT 1534.170 1400.840 1534.490 1400.900 ;
        RECT 1533.710 1366.020 1534.030 1366.080 ;
        RECT 1534.630 1366.020 1534.950 1366.080 ;
        RECT 1533.710 1365.880 1534.950 1366.020 ;
        RECT 1533.710 1365.820 1534.030 1365.880 ;
        RECT 1534.630 1365.820 1534.950 1365.880 ;
        RECT 1534.185 1352.420 1534.475 1352.465 ;
        RECT 1534.630 1352.420 1534.950 1352.480 ;
        RECT 1534.185 1352.280 1534.950 1352.420 ;
        RECT 1534.185 1352.235 1534.475 1352.280 ;
        RECT 1534.630 1352.220 1534.950 1352.280 ;
        RECT 1534.170 1304.480 1534.490 1304.540 ;
        RECT 1533.975 1304.340 1534.490 1304.480 ;
        RECT 1534.170 1304.280 1534.490 1304.340 ;
        RECT 1533.710 1269.460 1534.030 1269.520 ;
        RECT 1534.630 1269.460 1534.950 1269.520 ;
        RECT 1533.710 1269.320 1534.950 1269.460 ;
        RECT 1533.710 1269.260 1534.030 1269.320 ;
        RECT 1534.630 1269.260 1534.950 1269.320 ;
        RECT 1534.185 1255.860 1534.475 1255.905 ;
        RECT 1534.630 1255.860 1534.950 1255.920 ;
        RECT 1534.185 1255.720 1534.950 1255.860 ;
        RECT 1534.185 1255.675 1534.475 1255.720 ;
        RECT 1534.630 1255.660 1534.950 1255.720 ;
        RECT 1534.170 1207.580 1534.490 1207.640 ;
        RECT 1533.975 1207.440 1534.490 1207.580 ;
        RECT 1534.170 1207.380 1534.490 1207.440 ;
        RECT 1533.710 1076.340 1534.030 1076.400 ;
        RECT 1534.630 1076.340 1534.950 1076.400 ;
        RECT 1533.710 1076.200 1534.950 1076.340 ;
        RECT 1533.710 1076.140 1534.030 1076.200 ;
        RECT 1534.630 1076.140 1534.950 1076.200 ;
        RECT 1533.710 1014.460 1534.030 1014.520 ;
        RECT 1534.170 1014.460 1534.490 1014.520 ;
        RECT 1533.710 1014.320 1534.490 1014.460 ;
        RECT 1533.710 1014.260 1534.030 1014.320 ;
        RECT 1534.170 1014.260 1534.490 1014.320 ;
        RECT 1534.170 821.000 1534.490 821.060 ;
        RECT 1534.630 821.000 1534.950 821.060 ;
        RECT 1534.170 820.860 1534.950 821.000 ;
        RECT 1534.170 820.800 1534.490 820.860 ;
        RECT 1534.630 820.800 1534.950 820.860 ;
        RECT 1533.265 434.760 1533.555 434.805 ;
        RECT 1533.710 434.760 1534.030 434.820 ;
        RECT 1533.265 434.620 1534.030 434.760 ;
        RECT 1533.265 434.575 1533.555 434.620 ;
        RECT 1533.710 434.560 1534.030 434.620 ;
        RECT 1533.250 386.480 1533.570 386.540 ;
        RECT 1533.055 386.340 1533.570 386.480 ;
        RECT 1533.250 386.280 1533.570 386.340 ;
        RECT 1533.250 372.540 1533.570 372.600 ;
        RECT 1533.055 372.400 1533.570 372.540 ;
        RECT 1533.250 372.340 1533.570 372.400 ;
        RECT 1533.265 351.460 1533.555 351.505 ;
        RECT 1533.710 351.460 1534.030 351.520 ;
        RECT 1533.265 351.320 1534.030 351.460 ;
        RECT 1533.265 351.275 1533.555 351.320 ;
        RECT 1533.710 351.260 1534.030 351.320 ;
        RECT 1533.710 303.520 1534.030 303.580 ;
        RECT 1534.630 303.520 1534.950 303.580 ;
        RECT 1533.710 303.380 1534.950 303.520 ;
        RECT 1533.710 303.320 1534.030 303.380 ;
        RECT 1534.630 303.320 1534.950 303.380 ;
        RECT 1534.185 289.580 1534.475 289.625 ;
        RECT 1534.630 289.580 1534.950 289.640 ;
        RECT 1534.185 289.440 1534.950 289.580 ;
        RECT 1534.185 289.395 1534.475 289.440 ;
        RECT 1534.630 289.380 1534.950 289.440 ;
        RECT 1534.170 241.640 1534.490 241.700 ;
        RECT 1533.975 241.500 1534.490 241.640 ;
        RECT 1534.170 241.440 1534.490 241.500 ;
        RECT 1534.170 234.500 1534.490 234.560 ;
        RECT 1535.090 234.500 1535.410 234.560 ;
        RECT 1534.170 234.360 1535.410 234.500 ;
        RECT 1534.170 234.300 1534.490 234.360 ;
        RECT 1535.090 234.300 1535.410 234.360 ;
        RECT 1534.185 186.220 1534.475 186.265 ;
        RECT 1535.090 186.220 1535.410 186.280 ;
        RECT 1534.185 186.080 1535.410 186.220 ;
        RECT 1534.185 186.035 1534.475 186.080 ;
        RECT 1535.090 186.020 1535.410 186.080 ;
        RECT 1534.185 120.600 1534.475 120.645 ;
        RECT 1534.630 120.600 1534.950 120.660 ;
        RECT 1534.185 120.460 1534.950 120.600 ;
        RECT 1534.185 120.415 1534.475 120.460 ;
        RECT 1534.630 120.400 1534.950 120.460 ;
        RECT 1429.750 16.900 1430.070 16.960 ;
        RECT 1534.630 16.900 1534.950 16.960 ;
        RECT 1429.750 16.760 1534.950 16.900 ;
        RECT 1429.750 16.700 1430.070 16.760 ;
        RECT 1534.630 16.700 1534.950 16.760 ;
      LAYER via ;
        RECT 1534.660 1662.980 1534.920 1663.240 ;
        RECT 1536.960 1662.980 1537.220 1663.240 ;
        RECT 1534.200 1593.960 1534.460 1594.220 ;
        RECT 1534.660 1593.960 1534.920 1594.220 ;
        RECT 1535.120 1545.340 1535.380 1545.600 ;
        RECT 1535.580 1497.400 1535.840 1497.660 ;
        RECT 1535.580 1466.120 1535.840 1466.380 ;
        RECT 1534.200 1400.840 1534.460 1401.100 ;
        RECT 1533.740 1365.820 1534.000 1366.080 ;
        RECT 1534.660 1365.820 1534.920 1366.080 ;
        RECT 1534.660 1352.220 1534.920 1352.480 ;
        RECT 1534.200 1304.280 1534.460 1304.540 ;
        RECT 1533.740 1269.260 1534.000 1269.520 ;
        RECT 1534.660 1269.260 1534.920 1269.520 ;
        RECT 1534.660 1255.660 1534.920 1255.920 ;
        RECT 1534.200 1207.380 1534.460 1207.640 ;
        RECT 1533.740 1076.140 1534.000 1076.400 ;
        RECT 1534.660 1076.140 1534.920 1076.400 ;
        RECT 1533.740 1014.260 1534.000 1014.520 ;
        RECT 1534.200 1014.260 1534.460 1014.520 ;
        RECT 1534.200 820.800 1534.460 821.060 ;
        RECT 1534.660 820.800 1534.920 821.060 ;
        RECT 1533.740 434.560 1534.000 434.820 ;
        RECT 1533.280 386.280 1533.540 386.540 ;
        RECT 1533.280 372.340 1533.540 372.600 ;
        RECT 1533.740 351.260 1534.000 351.520 ;
        RECT 1533.740 303.320 1534.000 303.580 ;
        RECT 1534.660 303.320 1534.920 303.580 ;
        RECT 1534.660 289.380 1534.920 289.640 ;
        RECT 1534.200 241.440 1534.460 241.700 ;
        RECT 1534.200 234.300 1534.460 234.560 ;
        RECT 1535.120 234.300 1535.380 234.560 ;
        RECT 1535.120 186.020 1535.380 186.280 ;
        RECT 1534.660 120.400 1534.920 120.660 ;
        RECT 1429.780 16.700 1430.040 16.960 ;
        RECT 1534.660 16.700 1534.920 16.960 ;
      LAYER met2 ;
        RECT 1537.410 1700.410 1537.690 1704.000 ;
        RECT 1537.020 1700.270 1537.690 1700.410 ;
        RECT 1537.020 1663.270 1537.160 1700.270 ;
        RECT 1537.410 1700.000 1537.690 1700.270 ;
        RECT 1534.660 1662.950 1534.920 1663.270 ;
        RECT 1536.960 1662.950 1537.220 1663.270 ;
        RECT 1534.720 1594.250 1534.860 1662.950 ;
        RECT 1534.200 1593.930 1534.460 1594.250 ;
        RECT 1534.660 1593.930 1534.920 1594.250 ;
        RECT 1534.260 1593.765 1534.400 1593.930 ;
        RECT 1534.190 1593.395 1534.470 1593.765 ;
        RECT 1535.570 1593.395 1535.850 1593.765 ;
        RECT 1535.640 1546.050 1535.780 1593.395 ;
        RECT 1535.180 1545.910 1535.780 1546.050 ;
        RECT 1535.180 1545.630 1535.320 1545.910 ;
        RECT 1535.120 1545.310 1535.380 1545.630 ;
        RECT 1535.580 1497.370 1535.840 1497.690 ;
        RECT 1535.640 1466.410 1535.780 1497.370 ;
        RECT 1535.580 1466.090 1535.840 1466.410 ;
        RECT 1534.200 1400.810 1534.460 1401.130 ;
        RECT 1534.260 1366.530 1534.400 1400.810 ;
        RECT 1533.800 1366.390 1534.400 1366.530 ;
        RECT 1533.800 1366.110 1533.940 1366.390 ;
        RECT 1533.740 1365.790 1534.000 1366.110 ;
        RECT 1534.660 1365.790 1534.920 1366.110 ;
        RECT 1534.720 1352.510 1534.860 1365.790 ;
        RECT 1534.660 1352.190 1534.920 1352.510 ;
        RECT 1534.200 1304.250 1534.460 1304.570 ;
        RECT 1534.260 1269.970 1534.400 1304.250 ;
        RECT 1533.800 1269.830 1534.400 1269.970 ;
        RECT 1533.800 1269.550 1533.940 1269.830 ;
        RECT 1533.740 1269.230 1534.000 1269.550 ;
        RECT 1534.660 1269.230 1534.920 1269.550 ;
        RECT 1534.720 1255.950 1534.860 1269.230 ;
        RECT 1534.660 1255.630 1534.920 1255.950 ;
        RECT 1534.260 1207.670 1534.400 1207.825 ;
        RECT 1534.200 1207.410 1534.460 1207.670 ;
        RECT 1534.200 1207.350 1534.860 1207.410 ;
        RECT 1534.260 1207.270 1534.860 1207.350 ;
        RECT 1534.720 1124.450 1534.860 1207.270 ;
        RECT 1534.260 1124.310 1534.860 1124.450 ;
        RECT 1534.260 1076.850 1534.400 1124.310 ;
        RECT 1533.800 1076.710 1534.400 1076.850 ;
        RECT 1533.800 1076.430 1533.940 1076.710 ;
        RECT 1533.740 1076.110 1534.000 1076.430 ;
        RECT 1534.660 1076.110 1534.920 1076.430 ;
        RECT 1534.720 1062.685 1534.860 1076.110 ;
        RECT 1533.730 1062.315 1534.010 1062.685 ;
        RECT 1534.650 1062.315 1534.930 1062.685 ;
        RECT 1533.800 1014.550 1533.940 1062.315 ;
        RECT 1533.740 1014.230 1534.000 1014.550 ;
        RECT 1534.200 1014.230 1534.460 1014.550 ;
        RECT 1534.260 983.010 1534.400 1014.230 ;
        RECT 1534.260 982.870 1534.860 983.010 ;
        RECT 1534.720 931.330 1534.860 982.870 ;
        RECT 1534.260 931.190 1534.860 931.330 ;
        RECT 1534.260 862.650 1534.400 931.190 ;
        RECT 1534.260 862.510 1534.860 862.650 ;
        RECT 1534.720 834.770 1534.860 862.510 ;
        RECT 1534.260 834.630 1534.860 834.770 ;
        RECT 1534.260 821.090 1534.400 834.630 ;
        RECT 1534.200 820.770 1534.460 821.090 ;
        RECT 1534.660 820.770 1534.920 821.090 ;
        RECT 1534.720 738.210 1534.860 820.770 ;
        RECT 1534.260 738.070 1534.860 738.210 ;
        RECT 1534.260 700.130 1534.400 738.070 ;
        RECT 1533.340 699.990 1534.400 700.130 ;
        RECT 1533.340 676.445 1533.480 699.990 ;
        RECT 1533.270 676.075 1533.550 676.445 ;
        RECT 1534.650 676.075 1534.930 676.445 ;
        RECT 1534.720 641.650 1534.860 676.075 ;
        RECT 1534.260 641.510 1534.860 641.650 ;
        RECT 1534.260 627.880 1534.400 641.510 ;
        RECT 1533.340 627.740 1534.400 627.880 ;
        RECT 1533.340 579.885 1533.480 627.740 ;
        RECT 1533.270 579.515 1533.550 579.885 ;
        RECT 1534.650 579.515 1534.930 579.885 ;
        RECT 1534.720 545.090 1534.860 579.515 ;
        RECT 1534.260 544.950 1534.860 545.090 ;
        RECT 1534.260 507.010 1534.400 544.950 ;
        RECT 1533.340 506.870 1534.400 507.010 ;
        RECT 1533.340 483.325 1533.480 506.870 ;
        RECT 1533.270 482.955 1533.550 483.325 ;
        RECT 1534.650 482.955 1534.930 483.325 ;
        RECT 1534.720 448.530 1534.860 482.955 ;
        RECT 1533.800 448.390 1534.860 448.530 ;
        RECT 1533.800 434.850 1533.940 448.390 ;
        RECT 1533.740 434.530 1534.000 434.850 ;
        RECT 1533.280 386.250 1533.540 386.570 ;
        RECT 1533.340 372.630 1533.480 386.250 ;
        RECT 1533.280 372.310 1533.540 372.630 ;
        RECT 1533.740 351.230 1534.000 351.550 ;
        RECT 1533.800 303.610 1533.940 351.230 ;
        RECT 1533.740 303.290 1534.000 303.610 ;
        RECT 1534.660 303.290 1534.920 303.610 ;
        RECT 1534.720 289.670 1534.860 303.290 ;
        RECT 1534.660 289.350 1534.920 289.670 ;
        RECT 1534.200 241.410 1534.460 241.730 ;
        RECT 1534.260 234.590 1534.400 241.410 ;
        RECT 1534.200 234.270 1534.460 234.590 ;
        RECT 1535.120 234.270 1535.380 234.590 ;
        RECT 1535.180 186.310 1535.320 234.270 ;
        RECT 1535.120 185.990 1535.380 186.310 ;
        RECT 1534.660 120.370 1534.920 120.690 ;
        RECT 1534.720 16.990 1534.860 120.370 ;
        RECT 1429.780 16.670 1430.040 16.990 ;
        RECT 1534.660 16.670 1534.920 16.990 ;
        RECT 1429.840 2.400 1429.980 16.670 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 1534.190 1593.440 1534.470 1593.720 ;
        RECT 1535.570 1593.440 1535.850 1593.720 ;
        RECT 1533.730 1062.360 1534.010 1062.640 ;
        RECT 1534.650 1062.360 1534.930 1062.640 ;
        RECT 1533.270 676.120 1533.550 676.400 ;
        RECT 1534.650 676.120 1534.930 676.400 ;
        RECT 1533.270 579.560 1533.550 579.840 ;
        RECT 1534.650 579.560 1534.930 579.840 ;
        RECT 1533.270 483.000 1533.550 483.280 ;
        RECT 1534.650 483.000 1534.930 483.280 ;
      LAYER met3 ;
        RECT 1534.165 1593.730 1534.495 1593.745 ;
        RECT 1535.545 1593.730 1535.875 1593.745 ;
        RECT 1534.165 1593.430 1535.875 1593.730 ;
        RECT 1534.165 1593.415 1534.495 1593.430 ;
        RECT 1535.545 1593.415 1535.875 1593.430 ;
        RECT 1533.705 1062.650 1534.035 1062.665 ;
        RECT 1534.625 1062.650 1534.955 1062.665 ;
        RECT 1533.705 1062.350 1534.955 1062.650 ;
        RECT 1533.705 1062.335 1534.035 1062.350 ;
        RECT 1534.625 1062.335 1534.955 1062.350 ;
        RECT 1533.245 676.410 1533.575 676.425 ;
        RECT 1534.625 676.410 1534.955 676.425 ;
        RECT 1533.245 676.110 1534.955 676.410 ;
        RECT 1533.245 676.095 1533.575 676.110 ;
        RECT 1534.625 676.095 1534.955 676.110 ;
        RECT 1533.245 579.850 1533.575 579.865 ;
        RECT 1534.625 579.850 1534.955 579.865 ;
        RECT 1533.245 579.550 1534.955 579.850 ;
        RECT 1533.245 579.535 1533.575 579.550 ;
        RECT 1534.625 579.535 1534.955 579.550 ;
        RECT 1533.245 483.290 1533.575 483.305 ;
        RECT 1534.625 483.290 1534.955 483.305 ;
        RECT 1533.245 482.990 1534.955 483.290 ;
        RECT 1533.245 482.975 1533.575 482.990 ;
        RECT 1534.625 482.975 1534.955 482.990 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 0.300 ;
=======
      LAYER met1 ;
        RECT 1447.690 15.200 1448.010 15.260 ;
        RECT 1540.150 15.200 1540.470 15.260 ;
        RECT 1447.690 15.060 1540.470 15.200 ;
        RECT 1447.690 15.000 1448.010 15.060 ;
        RECT 1540.150 15.000 1540.470 15.060 ;
=======
      LAYER li1 ;
        RECT 1486.865 16.575 1487.035 18.275 ;
        RECT 1486.405 16.405 1487.035 16.575 ;
      LAYER mcon ;
        RECT 1486.865 18.105 1487.035 18.275 ;
      LAYER met1 ;
        RECT 1486.805 18.260 1487.095 18.305 ;
        RECT 1540.150 18.260 1540.470 18.320 ;
        RECT 1486.805 18.120 1540.470 18.260 ;
        RECT 1486.805 18.075 1487.095 18.120 ;
        RECT 1540.150 18.060 1540.470 18.120 ;
        RECT 1447.690 16.560 1448.010 16.620 ;
        RECT 1486.345 16.560 1486.635 16.605 ;
        RECT 1447.690 16.420 1486.635 16.560 ;
        RECT 1447.690 16.360 1448.010 16.420 ;
        RECT 1486.345 16.375 1486.635 16.420 ;
>>>>>>> re-updated local openlane
      LAYER via ;
        RECT 1540.180 18.060 1540.440 18.320 ;
        RECT 1447.720 16.360 1447.980 16.620 ;
      LAYER met2 ;
        RECT 1542.010 1700.410 1542.290 1704.000 ;
        RECT 1541.620 1700.270 1542.290 1700.410 ;
        RECT 1541.620 1656.210 1541.760 1700.270 ;
        RECT 1542.010 1700.000 1542.290 1700.270 ;
        RECT 1540.240 1656.070 1541.760 1656.210 ;
        RECT 1540.240 18.350 1540.380 1656.070 ;
        RECT 1540.180 18.030 1540.440 18.350 ;
        RECT 1447.720 16.330 1447.980 16.650 ;
        RECT 1447.780 2.400 1447.920 16.330 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 0.300 ;
=======
      LAYER li1 ;
        RECT 1488.245 16.065 1488.415 17.255 ;
      LAYER mcon ;
        RECT 1488.245 17.085 1488.415 17.255 ;
      LAYER met1 ;
        RECT 1488.185 17.240 1488.475 17.285 ;
        RECT 1546.130 17.240 1546.450 17.300 ;
        RECT 1488.185 17.100 1546.450 17.240 ;
        RECT 1488.185 17.055 1488.475 17.100 ;
        RECT 1546.130 17.040 1546.450 17.100 ;
        RECT 1465.630 16.220 1465.950 16.280 ;
        RECT 1488.185 16.220 1488.475 16.265 ;
        RECT 1465.630 16.080 1488.475 16.220 ;
        RECT 1465.630 16.020 1465.950 16.080 ;
        RECT 1488.185 16.035 1488.475 16.080 ;
      LAYER via ;
        RECT 1546.160 17.040 1546.420 17.300 ;
        RECT 1465.660 16.020 1465.920 16.280 ;
      LAYER met2 ;
        RECT 1545.690 1700.410 1545.970 1704.000 ;
        RECT 1545.690 1700.270 1546.360 1700.410 ;
        RECT 1545.690 1700.000 1545.970 1700.270 ;
        RECT 1546.220 17.330 1546.360 1700.270 ;
        RECT 1546.160 17.010 1546.420 17.330 ;
        RECT 1465.660 15.990 1465.920 16.310 ;
        RECT 1465.720 2.400 1465.860 15.990 ;
=======
      LAYER met1 ;
        RECT 1547.050 15.880 1547.370 15.940 ;
        RECT 1524.140 15.740 1547.370 15.880 ;
        RECT 1465.630 15.540 1465.950 15.600 ;
        RECT 1524.140 15.540 1524.280 15.740 ;
        RECT 1547.050 15.680 1547.370 15.740 ;
        RECT 1465.630 15.400 1524.280 15.540 ;
        RECT 1465.630 15.340 1465.950 15.400 ;
      LAYER via ;
        RECT 1465.660 15.340 1465.920 15.600 ;
        RECT 1547.080 15.680 1547.340 15.940 ;
      LAYER met2 ;
        RECT 1547.070 1700.000 1547.350 1704.000 ;
        RECT 1547.140 15.970 1547.280 1700.000 ;
        RECT 1547.080 15.650 1547.340 15.970 ;
        RECT 1465.660 15.310 1465.920 15.630 ;
        RECT 1465.720 2.400 1465.860 15.310 ;
>>>>>>> re-updated local openlane
        RECT 1465.510 -4.800 1466.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1546.590 1678.480 1546.910 1678.540 ;
        RECT 1550.730 1678.480 1551.050 1678.540 ;
        RECT 1546.590 1678.340 1551.050 1678.480 ;
        RECT 1546.590 1678.280 1546.910 1678.340 ;
        RECT 1550.730 1678.280 1551.050 1678.340 ;
        RECT 1483.570 14.180 1483.890 14.240 ;
        RECT 1546.590 14.180 1546.910 14.240 ;
        RECT 1483.570 14.040 1546.910 14.180 ;
        RECT 1483.570 13.980 1483.890 14.040 ;
        RECT 1546.590 13.980 1546.910 14.040 ;
      LAYER via ;
        RECT 1546.620 1678.280 1546.880 1678.540 ;
        RECT 1550.760 1678.280 1551.020 1678.540 ;
        RECT 1483.600 13.980 1483.860 14.240 ;
        RECT 1546.620 13.980 1546.880 14.240 ;
      LAYER met2 ;
        RECT 1552.130 1700.410 1552.410 1704.000 ;
        RECT 1550.820 1700.270 1552.410 1700.410 ;
        RECT 1550.820 1678.570 1550.960 1700.270 ;
        RECT 1552.130 1700.000 1552.410 1700.270 ;
        RECT 1546.620 1678.250 1546.880 1678.570 ;
        RECT 1550.760 1678.250 1551.020 1678.570 ;
        RECT 1546.680 14.270 1546.820 1678.250 ;
        RECT 1483.600 13.950 1483.860 14.270 ;
        RECT 1546.620 13.950 1546.880 14.270 ;
        RECT 1483.660 2.400 1483.800 13.950 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 0.300 ;
=======
      LAYER met1 ;
        RECT 1501.510 18.260 1501.830 18.320 ;
        RECT 1553.950 18.260 1554.270 18.320 ;
        RECT 1501.510 18.120 1554.270 18.260 ;
        RECT 1501.510 18.060 1501.830 18.120 ;
        RECT 1553.950 18.060 1554.270 18.120 ;
      LAYER via ;
        RECT 1501.540 18.060 1501.800 18.320 ;
        RECT 1553.980 18.060 1554.240 18.320 ;
      LAYER met2 ;
        RECT 1554.890 1700.410 1555.170 1704.000 ;
        RECT 1554.040 1700.270 1555.170 1700.410 ;
        RECT 1554.040 18.350 1554.180 1700.270 ;
        RECT 1554.890 1700.000 1555.170 1700.270 ;
        RECT 1501.540 18.030 1501.800 18.350 ;
        RECT 1553.980 18.030 1554.240 18.350 ;
        RECT 1501.600 2.400 1501.740 18.030 ;
=======
      LAYER li1 ;
        RECT 1511.245 17.085 1511.415 19.635 ;
      LAYER mcon ;
        RECT 1511.245 19.465 1511.415 19.635 ;
      LAYER met1 ;
        RECT 1553.950 20.300 1554.270 20.360 ;
        RECT 1528.740 20.160 1554.270 20.300 ;
        RECT 1511.185 19.620 1511.475 19.665 ;
        RECT 1528.740 19.620 1528.880 20.160 ;
        RECT 1553.950 20.100 1554.270 20.160 ;
        RECT 1511.185 19.480 1528.880 19.620 ;
        RECT 1511.185 19.435 1511.475 19.480 ;
        RECT 1501.510 17.240 1501.830 17.300 ;
        RECT 1511.185 17.240 1511.475 17.285 ;
        RECT 1501.510 17.100 1511.475 17.240 ;
        RECT 1501.510 17.040 1501.830 17.100 ;
        RECT 1511.185 17.055 1511.475 17.100 ;
      LAYER via ;
        RECT 1553.980 20.100 1554.240 20.360 ;
        RECT 1501.540 17.040 1501.800 17.300 ;
      LAYER met2 ;
        RECT 1556.730 1700.410 1557.010 1704.000 ;
        RECT 1555.880 1700.270 1557.010 1700.410 ;
        RECT 1555.880 1688.850 1556.020 1700.270 ;
        RECT 1556.730 1700.000 1557.010 1700.270 ;
        RECT 1554.040 1688.710 1556.020 1688.850 ;
        RECT 1554.040 20.390 1554.180 1688.710 ;
        RECT 1553.980 20.070 1554.240 20.390 ;
        RECT 1501.540 17.010 1501.800 17.330 ;
        RECT 1501.600 2.400 1501.740 17.010 ;
>>>>>>> re-updated local openlane
        RECT 1501.390 -4.800 1501.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 0.300 ;
=======
      LAYER met1 ;
        RECT 1518.990 17.920 1519.310 17.980 ;
        RECT 1561.310 17.920 1561.630 17.980 ;
        RECT 1518.990 17.780 1561.630 17.920 ;
        RECT 1518.990 17.720 1519.310 17.780 ;
        RECT 1561.310 17.720 1561.630 17.780 ;
      LAYER via ;
        RECT 1519.020 17.720 1519.280 17.980 ;
        RECT 1561.340 17.720 1561.600 17.980 ;
      LAYER met2 ;
        RECT 1561.790 1700.410 1562.070 1704.000 ;
        RECT 1561.400 1700.270 1562.070 1700.410 ;
        RECT 1561.400 18.010 1561.540 1700.270 ;
        RECT 1561.790 1700.000 1562.070 1700.270 ;
        RECT 1519.020 17.690 1519.280 18.010 ;
        RECT 1561.340 17.690 1561.600 18.010 ;
        RECT 1519.080 2.400 1519.220 17.690 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1338.670 1674.400 1338.990 1674.460 ;
        RECT 1342.810 1674.400 1343.130 1674.460 ;
        RECT 1338.670 1674.260 1343.130 1674.400 ;
        RECT 1338.670 1674.200 1338.990 1674.260 ;
        RECT 1342.810 1674.200 1343.130 1674.260 ;
        RECT 716.290 48.180 716.610 48.240 ;
        RECT 1338.670 48.180 1338.990 48.240 ;
        RECT 716.290 48.040 1338.990 48.180 ;
        RECT 716.290 47.980 716.610 48.040 ;
        RECT 1338.670 47.980 1338.990 48.040 ;
      LAYER via ;
        RECT 1338.700 1674.200 1338.960 1674.460 ;
        RECT 1342.840 1674.200 1343.100 1674.460 ;
        RECT 716.320 47.980 716.580 48.240 ;
        RECT 1338.700 47.980 1338.960 48.240 ;
      LAYER met2 ;
        RECT 1343.750 1700.410 1344.030 1704.000 ;
        RECT 1342.900 1700.270 1344.030 1700.410 ;
        RECT 1342.900 1674.490 1343.040 1700.270 ;
        RECT 1343.750 1700.000 1344.030 1700.270 ;
        RECT 1338.700 1674.170 1338.960 1674.490 ;
        RECT 1342.840 1674.170 1343.100 1674.490 ;
        RECT 1338.760 48.270 1338.900 1674.170 ;
        RECT 716.320 47.950 716.580 48.270 ;
        RECT 1338.700 47.950 1338.960 48.270 ;
        RECT 716.380 2.400 716.520 47.950 ;
        RECT 716.170 -4.800 716.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 0.300 ;
=======
      LAYER li1 ;
        RECT 1562.305 1490.645 1562.475 1529.915 ;
        RECT 1561.845 1200.625 1562.015 1248.735 ;
        RECT 1561.845 689.605 1562.015 724.455 ;
        RECT 1561.845 593.045 1562.015 627.895 ;
        RECT 1561.845 496.485 1562.015 531.335 ;
        RECT 1562.305 179.605 1562.475 227.715 ;
        RECT 1560.005 65.365 1560.175 110.755 ;
      LAYER mcon ;
        RECT 1562.305 1529.745 1562.475 1529.915 ;
        RECT 1561.845 1248.565 1562.015 1248.735 ;
        RECT 1561.845 724.285 1562.015 724.455 ;
        RECT 1561.845 627.725 1562.015 627.895 ;
        RECT 1561.845 531.165 1562.015 531.335 ;
        RECT 1562.305 227.545 1562.475 227.715 ;
        RECT 1560.005 110.585 1560.175 110.755 ;
      LAYER met1 ;
        RECT 1562.230 1692.080 1562.550 1692.140 ;
        RECT 1564.530 1692.080 1564.850 1692.140 ;
        RECT 1562.230 1691.940 1564.850 1692.080 ;
        RECT 1562.230 1691.880 1562.550 1691.940 ;
        RECT 1564.530 1691.880 1564.850 1691.940 ;
        RECT 1561.770 1594.160 1562.090 1594.220 ;
        RECT 1562.230 1594.160 1562.550 1594.220 ;
        RECT 1561.770 1594.020 1562.550 1594.160 ;
        RECT 1561.770 1593.960 1562.090 1594.020 ;
        RECT 1562.230 1593.960 1562.550 1594.020 ;
        RECT 1562.230 1529.900 1562.550 1529.960 ;
        RECT 1562.035 1529.760 1562.550 1529.900 ;
        RECT 1562.230 1529.700 1562.550 1529.760 ;
        RECT 1562.245 1490.800 1562.535 1490.845 ;
        RECT 1562.690 1490.800 1563.010 1490.860 ;
        RECT 1562.245 1490.660 1563.010 1490.800 ;
        RECT 1562.245 1490.615 1562.535 1490.660 ;
        RECT 1562.690 1490.600 1563.010 1490.660 ;
        RECT 1561.770 1442.180 1562.090 1442.240 ;
        RECT 1562.690 1442.180 1563.010 1442.240 ;
        RECT 1561.770 1442.040 1563.010 1442.180 ;
        RECT 1561.770 1441.980 1562.090 1442.040 ;
        RECT 1562.690 1441.980 1563.010 1442.040 ;
        RECT 1561.770 1414.440 1562.090 1414.700 ;
        RECT 1561.860 1414.300 1562.000 1414.440 ;
        RECT 1562.230 1414.300 1562.550 1414.360 ;
        RECT 1561.860 1414.160 1562.550 1414.300 ;
        RECT 1562.230 1414.100 1562.550 1414.160 ;
        RECT 1561.770 1248.720 1562.090 1248.780 ;
        RECT 1561.575 1248.580 1562.090 1248.720 ;
        RECT 1561.770 1248.520 1562.090 1248.580 ;
        RECT 1561.770 1200.780 1562.090 1200.840 ;
        RECT 1561.575 1200.640 1562.090 1200.780 ;
        RECT 1561.770 1200.580 1562.090 1200.640 ;
        RECT 1561.310 1124.960 1561.630 1125.020 ;
        RECT 1562.230 1124.960 1562.550 1125.020 ;
        RECT 1561.310 1124.820 1562.550 1124.960 ;
        RECT 1561.310 1124.760 1561.630 1124.820 ;
        RECT 1562.230 1124.760 1562.550 1124.820 ;
        RECT 1561.310 1028.400 1561.630 1028.460 ;
        RECT 1562.230 1028.400 1562.550 1028.460 ;
        RECT 1561.310 1028.260 1562.550 1028.400 ;
        RECT 1561.310 1028.200 1561.630 1028.260 ;
        RECT 1562.230 1028.200 1562.550 1028.260 ;
        RECT 1561.310 931.840 1561.630 931.900 ;
        RECT 1562.230 931.840 1562.550 931.900 ;
        RECT 1561.310 931.700 1562.550 931.840 ;
        RECT 1561.310 931.640 1561.630 931.700 ;
        RECT 1562.230 931.640 1562.550 931.700 ;
        RECT 1560.850 869.620 1561.170 869.680 ;
        RECT 1562.230 869.620 1562.550 869.680 ;
        RECT 1560.850 869.480 1562.550 869.620 ;
        RECT 1560.850 869.420 1561.170 869.480 ;
        RECT 1562.230 869.420 1562.550 869.480 ;
        RECT 1561.310 818.280 1561.630 818.340 ;
        RECT 1562.230 818.280 1562.550 818.340 ;
        RECT 1561.310 818.140 1562.550 818.280 ;
        RECT 1561.310 818.080 1561.630 818.140 ;
        RECT 1562.230 818.080 1562.550 818.140 ;
        RECT 1561.770 724.440 1562.090 724.500 ;
        RECT 1561.575 724.300 1562.090 724.440 ;
        RECT 1561.770 724.240 1562.090 724.300 ;
        RECT 1561.770 689.760 1562.090 689.820 ;
        RECT 1561.575 689.620 1562.090 689.760 ;
        RECT 1561.770 689.560 1562.090 689.620 ;
        RECT 1561.310 641.820 1561.630 641.880 ;
        RECT 1562.230 641.820 1562.550 641.880 ;
        RECT 1561.310 641.680 1562.550 641.820 ;
        RECT 1561.310 641.620 1561.630 641.680 ;
        RECT 1562.230 641.620 1562.550 641.680 ;
        RECT 1561.770 627.880 1562.090 627.940 ;
        RECT 1561.575 627.740 1562.090 627.880 ;
        RECT 1561.770 627.680 1562.090 627.740 ;
        RECT 1561.770 593.200 1562.090 593.260 ;
        RECT 1561.575 593.060 1562.090 593.200 ;
        RECT 1561.770 593.000 1562.090 593.060 ;
        RECT 1561.310 545.260 1561.630 545.320 ;
        RECT 1562.230 545.260 1562.550 545.320 ;
        RECT 1561.310 545.120 1562.550 545.260 ;
        RECT 1561.310 545.060 1561.630 545.120 ;
        RECT 1562.230 545.060 1562.550 545.120 ;
        RECT 1561.770 531.320 1562.090 531.380 ;
        RECT 1561.575 531.180 1562.090 531.320 ;
        RECT 1561.770 531.120 1562.090 531.180 ;
        RECT 1561.770 496.640 1562.090 496.700 ;
        RECT 1561.575 496.500 1562.090 496.640 ;
        RECT 1561.770 496.440 1562.090 496.500 ;
        RECT 1561.310 448.360 1561.630 448.420 ;
        RECT 1562.230 448.360 1562.550 448.420 ;
        RECT 1561.310 448.220 1562.550 448.360 ;
        RECT 1561.310 448.160 1561.630 448.220 ;
        RECT 1562.230 448.160 1562.550 448.220 ;
        RECT 1560.850 338.200 1561.170 338.260 ;
        RECT 1561.310 338.200 1561.630 338.260 ;
        RECT 1560.850 338.060 1561.630 338.200 ;
        RECT 1560.850 338.000 1561.170 338.060 ;
        RECT 1561.310 338.000 1561.630 338.060 ;
        RECT 1560.850 302.840 1561.170 302.900 ;
        RECT 1561.770 302.840 1562.090 302.900 ;
        RECT 1560.850 302.700 1562.090 302.840 ;
        RECT 1560.850 302.640 1561.170 302.700 ;
        RECT 1561.770 302.640 1562.090 302.700 ;
        RECT 1561.770 255.380 1562.090 255.640 ;
        RECT 1561.860 254.900 1562.000 255.380 ;
        RECT 1562.690 254.900 1563.010 254.960 ;
        RECT 1561.860 254.760 1563.010 254.900 ;
        RECT 1562.690 254.700 1563.010 254.760 ;
        RECT 1562.245 227.700 1562.535 227.745 ;
        RECT 1562.690 227.700 1563.010 227.760 ;
        RECT 1562.245 227.560 1563.010 227.700 ;
        RECT 1562.245 227.515 1562.535 227.560 ;
        RECT 1562.690 227.500 1563.010 227.560 ;
        RECT 1562.230 179.760 1562.550 179.820 ;
        RECT 1562.035 179.620 1562.550 179.760 ;
        RECT 1562.230 179.560 1562.550 179.620 ;
        RECT 1559.945 110.740 1560.235 110.785 ;
        RECT 1561.310 110.740 1561.630 110.800 ;
        RECT 1559.945 110.600 1561.630 110.740 ;
        RECT 1559.945 110.555 1560.235 110.600 ;
        RECT 1561.310 110.540 1561.630 110.600 ;
        RECT 1559.945 65.520 1560.235 65.565 ;
        RECT 1561.770 65.520 1562.090 65.580 ;
        RECT 1559.945 65.380 1562.090 65.520 ;
        RECT 1559.945 65.335 1560.235 65.380 ;
        RECT 1561.770 65.320 1562.090 65.380 ;
        RECT 1536.930 16.900 1537.250 16.960 ;
        RECT 1561.770 16.900 1562.090 16.960 ;
        RECT 1536.930 16.760 1562.090 16.900 ;
        RECT 1536.930 16.700 1537.250 16.760 ;
        RECT 1561.770 16.700 1562.090 16.760 ;
      LAYER via ;
        RECT 1562.260 1691.880 1562.520 1692.140 ;
        RECT 1564.560 1691.880 1564.820 1692.140 ;
        RECT 1561.800 1593.960 1562.060 1594.220 ;
        RECT 1562.260 1593.960 1562.520 1594.220 ;
        RECT 1562.260 1529.700 1562.520 1529.960 ;
        RECT 1562.720 1490.600 1562.980 1490.860 ;
        RECT 1561.800 1441.980 1562.060 1442.240 ;
        RECT 1562.720 1441.980 1562.980 1442.240 ;
        RECT 1561.800 1414.440 1562.060 1414.700 ;
        RECT 1562.260 1414.100 1562.520 1414.360 ;
        RECT 1561.800 1248.520 1562.060 1248.780 ;
        RECT 1561.800 1200.580 1562.060 1200.840 ;
        RECT 1561.340 1124.760 1561.600 1125.020 ;
        RECT 1562.260 1124.760 1562.520 1125.020 ;
        RECT 1561.340 1028.200 1561.600 1028.460 ;
        RECT 1562.260 1028.200 1562.520 1028.460 ;
        RECT 1561.340 931.640 1561.600 931.900 ;
        RECT 1562.260 931.640 1562.520 931.900 ;
        RECT 1560.880 869.420 1561.140 869.680 ;
        RECT 1562.260 869.420 1562.520 869.680 ;
        RECT 1561.340 818.080 1561.600 818.340 ;
        RECT 1562.260 818.080 1562.520 818.340 ;
        RECT 1561.800 724.240 1562.060 724.500 ;
        RECT 1561.800 689.560 1562.060 689.820 ;
        RECT 1561.340 641.620 1561.600 641.880 ;
        RECT 1562.260 641.620 1562.520 641.880 ;
        RECT 1561.800 627.680 1562.060 627.940 ;
        RECT 1561.800 593.000 1562.060 593.260 ;
        RECT 1561.340 545.060 1561.600 545.320 ;
        RECT 1562.260 545.060 1562.520 545.320 ;
        RECT 1561.800 531.120 1562.060 531.380 ;
        RECT 1561.800 496.440 1562.060 496.700 ;
        RECT 1561.340 448.160 1561.600 448.420 ;
        RECT 1562.260 448.160 1562.520 448.420 ;
        RECT 1560.880 338.000 1561.140 338.260 ;
        RECT 1561.340 338.000 1561.600 338.260 ;
        RECT 1560.880 302.640 1561.140 302.900 ;
        RECT 1561.800 302.640 1562.060 302.900 ;
        RECT 1561.800 255.380 1562.060 255.640 ;
        RECT 1562.720 254.700 1562.980 254.960 ;
        RECT 1562.720 227.500 1562.980 227.760 ;
        RECT 1562.260 179.560 1562.520 179.820 ;
        RECT 1561.340 110.540 1561.600 110.800 ;
        RECT 1561.800 65.320 1562.060 65.580 ;
        RECT 1536.960 16.700 1537.220 16.960 ;
        RECT 1561.800 16.700 1562.060 16.960 ;
      LAYER met2 ;
        RECT 1564.550 1700.000 1564.830 1704.000 ;
        RECT 1564.620 1692.170 1564.760 1700.000 ;
        RECT 1562.260 1691.850 1562.520 1692.170 ;
        RECT 1564.560 1691.850 1564.820 1692.170 ;
        RECT 1562.320 1594.250 1562.460 1691.850 ;
        RECT 1561.800 1593.930 1562.060 1594.250 ;
        RECT 1562.260 1593.930 1562.520 1594.250 ;
        RECT 1561.860 1559.650 1562.000 1593.930 ;
        RECT 1561.860 1559.510 1562.460 1559.650 ;
        RECT 1562.320 1529.990 1562.460 1559.510 ;
        RECT 1562.260 1529.670 1562.520 1529.990 ;
        RECT 1562.720 1490.570 1562.980 1490.890 ;
        RECT 1562.780 1442.270 1562.920 1490.570 ;
        RECT 1561.800 1441.950 1562.060 1442.270 ;
        RECT 1562.720 1441.950 1562.980 1442.270 ;
        RECT 1561.860 1414.730 1562.000 1441.950 ;
        RECT 1561.800 1414.410 1562.060 1414.730 ;
        RECT 1562.260 1414.070 1562.520 1414.390 ;
        RECT 1562.320 1316.890 1562.460 1414.070 ;
        RECT 1561.400 1316.750 1562.460 1316.890 ;
        RECT 1561.400 1248.890 1561.540 1316.750 ;
        RECT 1561.400 1248.810 1562.000 1248.890 ;
        RECT 1561.400 1248.750 1562.060 1248.810 ;
        RECT 1561.800 1248.490 1562.060 1248.750 ;
        RECT 1561.800 1200.550 1562.060 1200.870 ;
        RECT 1561.860 1173.410 1562.000 1200.550 ;
        RECT 1561.860 1173.270 1562.460 1173.410 ;
        RECT 1562.320 1125.050 1562.460 1173.270 ;
        RECT 1561.340 1124.730 1561.600 1125.050 ;
        RECT 1562.260 1124.730 1562.520 1125.050 ;
        RECT 1561.400 1124.450 1561.540 1124.730 ;
        RECT 1561.400 1124.310 1562.000 1124.450 ;
        RECT 1561.860 1076.850 1562.000 1124.310 ;
        RECT 1561.860 1076.710 1562.460 1076.850 ;
        RECT 1562.320 1028.490 1562.460 1076.710 ;
        RECT 1561.340 1028.170 1561.600 1028.490 ;
        RECT 1562.260 1028.170 1562.520 1028.490 ;
        RECT 1561.400 1027.890 1561.540 1028.170 ;
        RECT 1561.400 1027.750 1562.000 1027.890 ;
        RECT 1561.860 980.290 1562.000 1027.750 ;
        RECT 1561.860 980.150 1562.460 980.290 ;
        RECT 1562.320 931.930 1562.460 980.150 ;
        RECT 1561.340 931.610 1561.600 931.930 ;
        RECT 1562.260 931.610 1562.520 931.930 ;
        RECT 1561.400 931.330 1561.540 931.610 ;
        RECT 1561.400 931.190 1562.000 931.330 ;
        RECT 1561.860 917.845 1562.000 931.190 ;
        RECT 1560.870 917.475 1561.150 917.845 ;
        RECT 1561.790 917.475 1562.070 917.845 ;
        RECT 1560.940 869.710 1561.080 917.475 ;
        RECT 1560.880 869.390 1561.140 869.710 ;
        RECT 1562.260 869.390 1562.520 869.710 ;
        RECT 1562.320 818.370 1562.460 869.390 ;
        RECT 1561.340 818.050 1561.600 818.370 ;
        RECT 1562.260 818.050 1562.520 818.370 ;
        RECT 1561.400 787.170 1561.540 818.050 ;
        RECT 1560.940 787.030 1561.540 787.170 ;
        RECT 1560.940 766.090 1561.080 787.030 ;
        RECT 1560.940 765.950 1561.540 766.090 ;
        RECT 1561.400 738.210 1561.540 765.950 ;
        RECT 1561.400 738.070 1562.000 738.210 ;
        RECT 1561.860 724.530 1562.000 738.070 ;
        RECT 1561.800 724.210 1562.060 724.530 ;
        RECT 1561.800 689.530 1562.060 689.850 ;
        RECT 1561.860 676.330 1562.000 689.530 ;
        RECT 1561.860 676.190 1562.460 676.330 ;
        RECT 1562.320 641.910 1562.460 676.190 ;
        RECT 1561.340 641.650 1561.600 641.910 ;
        RECT 1561.340 641.590 1562.000 641.650 ;
        RECT 1562.260 641.590 1562.520 641.910 ;
        RECT 1561.400 641.510 1562.000 641.590 ;
        RECT 1561.860 627.970 1562.000 641.510 ;
        RECT 1561.800 627.650 1562.060 627.970 ;
        RECT 1561.800 592.970 1562.060 593.290 ;
        RECT 1561.860 579.770 1562.000 592.970 ;
        RECT 1561.860 579.630 1562.460 579.770 ;
        RECT 1562.320 545.350 1562.460 579.630 ;
        RECT 1561.340 545.090 1561.600 545.350 ;
        RECT 1561.340 545.030 1562.000 545.090 ;
        RECT 1562.260 545.030 1562.520 545.350 ;
        RECT 1561.400 544.950 1562.000 545.030 ;
        RECT 1561.860 531.410 1562.000 544.950 ;
        RECT 1561.800 531.090 1562.060 531.410 ;
        RECT 1561.800 496.410 1562.060 496.730 ;
        RECT 1561.860 483.210 1562.000 496.410 ;
        RECT 1561.860 483.070 1562.460 483.210 ;
        RECT 1562.320 448.450 1562.460 483.070 ;
        RECT 1561.340 448.130 1561.600 448.450 ;
        RECT 1562.260 448.130 1562.520 448.450 ;
        RECT 1561.400 400.930 1561.540 448.130 ;
        RECT 1560.940 400.790 1561.540 400.930 ;
        RECT 1560.940 400.250 1561.080 400.790 ;
        RECT 1560.940 400.110 1561.540 400.250 ;
        RECT 1561.400 338.290 1561.540 400.110 ;
        RECT 1560.880 337.970 1561.140 338.290 ;
        RECT 1561.340 337.970 1561.600 338.290 ;
        RECT 1560.940 302.930 1561.080 337.970 ;
        RECT 1560.880 302.610 1561.140 302.930 ;
        RECT 1561.800 302.610 1562.060 302.930 ;
        RECT 1561.860 255.670 1562.000 302.610 ;
        RECT 1561.800 255.350 1562.060 255.670 ;
        RECT 1562.720 254.670 1562.980 254.990 ;
        RECT 1562.780 227.790 1562.920 254.670 ;
        RECT 1562.720 227.470 1562.980 227.790 ;
        RECT 1562.260 179.530 1562.520 179.850 ;
        RECT 1562.320 154.770 1562.460 179.530 ;
        RECT 1561.400 154.630 1562.460 154.770 ;
        RECT 1561.400 110.830 1561.540 154.630 ;
        RECT 1561.340 110.510 1561.600 110.830 ;
        RECT 1561.800 65.290 1562.060 65.610 ;
        RECT 1561.860 16.990 1562.000 65.290 ;
        RECT 1536.960 16.670 1537.220 16.990 ;
        RECT 1561.800 16.670 1562.060 16.990 ;
        RECT 1537.020 2.400 1537.160 16.670 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
      LAYER via2 ;
        RECT 1560.870 917.520 1561.150 917.800 ;
        RECT 1561.790 917.520 1562.070 917.800 ;
      LAYER met3 ;
        RECT 1560.845 917.810 1561.175 917.825 ;
        RECT 1561.765 917.810 1562.095 917.825 ;
        RECT 1560.845 917.510 1562.095 917.810 ;
        RECT 1560.845 917.495 1561.175 917.510 ;
        RECT 1561.765 917.495 1562.095 917.510 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1555.790 1688.340 1556.110 1688.400 ;
        RECT 1566.370 1688.340 1566.690 1688.400 ;
        RECT 1555.790 1688.200 1566.690 1688.340 ;
        RECT 1555.790 1688.140 1556.110 1688.200 ;
        RECT 1566.370 1688.140 1566.690 1688.200 ;
        RECT 1536.930 19.960 1537.250 20.020 ;
        RECT 1555.790 19.960 1556.110 20.020 ;
        RECT 1536.930 19.820 1556.110 19.960 ;
        RECT 1536.930 19.760 1537.250 19.820 ;
        RECT 1555.790 19.760 1556.110 19.820 ;
      LAYER via ;
        RECT 1555.820 1688.140 1556.080 1688.400 ;
        RECT 1566.400 1688.140 1566.660 1688.400 ;
        RECT 1536.960 19.760 1537.220 20.020 ;
        RECT 1555.820 19.760 1556.080 20.020 ;
      LAYER met2 ;
        RECT 1566.390 1700.000 1566.670 1704.000 ;
        RECT 1566.460 1688.430 1566.600 1700.000 ;
        RECT 1555.820 1688.110 1556.080 1688.430 ;
        RECT 1566.400 1688.110 1566.660 1688.430 ;
        RECT 1555.880 20.050 1556.020 1688.110 ;
        RECT 1536.960 19.730 1537.220 20.050 ;
        RECT 1555.820 19.730 1556.080 20.050 ;
        RECT 1537.020 2.400 1537.160 19.730 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1568.670 1694.800 1568.990 1694.860 ;
        RECT 1571.430 1694.800 1571.750 1694.860 ;
        RECT 1568.670 1694.660 1571.750 1694.800 ;
        RECT 1568.670 1694.600 1568.990 1694.660 ;
        RECT 1571.430 1694.600 1571.750 1694.660 ;
        RECT 1554.870 20.300 1555.190 20.360 ;
        RECT 1567.750 20.300 1568.070 20.360 ;
        RECT 1554.870 20.160 1568.070 20.300 ;
        RECT 1554.870 20.100 1555.190 20.160 ;
        RECT 1567.750 20.100 1568.070 20.160 ;
      LAYER via ;
        RECT 1568.700 1694.600 1568.960 1694.860 ;
        RECT 1571.460 1694.600 1571.720 1694.860 ;
        RECT 1554.900 20.100 1555.160 20.360 ;
        RECT 1567.780 20.100 1568.040 20.360 ;
      LAYER met2 ;
        RECT 1571.450 1700.000 1571.730 1704.000 ;
        RECT 1571.520 1694.890 1571.660 1700.000 ;
        RECT 1568.700 1694.570 1568.960 1694.890 ;
        RECT 1571.460 1694.570 1571.720 1694.890 ;
        RECT 1568.760 1656.210 1568.900 1694.570 ;
        RECT 1567.840 1656.070 1568.900 1656.210 ;
        RECT 1567.840 20.390 1567.980 1656.070 ;
        RECT 1554.900 20.070 1555.160 20.390 ;
        RECT 1567.780 20.070 1568.040 20.390 ;
        RECT 1554.960 2.400 1555.100 20.070 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 0.300 ;
=======
      LAYER li1 ;
        RECT 1574.265 1442.025 1574.435 1490.475 ;
        RECT 1574.265 572.645 1574.435 620.755 ;
        RECT 1574.265 476.085 1574.435 524.195 ;
        RECT 1574.265 379.525 1574.435 427.635 ;
        RECT 1574.265 282.965 1574.435 331.075 ;
        RECT 1574.265 186.405 1574.435 234.515 ;
        RECT 1574.265 48.365 1574.435 137.955 ;
      LAYER mcon ;
        RECT 1574.265 1490.305 1574.435 1490.475 ;
        RECT 1574.265 620.585 1574.435 620.755 ;
        RECT 1574.265 524.025 1574.435 524.195 ;
        RECT 1574.265 427.465 1574.435 427.635 ;
        RECT 1574.265 330.905 1574.435 331.075 ;
        RECT 1574.265 234.345 1574.435 234.515 ;
        RECT 1574.265 137.785 1574.435 137.955 ;
      LAYER met1 ;
        RECT 1574.190 1498.080 1574.510 1498.340 ;
        RECT 1574.280 1497.660 1574.420 1498.080 ;
        RECT 1574.190 1497.400 1574.510 1497.660 ;
        RECT 1574.190 1490.460 1574.510 1490.520 ;
        RECT 1573.995 1490.320 1574.510 1490.460 ;
        RECT 1574.190 1490.260 1574.510 1490.320 ;
        RECT 1574.190 1442.180 1574.510 1442.240 ;
        RECT 1573.995 1442.040 1574.510 1442.180 ;
        RECT 1574.190 1441.980 1574.510 1442.040 ;
        RECT 1574.190 1401.520 1574.510 1401.780 ;
        RECT 1574.280 1401.100 1574.420 1401.520 ;
        RECT 1574.190 1400.840 1574.510 1401.100 ;
        RECT 1574.190 1345.620 1574.510 1345.680 ;
        RECT 1575.110 1345.620 1575.430 1345.680 ;
        RECT 1574.190 1345.480 1575.430 1345.620 ;
        RECT 1574.190 1345.420 1574.510 1345.480 ;
        RECT 1575.110 1345.420 1575.430 1345.480 ;
        RECT 1574.190 1304.960 1574.510 1305.220 ;
        RECT 1574.280 1304.540 1574.420 1304.960 ;
        RECT 1574.190 1304.280 1574.510 1304.540 ;
        RECT 1574.190 1249.060 1574.510 1249.120 ;
        RECT 1575.110 1249.060 1575.430 1249.120 ;
        RECT 1574.190 1248.920 1575.430 1249.060 ;
        RECT 1574.190 1248.860 1574.510 1248.920 ;
        RECT 1575.110 1248.860 1575.430 1248.920 ;
        RECT 1574.190 1207.580 1574.510 1207.640 ;
        RECT 1574.650 1207.580 1574.970 1207.640 ;
        RECT 1574.190 1207.440 1574.970 1207.580 ;
        RECT 1574.190 1207.380 1574.510 1207.440 ;
        RECT 1574.650 1207.380 1574.970 1207.440 ;
        RECT 1574.190 1152.500 1574.510 1152.560 ;
        RECT 1575.110 1152.500 1575.430 1152.560 ;
        RECT 1574.190 1152.360 1575.430 1152.500 ;
        RECT 1574.190 1152.300 1574.510 1152.360 ;
        RECT 1575.110 1152.300 1575.430 1152.360 ;
        RECT 1574.190 1007.320 1574.510 1007.380 ;
        RECT 1575.110 1007.320 1575.430 1007.380 ;
        RECT 1574.190 1007.180 1575.430 1007.320 ;
        RECT 1574.190 1007.120 1574.510 1007.180 ;
        RECT 1575.110 1007.120 1575.430 1007.180 ;
        RECT 1574.190 910.760 1574.510 910.820 ;
        RECT 1575.110 910.760 1575.430 910.820 ;
        RECT 1574.190 910.620 1575.430 910.760 ;
        RECT 1574.190 910.560 1574.510 910.620 ;
        RECT 1575.110 910.560 1575.430 910.620 ;
        RECT 1574.190 814.200 1574.510 814.260 ;
        RECT 1575.110 814.200 1575.430 814.260 ;
        RECT 1574.190 814.060 1575.430 814.200 ;
        RECT 1574.190 814.000 1574.510 814.060 ;
        RECT 1575.110 814.000 1575.430 814.060 ;
        RECT 1574.190 717.640 1574.510 717.700 ;
        RECT 1575.110 717.640 1575.430 717.700 ;
        RECT 1574.190 717.500 1575.430 717.640 ;
        RECT 1574.190 717.440 1574.510 717.500 ;
        RECT 1575.110 717.440 1575.430 717.500 ;
        RECT 1574.190 620.740 1574.510 620.800 ;
        RECT 1573.995 620.600 1574.510 620.740 ;
        RECT 1574.190 620.540 1574.510 620.600 ;
        RECT 1574.190 572.800 1574.510 572.860 ;
        RECT 1573.995 572.660 1574.510 572.800 ;
        RECT 1574.190 572.600 1574.510 572.660 ;
        RECT 1574.190 524.180 1574.510 524.240 ;
        RECT 1573.995 524.040 1574.510 524.180 ;
        RECT 1574.190 523.980 1574.510 524.040 ;
        RECT 1574.190 476.240 1574.510 476.300 ;
        RECT 1573.995 476.100 1574.510 476.240 ;
        RECT 1574.190 476.040 1574.510 476.100 ;
        RECT 1574.190 427.620 1574.510 427.680 ;
        RECT 1573.995 427.480 1574.510 427.620 ;
        RECT 1574.190 427.420 1574.510 427.480 ;
        RECT 1574.190 379.680 1574.510 379.740 ;
        RECT 1573.995 379.540 1574.510 379.680 ;
        RECT 1574.190 379.480 1574.510 379.540 ;
        RECT 1574.190 331.060 1574.510 331.120 ;
        RECT 1573.995 330.920 1574.510 331.060 ;
        RECT 1574.190 330.860 1574.510 330.920 ;
        RECT 1574.205 283.120 1574.495 283.165 ;
        RECT 1574.650 283.120 1574.970 283.180 ;
        RECT 1574.205 282.980 1574.970 283.120 ;
        RECT 1574.205 282.935 1574.495 282.980 ;
        RECT 1574.650 282.920 1574.970 282.980 ;
        RECT 1574.190 234.500 1574.510 234.560 ;
        RECT 1573.995 234.360 1574.510 234.500 ;
        RECT 1574.190 234.300 1574.510 234.360 ;
        RECT 1574.205 186.560 1574.495 186.605 ;
        RECT 1574.650 186.560 1574.970 186.620 ;
        RECT 1574.205 186.420 1574.970 186.560 ;
        RECT 1574.205 186.375 1574.495 186.420 ;
        RECT 1574.650 186.360 1574.970 186.420 ;
        RECT 1574.190 137.940 1574.510 138.000 ;
        RECT 1573.995 137.800 1574.510 137.940 ;
        RECT 1574.190 137.740 1574.510 137.800 ;
        RECT 1574.205 48.520 1574.495 48.565 ;
        RECT 1574.650 48.520 1574.970 48.580 ;
        RECT 1574.205 48.380 1574.970 48.520 ;
        RECT 1574.205 48.335 1574.495 48.380 ;
        RECT 1574.650 48.320 1574.970 48.380 ;
        RECT 1572.810 20.300 1573.130 20.360 ;
        RECT 1574.650 20.300 1574.970 20.360 ;
        RECT 1572.810 20.160 1574.970 20.300 ;
        RECT 1572.810 20.100 1573.130 20.160 ;
        RECT 1574.650 20.100 1574.970 20.160 ;
      LAYER via ;
        RECT 1574.220 1498.080 1574.480 1498.340 ;
        RECT 1574.220 1497.400 1574.480 1497.660 ;
        RECT 1574.220 1490.260 1574.480 1490.520 ;
        RECT 1574.220 1441.980 1574.480 1442.240 ;
        RECT 1574.220 1401.520 1574.480 1401.780 ;
        RECT 1574.220 1400.840 1574.480 1401.100 ;
        RECT 1574.220 1345.420 1574.480 1345.680 ;
        RECT 1575.140 1345.420 1575.400 1345.680 ;
        RECT 1574.220 1304.960 1574.480 1305.220 ;
        RECT 1574.220 1304.280 1574.480 1304.540 ;
        RECT 1574.220 1248.860 1574.480 1249.120 ;
        RECT 1575.140 1248.860 1575.400 1249.120 ;
        RECT 1574.220 1207.380 1574.480 1207.640 ;
        RECT 1574.680 1207.380 1574.940 1207.640 ;
        RECT 1574.220 1152.300 1574.480 1152.560 ;
        RECT 1575.140 1152.300 1575.400 1152.560 ;
        RECT 1574.220 1007.120 1574.480 1007.380 ;
        RECT 1575.140 1007.120 1575.400 1007.380 ;
        RECT 1574.220 910.560 1574.480 910.820 ;
        RECT 1575.140 910.560 1575.400 910.820 ;
        RECT 1574.220 814.000 1574.480 814.260 ;
        RECT 1575.140 814.000 1575.400 814.260 ;
        RECT 1574.220 717.440 1574.480 717.700 ;
        RECT 1575.140 717.440 1575.400 717.700 ;
        RECT 1574.220 620.540 1574.480 620.800 ;
        RECT 1574.220 572.600 1574.480 572.860 ;
        RECT 1574.220 523.980 1574.480 524.240 ;
        RECT 1574.220 476.040 1574.480 476.300 ;
        RECT 1574.220 427.420 1574.480 427.680 ;
        RECT 1574.220 379.480 1574.480 379.740 ;
        RECT 1574.220 330.860 1574.480 331.120 ;
        RECT 1574.680 282.920 1574.940 283.180 ;
        RECT 1574.220 234.300 1574.480 234.560 ;
        RECT 1574.680 186.360 1574.940 186.620 ;
        RECT 1574.220 137.740 1574.480 138.000 ;
        RECT 1574.680 48.320 1574.940 48.580 ;
        RECT 1572.840 20.100 1573.100 20.360 ;
        RECT 1574.680 20.100 1574.940 20.360 ;
      LAYER met2 ;
        RECT 1576.050 1700.410 1576.330 1704.000 ;
        RECT 1575.660 1700.270 1576.330 1700.410 ;
        RECT 1575.660 1677.970 1575.800 1700.270 ;
        RECT 1576.050 1700.000 1576.330 1700.270 ;
        RECT 1574.280 1677.830 1575.800 1677.970 ;
        RECT 1574.280 1498.370 1574.420 1677.830 ;
        RECT 1574.220 1498.050 1574.480 1498.370 ;
        RECT 1574.220 1497.370 1574.480 1497.690 ;
        RECT 1574.280 1490.550 1574.420 1497.370 ;
        RECT 1574.220 1490.230 1574.480 1490.550 ;
        RECT 1574.220 1441.950 1574.480 1442.270 ;
        RECT 1574.280 1401.810 1574.420 1441.950 ;
        RECT 1574.220 1401.490 1574.480 1401.810 ;
        RECT 1574.220 1400.810 1574.480 1401.130 ;
        RECT 1574.280 1393.845 1574.420 1400.810 ;
        RECT 1574.210 1393.475 1574.490 1393.845 ;
        RECT 1575.130 1393.475 1575.410 1393.845 ;
        RECT 1575.200 1345.710 1575.340 1393.475 ;
        RECT 1574.220 1345.390 1574.480 1345.710 ;
        RECT 1575.140 1345.390 1575.400 1345.710 ;
        RECT 1574.280 1305.250 1574.420 1345.390 ;
        RECT 1574.220 1304.930 1574.480 1305.250 ;
        RECT 1574.220 1304.250 1574.480 1304.570 ;
        RECT 1574.280 1297.285 1574.420 1304.250 ;
        RECT 1574.210 1296.915 1574.490 1297.285 ;
        RECT 1575.130 1296.915 1575.410 1297.285 ;
        RECT 1575.200 1249.150 1575.340 1296.915 ;
        RECT 1574.220 1248.830 1574.480 1249.150 ;
        RECT 1575.140 1248.830 1575.400 1249.150 ;
        RECT 1574.280 1208.770 1574.420 1248.830 ;
        RECT 1574.280 1208.630 1574.880 1208.770 ;
        RECT 1574.740 1207.670 1574.880 1208.630 ;
        RECT 1574.220 1207.350 1574.480 1207.670 ;
        RECT 1574.680 1207.350 1574.940 1207.670 ;
        RECT 1574.280 1200.725 1574.420 1207.350 ;
        RECT 1574.210 1200.355 1574.490 1200.725 ;
        RECT 1575.130 1200.355 1575.410 1200.725 ;
        RECT 1575.200 1152.590 1575.340 1200.355 ;
        RECT 1574.220 1152.270 1574.480 1152.590 ;
        RECT 1575.140 1152.270 1575.400 1152.590 ;
        RECT 1574.280 1104.165 1574.420 1152.270 ;
        RECT 1574.210 1103.795 1574.490 1104.165 ;
        RECT 1575.130 1103.795 1575.410 1104.165 ;
        RECT 1575.200 1055.885 1575.340 1103.795 ;
        RECT 1574.210 1055.515 1574.490 1055.885 ;
        RECT 1575.130 1055.515 1575.410 1055.885 ;
        RECT 1574.280 1007.410 1574.420 1055.515 ;
        RECT 1574.220 1007.090 1574.480 1007.410 ;
        RECT 1575.140 1007.090 1575.400 1007.410 ;
        RECT 1575.200 959.325 1575.340 1007.090 ;
        RECT 1574.210 958.955 1574.490 959.325 ;
        RECT 1575.130 958.955 1575.410 959.325 ;
        RECT 1574.280 910.850 1574.420 958.955 ;
        RECT 1574.220 910.530 1574.480 910.850 ;
        RECT 1575.140 910.530 1575.400 910.850 ;
        RECT 1575.200 862.765 1575.340 910.530 ;
        RECT 1574.210 862.395 1574.490 862.765 ;
        RECT 1575.130 862.395 1575.410 862.765 ;
        RECT 1574.280 814.290 1574.420 862.395 ;
        RECT 1574.220 813.970 1574.480 814.290 ;
        RECT 1575.140 813.970 1575.400 814.290 ;
        RECT 1575.200 766.205 1575.340 813.970 ;
        RECT 1574.210 765.835 1574.490 766.205 ;
        RECT 1575.130 765.835 1575.410 766.205 ;
        RECT 1574.280 717.730 1574.420 765.835 ;
        RECT 1574.220 717.410 1574.480 717.730 ;
        RECT 1575.140 717.410 1575.400 717.730 ;
        RECT 1575.200 669.645 1575.340 717.410 ;
        RECT 1574.210 669.275 1574.490 669.645 ;
        RECT 1575.130 669.275 1575.410 669.645 ;
        RECT 1574.280 620.830 1574.420 669.275 ;
        RECT 1574.220 620.510 1574.480 620.830 ;
        RECT 1574.220 572.570 1574.480 572.890 ;
        RECT 1574.280 532.285 1574.420 572.570 ;
        RECT 1574.210 531.915 1574.490 532.285 ;
        RECT 1574.210 531.235 1574.490 531.605 ;
        RECT 1574.280 524.270 1574.420 531.235 ;
        RECT 1574.220 523.950 1574.480 524.270 ;
        RECT 1574.220 476.010 1574.480 476.330 ;
        RECT 1574.280 435.725 1574.420 476.010 ;
        RECT 1574.210 435.355 1574.490 435.725 ;
        RECT 1574.210 434.675 1574.490 435.045 ;
        RECT 1574.280 427.710 1574.420 434.675 ;
        RECT 1574.220 427.390 1574.480 427.710 ;
        RECT 1574.220 379.450 1574.480 379.770 ;
        RECT 1574.280 331.150 1574.420 379.450 ;
        RECT 1574.220 330.830 1574.480 331.150 ;
        RECT 1574.680 282.890 1574.940 283.210 ;
        RECT 1574.740 241.810 1574.880 282.890 ;
        RECT 1574.280 241.670 1574.880 241.810 ;
        RECT 1574.280 234.590 1574.420 241.670 ;
        RECT 1574.220 234.270 1574.480 234.590 ;
        RECT 1574.680 186.330 1574.940 186.650 ;
        RECT 1574.740 145.250 1574.880 186.330 ;
        RECT 1574.280 145.110 1574.880 145.250 ;
        RECT 1574.280 138.030 1574.420 145.110 ;
        RECT 1574.220 137.710 1574.480 138.030 ;
        RECT 1574.680 48.290 1574.940 48.610 ;
        RECT 1574.740 20.390 1574.880 48.290 ;
        RECT 1572.840 20.070 1573.100 20.390 ;
        RECT 1574.680 20.070 1574.940 20.390 ;
        RECT 1572.900 2.400 1573.040 20.070 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
      LAYER via2 ;
        RECT 1574.210 1393.520 1574.490 1393.800 ;
        RECT 1575.130 1393.520 1575.410 1393.800 ;
        RECT 1574.210 1296.960 1574.490 1297.240 ;
        RECT 1575.130 1296.960 1575.410 1297.240 ;
        RECT 1574.210 1200.400 1574.490 1200.680 ;
        RECT 1575.130 1200.400 1575.410 1200.680 ;
        RECT 1574.210 1103.840 1574.490 1104.120 ;
        RECT 1575.130 1103.840 1575.410 1104.120 ;
        RECT 1574.210 1055.560 1574.490 1055.840 ;
        RECT 1575.130 1055.560 1575.410 1055.840 ;
        RECT 1574.210 959.000 1574.490 959.280 ;
        RECT 1575.130 959.000 1575.410 959.280 ;
        RECT 1574.210 862.440 1574.490 862.720 ;
        RECT 1575.130 862.440 1575.410 862.720 ;
        RECT 1574.210 765.880 1574.490 766.160 ;
        RECT 1575.130 765.880 1575.410 766.160 ;
        RECT 1574.210 669.320 1574.490 669.600 ;
        RECT 1575.130 669.320 1575.410 669.600 ;
        RECT 1574.210 531.960 1574.490 532.240 ;
        RECT 1574.210 531.280 1574.490 531.560 ;
        RECT 1574.210 435.400 1574.490 435.680 ;
        RECT 1574.210 434.720 1574.490 435.000 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1572.805 1200.690 1573.135 1200.705 ;
        RECT 1573.725 1200.690 1574.055 1200.705 ;
        RECT 1572.805 1200.390 1574.055 1200.690 ;
        RECT 1572.805 1200.375 1573.135 1200.390 ;
        RECT 1573.725 1200.375 1574.055 1200.390 ;
        RECT 1572.805 1104.130 1573.135 1104.145 ;
        RECT 1573.725 1104.130 1574.055 1104.145 ;
        RECT 1572.805 1103.830 1574.055 1104.130 ;
        RECT 1572.805 1103.815 1573.135 1103.830 ;
        RECT 1573.725 1103.815 1574.055 1103.830 ;
        RECT 1572.805 1055.850 1573.135 1055.865 ;
        RECT 1573.725 1055.850 1574.055 1055.865 ;
        RECT 1572.805 1055.550 1574.055 1055.850 ;
        RECT 1572.805 1055.535 1573.135 1055.550 ;
        RECT 1573.725 1055.535 1574.055 1055.550 ;
        RECT 1572.805 959.290 1573.135 959.305 ;
        RECT 1573.725 959.290 1574.055 959.305 ;
        RECT 1572.805 958.990 1574.055 959.290 ;
        RECT 1572.805 958.975 1573.135 958.990 ;
        RECT 1573.725 958.975 1574.055 958.990 ;
        RECT 1572.805 862.730 1573.135 862.745 ;
        RECT 1573.725 862.730 1574.055 862.745 ;
        RECT 1572.805 862.430 1574.055 862.730 ;
        RECT 1572.805 862.415 1573.135 862.430 ;
        RECT 1573.725 862.415 1574.055 862.430 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1574.185 1393.810 1574.515 1393.825 ;
        RECT 1575.105 1393.810 1575.435 1393.825 ;
        RECT 1574.185 1393.510 1575.435 1393.810 ;
        RECT 1574.185 1393.495 1574.515 1393.510 ;
        RECT 1575.105 1393.495 1575.435 1393.510 ;
        RECT 1574.185 1297.250 1574.515 1297.265 ;
        RECT 1575.105 1297.250 1575.435 1297.265 ;
        RECT 1574.185 1296.950 1575.435 1297.250 ;
        RECT 1574.185 1296.935 1574.515 1296.950 ;
        RECT 1575.105 1296.935 1575.435 1296.950 ;
        RECT 1574.185 1200.690 1574.515 1200.705 ;
        RECT 1575.105 1200.690 1575.435 1200.705 ;
        RECT 1574.185 1200.390 1575.435 1200.690 ;
        RECT 1574.185 1200.375 1574.515 1200.390 ;
        RECT 1575.105 1200.375 1575.435 1200.390 ;
        RECT 1574.185 1104.130 1574.515 1104.145 ;
        RECT 1575.105 1104.130 1575.435 1104.145 ;
        RECT 1574.185 1103.830 1575.435 1104.130 ;
        RECT 1574.185 1103.815 1574.515 1103.830 ;
        RECT 1575.105 1103.815 1575.435 1103.830 ;
        RECT 1574.185 1055.850 1574.515 1055.865 ;
        RECT 1575.105 1055.850 1575.435 1055.865 ;
        RECT 1574.185 1055.550 1575.435 1055.850 ;
        RECT 1574.185 1055.535 1574.515 1055.550 ;
        RECT 1575.105 1055.535 1575.435 1055.550 ;
        RECT 1574.185 959.290 1574.515 959.305 ;
        RECT 1575.105 959.290 1575.435 959.305 ;
        RECT 1574.185 958.990 1575.435 959.290 ;
        RECT 1574.185 958.975 1574.515 958.990 ;
        RECT 1575.105 958.975 1575.435 958.990 ;
        RECT 1574.185 862.730 1574.515 862.745 ;
        RECT 1575.105 862.730 1575.435 862.745 ;
        RECT 1574.185 862.430 1575.435 862.730 ;
        RECT 1574.185 862.415 1574.515 862.430 ;
        RECT 1575.105 862.415 1575.435 862.430 ;
        RECT 1574.185 766.170 1574.515 766.185 ;
        RECT 1575.105 766.170 1575.435 766.185 ;
        RECT 1574.185 765.870 1575.435 766.170 ;
        RECT 1574.185 765.855 1574.515 765.870 ;
        RECT 1575.105 765.855 1575.435 765.870 ;
        RECT 1574.185 669.610 1574.515 669.625 ;
        RECT 1575.105 669.610 1575.435 669.625 ;
        RECT 1574.185 669.310 1575.435 669.610 ;
        RECT 1574.185 669.295 1574.515 669.310 ;
        RECT 1575.105 669.295 1575.435 669.310 ;
        RECT 1574.185 532.250 1574.515 532.265 ;
        RECT 1573.510 531.950 1574.515 532.250 ;
        RECT 1573.510 531.570 1573.810 531.950 ;
        RECT 1574.185 531.935 1574.515 531.950 ;
        RECT 1574.185 531.570 1574.515 531.585 ;
        RECT 1573.510 531.270 1574.515 531.570 ;
        RECT 1574.185 531.255 1574.515 531.270 ;
        RECT 1574.185 435.690 1574.515 435.705 ;
        RECT 1573.510 435.390 1574.515 435.690 ;
        RECT 1573.510 435.010 1573.810 435.390 ;
        RECT 1574.185 435.375 1574.515 435.390 ;
        RECT 1574.185 435.010 1574.515 435.025 ;
        RECT 1573.510 434.710 1574.515 435.010 ;
        RECT 1574.185 434.695 1574.515 434.710 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1581.090 1684.260 1581.410 1684.320 ;
        RECT 1585.690 1684.260 1586.010 1684.320 ;
        RECT 1581.090 1684.120 1586.010 1684.260 ;
        RECT 1581.090 1684.060 1581.410 1684.120 ;
        RECT 1585.690 1684.060 1586.010 1684.120 ;
        RECT 1585.690 20.640 1586.010 20.700 ;
        RECT 1590.290 20.640 1590.610 20.700 ;
        RECT 1585.690 20.500 1590.610 20.640 ;
        RECT 1585.690 20.440 1586.010 20.500 ;
        RECT 1590.290 20.440 1590.610 20.500 ;
      LAYER via ;
        RECT 1581.120 1684.060 1581.380 1684.320 ;
        RECT 1585.720 1684.060 1585.980 1684.320 ;
        RECT 1585.720 20.440 1585.980 20.700 ;
        RECT 1590.320 20.440 1590.580 20.700 ;
      LAYER met2 ;
        RECT 1581.110 1700.000 1581.390 1704.000 ;
        RECT 1581.180 1684.350 1581.320 1700.000 ;
        RECT 1581.120 1684.030 1581.380 1684.350 ;
        RECT 1585.720 1684.030 1585.980 1684.350 ;
        RECT 1585.780 20.730 1585.920 1684.030 ;
        RECT 1585.720 20.410 1585.980 20.730 ;
        RECT 1590.320 20.410 1590.580 20.730 ;
        RECT 1590.380 2.400 1590.520 20.410 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 0.300 ;
=======
      LAYER met1 ;
        RECT 1586.150 15.880 1586.470 15.940 ;
        RECT 1608.230 15.880 1608.550 15.940 ;
        RECT 1586.150 15.740 1608.550 15.880 ;
        RECT 1586.150 15.680 1586.470 15.740 ;
        RECT 1608.230 15.680 1608.550 15.740 ;
      LAYER via ;
        RECT 1586.180 15.680 1586.440 15.940 ;
        RECT 1608.260 15.680 1608.520 15.940 ;
      LAYER met2 ;
        RECT 1585.710 1700.410 1585.990 1704.000 ;
        RECT 1585.710 1700.270 1586.380 1700.410 ;
        RECT 1585.710 1700.000 1585.990 1700.270 ;
        RECT 1586.240 15.970 1586.380 1700.270 ;
        RECT 1586.180 15.650 1586.440 15.970 ;
        RECT 1608.260 15.650 1608.520 15.970 ;
        RECT 1608.320 2.400 1608.460 15.650 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1590.750 1684.600 1591.070 1684.660 ;
        RECT 1593.510 1684.600 1593.830 1684.660 ;
        RECT 1590.750 1684.460 1593.830 1684.600 ;
        RECT 1590.750 1684.400 1591.070 1684.460 ;
        RECT 1593.510 1684.400 1593.830 1684.460 ;
        RECT 1593.510 14.520 1593.830 14.580 ;
        RECT 1626.170 14.520 1626.490 14.580 ;
        RECT 1593.510 14.380 1626.490 14.520 ;
        RECT 1593.510 14.320 1593.830 14.380 ;
        RECT 1626.170 14.320 1626.490 14.380 ;
      LAYER via ;
        RECT 1590.780 1684.400 1591.040 1684.660 ;
        RECT 1593.540 1684.400 1593.800 1684.660 ;
        RECT 1593.540 14.320 1593.800 14.580 ;
        RECT 1626.200 14.320 1626.460 14.580 ;
      LAYER met2 ;
        RECT 1590.770 1700.000 1591.050 1704.000 ;
        RECT 1590.840 1684.690 1590.980 1700.000 ;
        RECT 1590.780 1684.370 1591.040 1684.690 ;
        RECT 1593.540 1684.370 1593.800 1684.690 ;
        RECT 1593.600 14.610 1593.740 1684.370 ;
        RECT 1593.540 14.290 1593.800 14.610 ;
        RECT 1626.200 14.290 1626.460 14.610 ;
        RECT 1626.260 2.400 1626.400 14.290 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1595.350 1685.620 1595.670 1685.680 ;
        RECT 1617.890 1685.620 1618.210 1685.680 ;
        RECT 1595.350 1685.480 1618.210 1685.620 ;
        RECT 1595.350 1685.420 1595.670 1685.480 ;
        RECT 1617.890 1685.420 1618.210 1685.480 ;
        RECT 1617.890 20.640 1618.210 20.700 ;
        RECT 1644.110 20.640 1644.430 20.700 ;
        RECT 1617.890 20.500 1644.430 20.640 ;
        RECT 1617.890 20.440 1618.210 20.500 ;
        RECT 1644.110 20.440 1644.430 20.500 ;
      LAYER via ;
        RECT 1595.380 1685.420 1595.640 1685.680 ;
        RECT 1617.920 1685.420 1618.180 1685.680 ;
        RECT 1617.920 20.440 1618.180 20.700 ;
        RECT 1644.140 20.440 1644.400 20.700 ;
      LAYER met2 ;
        RECT 1595.370 1700.000 1595.650 1704.000 ;
        RECT 1595.440 1685.710 1595.580 1700.000 ;
        RECT 1595.380 1685.390 1595.640 1685.710 ;
        RECT 1617.920 1685.390 1618.180 1685.710 ;
        RECT 1617.980 20.730 1618.120 1685.390 ;
        RECT 1617.920 20.410 1618.180 20.730 ;
        RECT 1644.140 20.410 1644.400 20.730 ;
        RECT 1644.200 2.400 1644.340 20.410 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1599.490 19.280 1599.810 19.340 ;
        RECT 1662.050 19.280 1662.370 19.340 ;
        RECT 1599.490 19.140 1662.370 19.280 ;
        RECT 1599.490 19.080 1599.810 19.140 ;
        RECT 1662.050 19.080 1662.370 19.140 ;
      LAYER via ;
        RECT 1599.520 19.080 1599.780 19.340 ;
        RECT 1662.080 19.080 1662.340 19.340 ;
      LAYER met2 ;
        RECT 1598.590 1700.410 1598.870 1704.000 ;
        RECT 1598.590 1700.270 1599.720 1700.410 ;
        RECT 1598.590 1700.000 1598.870 1700.270 ;
        RECT 1599.580 19.370 1599.720 1700.270 ;
        RECT 1599.520 19.050 1599.780 19.370 ;
        RECT 1662.080 19.050 1662.340 19.370 ;
        RECT 1662.140 2.400 1662.280 19.050 ;
=======
      LAYER li1 ;
        RECT 1652.925 14.025 1653.095 18.955 ;
      LAYER mcon ;
        RECT 1652.925 18.785 1653.095 18.955 ;
      LAYER met1 ;
        RECT 1600.410 1689.020 1600.730 1689.080 ;
        RECT 1611.450 1689.020 1611.770 1689.080 ;
        RECT 1600.410 1688.880 1611.770 1689.020 ;
        RECT 1600.410 1688.820 1600.730 1688.880 ;
        RECT 1611.450 1688.820 1611.770 1688.880 ;
        RECT 1652.865 18.940 1653.155 18.985 ;
        RECT 1645.120 18.800 1653.155 18.940 ;
        RECT 1611.450 18.600 1611.770 18.660 ;
        RECT 1645.120 18.600 1645.260 18.800 ;
        RECT 1652.865 18.755 1653.155 18.800 ;
        RECT 1611.450 18.460 1645.260 18.600 ;
        RECT 1611.450 18.400 1611.770 18.460 ;
        RECT 1652.865 14.180 1653.155 14.225 ;
        RECT 1662.050 14.180 1662.370 14.240 ;
        RECT 1652.865 14.040 1662.370 14.180 ;
        RECT 1652.865 13.995 1653.155 14.040 ;
        RECT 1662.050 13.980 1662.370 14.040 ;
      LAYER via ;
        RECT 1600.440 1688.820 1600.700 1689.080 ;
        RECT 1611.480 1688.820 1611.740 1689.080 ;
        RECT 1611.480 18.400 1611.740 18.660 ;
        RECT 1662.080 13.980 1662.340 14.240 ;
      LAYER met2 ;
        RECT 1600.430 1700.000 1600.710 1704.000 ;
        RECT 1600.500 1689.110 1600.640 1700.000 ;
        RECT 1600.440 1688.790 1600.700 1689.110 ;
        RECT 1611.480 1688.790 1611.740 1689.110 ;
        RECT 1611.540 18.690 1611.680 1688.790 ;
        RECT 1611.480 18.370 1611.740 18.690 ;
        RECT 1662.080 13.950 1662.340 14.270 ;
        RECT 1662.140 2.400 1662.280 13.950 ;
>>>>>>> re-updated local openlane
        RECT 1661.930 -4.800 1662.490 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 0.300 ;
=======
      LAYER met1 ;
        RECT 1603.170 1687.660 1603.490 1687.720 ;
        RECT 1673.090 1687.660 1673.410 1687.720 ;
        RECT 1603.170 1687.520 1673.410 1687.660 ;
        RECT 1603.170 1687.460 1603.490 1687.520 ;
        RECT 1673.090 1687.460 1673.410 1687.520 ;
        RECT 1673.090 20.640 1673.410 20.700 ;
        RECT 1679.530 20.640 1679.850 20.700 ;
        RECT 1673.090 20.500 1679.850 20.640 ;
        RECT 1673.090 20.440 1673.410 20.500 ;
        RECT 1679.530 20.440 1679.850 20.500 ;
      LAYER via ;
        RECT 1603.200 1687.460 1603.460 1687.720 ;
        RECT 1673.120 1687.460 1673.380 1687.720 ;
        RECT 1673.120 20.440 1673.380 20.700 ;
        RECT 1679.560 20.440 1679.820 20.700 ;
      LAYER met2 ;
        RECT 1603.190 1700.000 1603.470 1704.000 ;
        RECT 1603.260 1687.750 1603.400 1700.000 ;
        RECT 1603.200 1687.430 1603.460 1687.750 ;
        RECT 1673.120 1687.430 1673.380 1687.750 ;
        RECT 1673.180 20.730 1673.320 1687.430 ;
        RECT 1673.120 20.410 1673.380 20.730 ;
        RECT 1679.560 20.410 1679.820 20.730 ;
        RECT 1679.620 2.400 1679.760 20.410 ;
=======
      LAYER li1 ;
        RECT 1655.685 18.105 1656.775 18.275 ;
      LAYER mcon ;
        RECT 1656.605 18.105 1656.775 18.275 ;
      LAYER met1 ;
        RECT 1605.010 1686.640 1605.330 1686.700 ;
        RECT 1638.590 1686.640 1638.910 1686.700 ;
        RECT 1605.010 1686.500 1638.910 1686.640 ;
        RECT 1605.010 1686.440 1605.330 1686.500 ;
        RECT 1638.590 1686.440 1638.910 1686.500 ;
        RECT 1638.590 18.260 1638.910 18.320 ;
        RECT 1655.625 18.260 1655.915 18.305 ;
        RECT 1638.590 18.120 1655.915 18.260 ;
        RECT 1638.590 18.060 1638.910 18.120 ;
        RECT 1655.625 18.075 1655.915 18.120 ;
        RECT 1656.545 18.260 1656.835 18.305 ;
        RECT 1678.610 18.260 1678.930 18.320 ;
        RECT 1656.545 18.120 1678.930 18.260 ;
        RECT 1656.545 18.075 1656.835 18.120 ;
        RECT 1678.610 18.060 1678.930 18.120 ;
      LAYER via ;
        RECT 1605.040 1686.440 1605.300 1686.700 ;
        RECT 1638.620 1686.440 1638.880 1686.700 ;
        RECT 1638.620 18.060 1638.880 18.320 ;
        RECT 1678.640 18.060 1678.900 18.320 ;
      LAYER met2 ;
        RECT 1605.030 1700.000 1605.310 1704.000 ;
        RECT 1605.100 1686.730 1605.240 1700.000 ;
        RECT 1605.040 1686.410 1605.300 1686.730 ;
        RECT 1638.620 1686.410 1638.880 1686.730 ;
        RECT 1638.680 18.350 1638.820 1686.410 ;
        RECT 1678.700 18.630 1679.760 18.770 ;
        RECT 1678.700 18.350 1678.840 18.630 ;
        RECT 1638.620 18.030 1638.880 18.350 ;
        RECT 1678.640 18.030 1678.900 18.350 ;
        RECT 1679.620 2.400 1679.760 18.630 ;
>>>>>>> re-updated local openlane
        RECT 1679.410 -4.800 1679.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 0.300 ;
=======
      LAYER met1 ;
        RECT 1610.070 1684.600 1610.390 1684.660 ;
        RECT 1631.690 1684.600 1632.010 1684.660 ;
        RECT 1610.070 1684.460 1632.010 1684.600 ;
        RECT 1610.070 1684.400 1610.390 1684.460 ;
        RECT 1631.690 1684.400 1632.010 1684.460 ;
        RECT 1631.690 14.520 1632.010 14.580 ;
        RECT 1697.470 14.520 1697.790 14.580 ;
        RECT 1631.690 14.380 1697.790 14.520 ;
        RECT 1631.690 14.320 1632.010 14.380 ;
        RECT 1697.470 14.320 1697.790 14.380 ;
      LAYER via ;
        RECT 1610.100 1684.400 1610.360 1684.660 ;
        RECT 1631.720 1684.400 1631.980 1684.660 ;
        RECT 1631.720 14.320 1631.980 14.580 ;
        RECT 1697.500 14.320 1697.760 14.580 ;
      LAYER met2 ;
        RECT 1610.090 1700.000 1610.370 1704.000 ;
        RECT 1610.160 1684.690 1610.300 1700.000 ;
        RECT 1610.100 1684.370 1610.360 1684.690 ;
        RECT 1631.720 1684.370 1631.980 1684.690 ;
        RECT 1631.780 14.610 1631.920 1684.370 ;
        RECT 1631.720 14.290 1631.980 14.610 ;
        RECT 1697.500 14.290 1697.760 14.610 ;
        RECT 1697.560 2.400 1697.700 14.290 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 0.300 ;
=======
      LAYER met1 ;
        RECT 734.230 44.440 734.550 44.500 ;
        RECT 1347.870 44.440 1348.190 44.500 ;
        RECT 734.230 44.300 1348.190 44.440 ;
        RECT 734.230 44.240 734.550 44.300 ;
        RECT 1347.870 44.240 1348.190 44.300 ;
      LAYER via ;
        RECT 734.260 44.240 734.520 44.500 ;
        RECT 1347.900 44.240 1348.160 44.500 ;
      LAYER met2 ;
        RECT 1348.810 1700.410 1349.090 1704.000 ;
        RECT 1347.960 1700.270 1349.090 1700.410 ;
        RECT 1347.960 44.530 1348.100 1700.270 ;
        RECT 1348.810 1700.000 1349.090 1700.270 ;
        RECT 734.260 44.210 734.520 44.530 ;
        RECT 1347.900 44.210 1348.160 44.530 ;
        RECT 734.320 2.400 734.460 44.210 ;
        RECT 734.110 -4.800 734.670 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 0.300 ;
=======
      LAYER li1 ;
        RECT 1652.925 15.385 1653.095 16.575 ;
      LAYER mcon ;
        RECT 1652.925 16.405 1653.095 16.575 ;
      LAYER met1 ;
        RECT 1613.290 16.900 1613.610 16.960 ;
        RECT 1613.290 16.760 1620.880 16.900 ;
        RECT 1613.290 16.700 1613.610 16.760 ;
        RECT 1620.740 16.560 1620.880 16.760 ;
        RECT 1652.865 16.560 1653.155 16.605 ;
        RECT 1620.740 16.420 1653.155 16.560 ;
        RECT 1652.865 16.375 1653.155 16.420 ;
        RECT 1652.865 15.540 1653.155 15.585 ;
=======
      LAYER met1 ;
        RECT 1614.670 1684.260 1614.990 1684.320 ;
        RECT 1620.190 1684.260 1620.510 1684.320 ;
        RECT 1614.670 1684.120 1620.510 1684.260 ;
        RECT 1614.670 1684.060 1614.990 1684.120 ;
        RECT 1620.190 1684.060 1620.510 1684.120 ;
>>>>>>> re-updated local openlane
        RECT 1715.410 15.540 1715.730 15.600 ;
        RECT 1652.020 15.400 1715.730 15.540 ;
        RECT 1619.730 15.200 1620.050 15.260 ;
        RECT 1652.020 15.200 1652.160 15.400 ;
        RECT 1715.410 15.340 1715.730 15.400 ;
        RECT 1619.730 15.060 1652.160 15.200 ;
        RECT 1619.730 15.000 1620.050 15.060 ;
      LAYER via ;
        RECT 1614.700 1684.060 1614.960 1684.320 ;
        RECT 1620.220 1684.060 1620.480 1684.320 ;
        RECT 1619.760 15.000 1620.020 15.260 ;
        RECT 1715.440 15.340 1715.700 15.600 ;
      LAYER met2 ;
        RECT 1614.690 1700.000 1614.970 1704.000 ;
        RECT 1614.760 1684.350 1614.900 1700.000 ;
        RECT 1614.700 1684.030 1614.960 1684.350 ;
        RECT 1620.220 1684.030 1620.480 1684.350 ;
        RECT 1620.280 20.130 1620.420 1684.030 ;
        RECT 1619.820 19.990 1620.420 20.130 ;
        RECT 1619.820 15.290 1619.960 19.990 ;
        RECT 1715.440 15.310 1715.700 15.630 ;
        RECT 1619.760 14.970 1620.020 15.290 ;
        RECT 1715.500 2.400 1715.640 15.310 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 0.300 ;
=======
      LAYER met1 ;
        RECT 1617.890 1688.680 1618.210 1688.740 ;
        RECT 1620.190 1688.680 1620.510 1688.740 ;
        RECT 1617.890 1688.540 1620.510 1688.680 ;
        RECT 1617.890 1688.480 1618.210 1688.540 ;
        RECT 1620.190 1688.480 1620.510 1688.540 ;
        RECT 1619.730 14.860 1620.050 14.920 ;
        RECT 1733.350 14.860 1733.670 14.920 ;
        RECT 1619.730 14.720 1733.670 14.860 ;
        RECT 1619.730 14.660 1620.050 14.720 ;
        RECT 1733.350 14.660 1733.670 14.720 ;
      LAYER via ;
        RECT 1617.920 1688.480 1618.180 1688.740 ;
        RECT 1620.220 1688.480 1620.480 1688.740 ;
        RECT 1619.760 14.660 1620.020 14.920 ;
        RECT 1733.380 14.660 1733.640 14.920 ;
      LAYER met2 ;
        RECT 1617.910 1700.000 1618.190 1704.000 ;
        RECT 1617.980 1688.770 1618.120 1700.000 ;
        RECT 1617.920 1688.450 1618.180 1688.770 ;
        RECT 1620.220 1688.450 1620.480 1688.770 ;
        RECT 1620.280 20.130 1620.420 1688.450 ;
        RECT 1619.820 19.990 1620.420 20.130 ;
        RECT 1619.820 14.950 1619.960 19.990 ;
        RECT 1619.760 14.630 1620.020 14.950 ;
        RECT 1733.380 14.630 1733.640 14.950 ;
        RECT 1733.440 2.400 1733.580 14.630 ;
=======
      LAYER li1 ;
        RECT 1651.085 15.725 1651.255 16.575 ;
      LAYER mcon ;
        RECT 1651.085 16.405 1651.255 16.575 ;
      LAYER met1 ;
        RECT 1651.025 16.560 1651.315 16.605 ;
        RECT 1733.350 16.560 1733.670 16.620 ;
        RECT 1651.025 16.420 1733.670 16.560 ;
        RECT 1651.025 16.375 1651.315 16.420 ;
        RECT 1733.350 16.360 1733.670 16.420 ;
        RECT 1620.650 15.880 1620.970 15.940 ;
        RECT 1651.025 15.880 1651.315 15.925 ;
        RECT 1620.650 15.740 1651.315 15.880 ;
        RECT 1620.650 15.680 1620.970 15.740 ;
        RECT 1651.025 15.695 1651.315 15.740 ;
      LAYER via ;
        RECT 1733.380 16.360 1733.640 16.620 ;
        RECT 1620.680 15.680 1620.940 15.940 ;
      LAYER met2 ;
        RECT 1619.750 1700.410 1620.030 1704.000 ;
        RECT 1619.750 1700.270 1620.880 1700.410 ;
        RECT 1619.750 1700.000 1620.030 1700.270 ;
        RECT 1620.740 15.970 1620.880 1700.270 ;
        RECT 1733.380 16.330 1733.640 16.650 ;
        RECT 1620.680 15.650 1620.940 15.970 ;
        RECT 1733.440 2.400 1733.580 16.330 ;
>>>>>>> re-updated local openlane
        RECT 1733.230 -4.800 1733.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 0.300 ;
=======
      LAYER met1 ;
        RECT 1624.330 1683.920 1624.650 1683.980 ;
        RECT 1627.550 1683.920 1627.870 1683.980 ;
        RECT 1624.330 1683.780 1627.870 1683.920 ;
        RECT 1624.330 1683.720 1624.650 1683.780 ;
        RECT 1627.550 1683.720 1627.870 1683.780 ;
        RECT 1751.290 16.900 1751.610 16.960 ;
        RECT 1650.640 16.760 1751.610 16.900 ;
        RECT 1627.550 16.560 1627.870 16.620 ;
        RECT 1650.640 16.560 1650.780 16.760 ;
        RECT 1751.290 16.700 1751.610 16.760 ;
        RECT 1627.550 16.420 1650.780 16.560 ;
        RECT 1627.550 16.360 1627.870 16.420 ;
      LAYER via ;
        RECT 1624.360 1683.720 1624.620 1683.980 ;
        RECT 1627.580 1683.720 1627.840 1683.980 ;
        RECT 1627.580 16.360 1627.840 16.620 ;
        RECT 1751.320 16.700 1751.580 16.960 ;
      LAYER met2 ;
        RECT 1624.350 1700.000 1624.630 1704.000 ;
        RECT 1624.420 1684.010 1624.560 1700.000 ;
        RECT 1624.360 1683.690 1624.620 1684.010 ;
        RECT 1627.580 1683.690 1627.840 1684.010 ;
        RECT 1627.640 16.650 1627.780 1683.690 ;
        RECT 1751.320 16.670 1751.580 16.990 ;
        RECT 1627.580 16.330 1627.840 16.650 ;
        RECT 1751.380 2.400 1751.520 16.670 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 0.300 ;
=======
      LAYER met1 ;
        RECT 1629.390 1684.260 1629.710 1684.320 ;
        RECT 1633.990 1684.260 1634.310 1684.320 ;
        RECT 1629.390 1684.120 1634.310 1684.260 ;
        RECT 1629.390 1684.060 1629.710 1684.120 ;
        RECT 1633.990 1684.060 1634.310 1684.120 ;
        RECT 1633.990 20.300 1634.310 20.360 ;
        RECT 1768.770 20.300 1769.090 20.360 ;
        RECT 1633.990 20.160 1769.090 20.300 ;
        RECT 1633.990 20.100 1634.310 20.160 ;
        RECT 1768.770 20.100 1769.090 20.160 ;
      LAYER via ;
        RECT 1629.420 1684.060 1629.680 1684.320 ;
        RECT 1634.020 1684.060 1634.280 1684.320 ;
        RECT 1634.020 20.100 1634.280 20.360 ;
        RECT 1768.800 20.100 1769.060 20.360 ;
      LAYER met2 ;
        RECT 1629.410 1700.000 1629.690 1704.000 ;
        RECT 1629.480 1684.350 1629.620 1700.000 ;
        RECT 1629.420 1684.030 1629.680 1684.350 ;
        RECT 1634.020 1684.030 1634.280 1684.350 ;
        RECT 1634.080 20.390 1634.220 1684.030 ;
        RECT 1634.020 20.070 1634.280 20.390 ;
        RECT 1768.800 20.070 1769.060 20.390 ;
        RECT 1768.860 2.400 1769.000 20.070 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 0.300 ;
=======
      LAYER li1 ;
        RECT 1675.005 14.365 1675.175 19.975 ;
      LAYER mcon ;
        RECT 1675.005 19.805 1675.175 19.975 ;
      LAYER met1 ;
        RECT 1632.150 1688.680 1632.470 1688.740 ;
        RECT 1634.450 1688.680 1634.770 1688.740 ;
        RECT 1632.150 1688.540 1634.770 1688.680 ;
        RECT 1632.150 1688.480 1632.470 1688.540 ;
        RECT 1634.450 1688.480 1634.770 1688.540 ;
        RECT 1674.945 19.960 1675.235 20.005 ;
        RECT 1786.710 19.960 1787.030 20.020 ;
        RECT 1674.945 19.820 1787.030 19.960 ;
        RECT 1674.945 19.775 1675.235 19.820 ;
        RECT 1786.710 19.760 1787.030 19.820 ;
        RECT 1634.450 14.520 1634.770 14.580 ;
        RECT 1674.945 14.520 1675.235 14.565 ;
        RECT 1634.450 14.380 1675.235 14.520 ;
        RECT 1634.450 14.320 1634.770 14.380 ;
        RECT 1674.945 14.335 1675.235 14.380 ;
      LAYER via ;
        RECT 1632.180 1688.480 1632.440 1688.740 ;
        RECT 1634.480 1688.480 1634.740 1688.740 ;
        RECT 1786.740 19.760 1787.000 20.020 ;
        RECT 1634.480 14.320 1634.740 14.580 ;
      LAYER met2 ;
        RECT 1632.170 1700.000 1632.450 1704.000 ;
        RECT 1632.240 1688.770 1632.380 1700.000 ;
        RECT 1632.180 1688.450 1632.440 1688.770 ;
        RECT 1634.480 1688.450 1634.740 1688.770 ;
        RECT 1634.540 14.610 1634.680 1688.450 ;
        RECT 1786.740 19.730 1787.000 20.050 ;
        RECT 1634.480 14.290 1634.740 14.610 ;
        RECT 1786.800 2.400 1786.940 19.730 ;
=======
      LAYER met1 ;
        RECT 1634.450 19.620 1634.770 19.680 ;
        RECT 1786.710 19.620 1787.030 19.680 ;
        RECT 1634.450 19.480 1787.030 19.620 ;
        RECT 1634.450 19.420 1634.770 19.480 ;
        RECT 1786.710 19.420 1787.030 19.480 ;
      LAYER via ;
        RECT 1634.480 19.420 1634.740 19.680 ;
        RECT 1786.740 19.420 1787.000 19.680 ;
      LAYER met2 ;
        RECT 1634.010 1700.410 1634.290 1704.000 ;
        RECT 1634.010 1700.270 1634.680 1700.410 ;
        RECT 1634.010 1700.000 1634.290 1700.270 ;
        RECT 1634.540 19.710 1634.680 1700.270 ;
        RECT 1634.480 19.390 1634.740 19.710 ;
        RECT 1786.740 19.390 1787.000 19.710 ;
        RECT 1786.800 2.400 1786.940 19.390 ;
>>>>>>> re-updated local openlane
        RECT 1786.590 -4.800 1787.150 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 0.300 ;
=======
      LAYER li1 ;
        RECT 1641.425 1256.045 1641.595 1257.575 ;
        RECT 1662.585 16.065 1662.755 19.295 ;
      LAYER mcon ;
        RECT 1641.425 1257.405 1641.595 1257.575 ;
        RECT 1662.585 19.125 1662.755 19.295 ;
      LAYER met1 ;
        RECT 1637.210 1688.340 1637.530 1688.400 ;
        RECT 1641.350 1688.340 1641.670 1688.400 ;
        RECT 1637.210 1688.200 1641.670 1688.340 ;
        RECT 1637.210 1688.140 1637.530 1688.200 ;
        RECT 1641.350 1688.140 1641.670 1688.200 ;
        RECT 1641.350 1257.560 1641.670 1257.620 ;
        RECT 1641.155 1257.420 1641.670 1257.560 ;
        RECT 1641.350 1257.360 1641.670 1257.420 ;
        RECT 1641.350 1256.200 1641.670 1256.260 ;
        RECT 1641.155 1256.060 1641.670 1256.200 ;
        RECT 1641.350 1256.000 1641.670 1256.060 ;
        RECT 1641.350 435.920 1641.670 436.180 ;
        RECT 1641.440 435.160 1641.580 435.920 ;
        RECT 1641.350 434.900 1641.670 435.160 ;
        RECT 1641.350 146.240 1641.670 146.500 ;
        RECT 1641.440 145.140 1641.580 146.240 ;
        RECT 1641.350 144.880 1641.670 145.140 ;
        RECT 1662.525 19.280 1662.815 19.325 ;
=======
      LAYER met1 ;
        RECT 1639.050 1683.920 1639.370 1683.980 ;
        RECT 1641.810 1683.920 1642.130 1683.980 ;
        RECT 1639.050 1683.780 1642.130 1683.920 ;
        RECT 1639.050 1683.720 1639.370 1683.780 ;
        RECT 1641.810 1683.720 1642.130 1683.780 ;
        RECT 1641.810 19.280 1642.130 19.340 ;
>>>>>>> re-updated local openlane
        RECT 1804.650 19.280 1804.970 19.340 ;
        RECT 1641.810 19.140 1804.970 19.280 ;
        RECT 1641.810 19.080 1642.130 19.140 ;
        RECT 1804.650 19.080 1804.970 19.140 ;
      LAYER via ;
        RECT 1639.080 1683.720 1639.340 1683.980 ;
        RECT 1641.840 1683.720 1642.100 1683.980 ;
        RECT 1641.840 19.080 1642.100 19.340 ;
        RECT 1804.680 19.080 1804.940 19.340 ;
      LAYER met2 ;
        RECT 1639.070 1700.000 1639.350 1704.000 ;
        RECT 1639.140 1684.010 1639.280 1700.000 ;
        RECT 1639.080 1683.690 1639.340 1684.010 ;
        RECT 1641.840 1683.690 1642.100 1684.010 ;
        RECT 1641.900 19.370 1642.040 1683.690 ;
        RECT 1641.840 19.050 1642.100 19.370 ;
        RECT 1804.680 19.050 1804.940 19.370 ;
        RECT 1804.740 2.400 1804.880 19.050 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 0.300 ;
=======
      LAYER met1 ;
        RECT 1643.650 1684.600 1643.970 1684.660 ;
        RECT 1648.710 1684.600 1649.030 1684.660 ;
        RECT 1643.650 1684.460 1649.030 1684.600 ;
        RECT 1643.650 1684.400 1643.970 1684.460 ;
        RECT 1648.710 1684.400 1649.030 1684.460 ;
        RECT 1822.590 18.940 1822.910 19.000 ;
        RECT 1680.080 18.800 1822.910 18.940 ;
        RECT 1648.710 18.600 1649.030 18.660 ;
        RECT 1680.080 18.600 1680.220 18.800 ;
        RECT 1822.590 18.740 1822.910 18.800 ;
        RECT 1648.710 18.460 1680.220 18.600 ;
        RECT 1648.710 18.400 1649.030 18.460 ;
      LAYER via ;
        RECT 1643.680 1684.400 1643.940 1684.660 ;
        RECT 1648.740 1684.400 1649.000 1684.660 ;
        RECT 1648.740 18.400 1649.000 18.660 ;
        RECT 1822.620 18.740 1822.880 19.000 ;
      LAYER met2 ;
        RECT 1643.670 1700.000 1643.950 1704.000 ;
        RECT 1643.740 1684.690 1643.880 1700.000 ;
        RECT 1643.680 1684.370 1643.940 1684.690 ;
        RECT 1648.740 1684.370 1649.000 1684.690 ;
        RECT 1648.800 18.690 1648.940 1684.370 ;
        RECT 1822.620 18.710 1822.880 19.030 ;
        RECT 1648.740 18.370 1649.000 18.690 ;
        RECT 1822.680 2.400 1822.820 18.710 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1641.830 16.520 1642.110 16.800 ;
        RECT 1822.610 16.520 1822.890 16.800 ;
      LAYER met3 ;
        RECT 1641.805 16.810 1642.135 16.825 ;
        RECT 1822.585 16.810 1822.915 16.825 ;
        RECT 1641.805 16.510 1822.915 16.810 ;
        RECT 1641.805 16.495 1642.135 16.510 ;
        RECT 1822.585 16.495 1822.915 16.510 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 0.300 ;
=======
      LAYER li1 ;
        RECT 1700.765 17.425 1700.935 20.315 ;
        RECT 1820.365 17.425 1820.535 18.955 ;
      LAYER mcon ;
        RECT 1700.765 20.145 1700.935 20.315 ;
        RECT 1820.365 18.785 1820.535 18.955 ;
      LAYER met1 ;
        RECT 1646.870 1685.620 1647.190 1685.680 ;
        RECT 1648.710 1685.620 1649.030 1685.680 ;
        RECT 1646.870 1685.480 1649.030 1685.620 ;
        RECT 1646.870 1685.420 1647.190 1685.480 ;
        RECT 1648.710 1685.420 1649.030 1685.480 ;
        RECT 1700.705 20.300 1700.995 20.345 ;
        RECT 1674.560 20.160 1700.995 20.300 ;
        RECT 1648.710 19.960 1649.030 20.020 ;
        RECT 1674.560 19.960 1674.700 20.160 ;
        RECT 1700.705 20.115 1700.995 20.160 ;
        RECT 1648.710 19.820 1674.700 19.960 ;
        RECT 1648.710 19.760 1649.030 19.820 ;
        RECT 1820.305 18.940 1820.595 18.985 ;
        RECT 1840.070 18.940 1840.390 19.000 ;
        RECT 1820.305 18.800 1840.390 18.940 ;
        RECT 1820.305 18.755 1820.595 18.800 ;
        RECT 1840.070 18.740 1840.390 18.800 ;
        RECT 1700.705 17.580 1700.995 17.625 ;
        RECT 1820.305 17.580 1820.595 17.625 ;
        RECT 1700.705 17.440 1820.595 17.580 ;
        RECT 1700.705 17.395 1700.995 17.440 ;
        RECT 1820.305 17.395 1820.595 17.440 ;
      LAYER via ;
        RECT 1646.900 1685.420 1647.160 1685.680 ;
        RECT 1648.740 1685.420 1649.000 1685.680 ;
        RECT 1648.740 19.760 1649.000 20.020 ;
        RECT 1840.100 18.740 1840.360 19.000 ;
=======
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1648.730 1700.410 1649.010 1704.000 ;
        RECT 1648.340 1700.270 1649.010 1700.410 ;
        RECT 1648.340 16.845 1648.480 1700.270 ;
        RECT 1648.730 1700.000 1649.010 1700.270 ;
        RECT 1648.270 16.475 1648.550 16.845 ;
        RECT 1840.090 16.475 1840.370 16.845 ;
        RECT 1840.160 2.400 1840.300 16.475 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 1648.270 16.520 1648.550 16.800 ;
        RECT 1840.090 16.520 1840.370 16.800 ;
      LAYER met3 ;
        RECT 1648.245 16.810 1648.575 16.825 ;
        RECT 1840.065 16.810 1840.395 16.825 ;
        RECT 1648.245 16.510 1840.395 16.810 ;
        RECT 1648.245 16.495 1648.575 16.510 ;
        RECT 1840.065 16.495 1840.395 16.510 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 0.300 ;
=======
      LAYER met1 ;
        RECT 1651.470 1688.680 1651.790 1688.740 ;
        RECT 1655.610 1688.680 1655.930 1688.740 ;
        RECT 1651.470 1688.540 1655.930 1688.680 ;
        RECT 1651.470 1688.480 1651.790 1688.540 ;
        RECT 1655.610 1688.480 1655.930 1688.540 ;
        RECT 1655.610 17.240 1655.930 17.300 ;
        RECT 1858.010 17.240 1858.330 17.300 ;
        RECT 1655.610 17.100 1858.330 17.240 ;
        RECT 1655.610 17.040 1655.930 17.100 ;
        RECT 1858.010 17.040 1858.330 17.100 ;
      LAYER via ;
        RECT 1651.500 1688.480 1651.760 1688.740 ;
        RECT 1655.640 1688.480 1655.900 1688.740 ;
        RECT 1655.640 17.040 1655.900 17.300 ;
        RECT 1858.040 17.040 1858.300 17.300 ;
      LAYER met2 ;
        RECT 1651.490 1700.000 1651.770 1704.000 ;
        RECT 1651.560 1688.770 1651.700 1700.000 ;
        RECT 1651.500 1688.450 1651.760 1688.770 ;
        RECT 1655.640 1688.450 1655.900 1688.770 ;
        RECT 1655.700 17.330 1655.840 1688.450 ;
        RECT 1655.640 17.010 1655.900 17.330 ;
        RECT 1858.040 17.010 1858.300 17.330 ;
        RECT 1858.100 2.400 1858.240 17.010 ;
=======
      LAYER li1 ;
        RECT 1679.605 18.105 1679.775 18.955 ;
      LAYER mcon ;
        RECT 1679.605 18.785 1679.775 18.955 ;
      LAYER met1 ;
        RECT 1653.310 1683.920 1653.630 1683.980 ;
        RECT 1655.610 1683.920 1655.930 1683.980 ;
        RECT 1653.310 1683.780 1655.930 1683.920 ;
        RECT 1653.310 1683.720 1653.630 1683.780 ;
        RECT 1655.610 1683.720 1655.930 1683.780 ;
        RECT 1655.610 18.940 1655.930 19.000 ;
        RECT 1679.545 18.940 1679.835 18.985 ;
        RECT 1655.610 18.800 1679.835 18.940 ;
        RECT 1655.610 18.740 1655.930 18.800 ;
        RECT 1679.545 18.755 1679.835 18.800 ;
        RECT 1858.010 18.600 1858.330 18.660 ;
        RECT 1680.540 18.460 1858.330 18.600 ;
        RECT 1679.545 18.260 1679.835 18.305 ;
        RECT 1680.540 18.260 1680.680 18.460 ;
        RECT 1858.010 18.400 1858.330 18.460 ;
        RECT 1679.545 18.120 1680.680 18.260 ;
        RECT 1679.545 18.075 1679.835 18.120 ;
      LAYER via ;
        RECT 1653.340 1683.720 1653.600 1683.980 ;
        RECT 1655.640 1683.720 1655.900 1683.980 ;
        RECT 1655.640 18.740 1655.900 19.000 ;
        RECT 1858.040 18.400 1858.300 18.660 ;
      LAYER met2 ;
        RECT 1653.330 1700.000 1653.610 1704.000 ;
        RECT 1653.400 1684.010 1653.540 1700.000 ;
        RECT 1653.340 1683.690 1653.600 1684.010 ;
        RECT 1655.640 1683.690 1655.900 1684.010 ;
        RECT 1655.700 19.030 1655.840 1683.690 ;
        RECT 1655.640 18.710 1655.900 19.030 ;
        RECT 1858.040 18.370 1858.300 18.690 ;
        RECT 1858.100 2.400 1858.240 18.370 ;
>>>>>>> re-updated local openlane
        RECT 1857.890 -4.800 1858.450 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 0.300 ;
=======
      LAYER li1 ;
        RECT 1680.985 14.025 1681.155 18.275 ;
      LAYER mcon ;
        RECT 1680.985 18.105 1681.155 18.275 ;
      LAYER met1 ;
        RECT 1658.370 1684.600 1658.690 1684.660 ;
        RECT 1662.510 1684.600 1662.830 1684.660 ;
        RECT 1658.370 1684.460 1662.830 1684.600 ;
        RECT 1658.370 1684.400 1658.690 1684.460 ;
        RECT 1662.510 1684.400 1662.830 1684.460 ;
        RECT 1680.925 18.260 1681.215 18.305 ;
        RECT 1875.950 18.260 1876.270 18.320 ;
        RECT 1680.925 18.120 1876.270 18.260 ;
        RECT 1680.925 18.075 1681.215 18.120 ;
        RECT 1875.950 18.060 1876.270 18.120 ;
        RECT 1662.510 14.180 1662.830 14.240 ;
        RECT 1680.925 14.180 1681.215 14.225 ;
        RECT 1662.510 14.040 1681.215 14.180 ;
        RECT 1662.510 13.980 1662.830 14.040 ;
        RECT 1680.925 13.995 1681.215 14.040 ;
      LAYER via ;
        RECT 1658.400 1684.400 1658.660 1684.660 ;
        RECT 1662.540 1684.400 1662.800 1684.660 ;
        RECT 1875.980 18.060 1876.240 18.320 ;
        RECT 1662.540 13.980 1662.800 14.240 ;
      LAYER met2 ;
        RECT 1658.390 1700.000 1658.670 1704.000 ;
        RECT 1658.460 1684.690 1658.600 1700.000 ;
        RECT 1658.400 1684.370 1658.660 1684.690 ;
        RECT 1662.540 1684.370 1662.800 1684.690 ;
        RECT 1662.600 14.270 1662.740 1684.370 ;
        RECT 1875.980 18.030 1876.240 18.350 ;
        RECT 1662.540 13.950 1662.800 14.270 ;
        RECT 1876.040 2.400 1876.180 18.030 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 0.300 ;
=======
      LAYER met1 ;
        RECT 752.170 44.100 752.490 44.160 ;
        RECT 1353.390 44.100 1353.710 44.160 ;
        RECT 752.170 43.960 1353.710 44.100 ;
        RECT 752.170 43.900 752.490 43.960 ;
        RECT 1353.390 43.900 1353.710 43.960 ;
      LAYER via ;
        RECT 752.200 43.900 752.460 44.160 ;
        RECT 1353.420 43.900 1353.680 44.160 ;
      LAYER met2 ;
        RECT 1353.410 1700.000 1353.690 1704.000 ;
        RECT 1353.480 44.190 1353.620 1700.000 ;
        RECT 752.200 43.870 752.460 44.190 ;
        RECT 1353.420 43.870 1353.680 44.190 ;
        RECT 752.260 2.400 752.400 43.870 ;
        RECT 752.050 -4.800 752.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1662.970 1683.920 1663.290 1683.980 ;
        RECT 1662.970 1683.780 1667.800 1683.920 ;
        RECT 1662.970 1683.720 1663.290 1683.780 ;
        RECT 1667.660 1683.240 1667.800 1683.780 ;
        RECT 1669.410 1683.240 1669.730 1683.300 ;
        RECT 1667.660 1683.100 1669.730 1683.240 ;
        RECT 1669.410 1683.040 1669.730 1683.100 ;
        RECT 1669.410 17.920 1669.730 17.980 ;
        RECT 1893.890 17.920 1894.210 17.980 ;
        RECT 1669.410 17.780 1894.210 17.920 ;
        RECT 1669.410 17.720 1669.730 17.780 ;
        RECT 1893.890 17.720 1894.210 17.780 ;
      LAYER via ;
        RECT 1663.000 1683.720 1663.260 1683.980 ;
        RECT 1669.440 1683.040 1669.700 1683.300 ;
        RECT 1669.440 17.720 1669.700 17.980 ;
        RECT 1893.920 17.720 1894.180 17.980 ;
      LAYER met2 ;
        RECT 1662.990 1700.000 1663.270 1704.000 ;
        RECT 1663.060 1684.010 1663.200 1700.000 ;
        RECT 1663.000 1683.690 1663.260 1684.010 ;
        RECT 1669.440 1683.010 1669.700 1683.330 ;
        RECT 1669.500 18.010 1669.640 1683.010 ;
        RECT 1669.440 17.690 1669.700 18.010 ;
        RECT 1893.920 17.690 1894.180 18.010 ;
        RECT 1893.980 2.400 1894.120 17.690 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1668.950 17.580 1669.270 17.640 ;
        RECT 1911.830 17.580 1912.150 17.640 ;
        RECT 1668.950 17.440 1912.150 17.580 ;
        RECT 1668.950 17.380 1669.270 17.440 ;
        RECT 1911.830 17.380 1912.150 17.440 ;
      LAYER via ;
        RECT 1668.980 17.380 1669.240 17.640 ;
        RECT 1911.860 17.380 1912.120 17.640 ;
      LAYER met2 ;
        RECT 1668.050 1700.410 1668.330 1704.000 ;
        RECT 1668.050 1700.270 1669.180 1700.410 ;
        RECT 1668.050 1700.000 1668.330 1700.270 ;
        RECT 1669.040 17.670 1669.180 1700.270 ;
        RECT 1668.980 17.350 1669.240 17.670 ;
        RECT 1911.860 17.350 1912.120 17.670 ;
        RECT 1911.920 2.400 1912.060 17.350 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1672.630 1684.600 1672.950 1684.660 ;
        RECT 1676.310 1684.600 1676.630 1684.660 ;
        RECT 1672.630 1684.460 1676.630 1684.600 ;
        RECT 1672.630 1684.400 1672.950 1684.460 ;
        RECT 1676.310 1684.400 1676.630 1684.460 ;
        RECT 1676.310 17.240 1676.630 17.300 ;
        RECT 1929.310 17.240 1929.630 17.300 ;
        RECT 1676.310 17.100 1929.630 17.240 ;
        RECT 1676.310 17.040 1676.630 17.100 ;
        RECT 1929.310 17.040 1929.630 17.100 ;
      LAYER via ;
        RECT 1672.660 1684.400 1672.920 1684.660 ;
        RECT 1676.340 1684.400 1676.600 1684.660 ;
        RECT 1676.340 17.040 1676.600 17.300 ;
        RECT 1929.340 17.040 1929.600 17.300 ;
      LAYER met2 ;
        RECT 1672.650 1700.000 1672.930 1704.000 ;
        RECT 1672.720 1684.690 1672.860 1700.000 ;
        RECT 1672.660 1684.370 1672.920 1684.690 ;
        RECT 1676.340 1684.370 1676.600 1684.690 ;
        RECT 1676.400 17.330 1676.540 1684.370 ;
        RECT 1676.340 17.010 1676.600 17.330 ;
        RECT 1929.340 17.010 1929.600 17.330 ;
        RECT 1929.400 2.400 1929.540 17.010 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1947.130 -4.800 1947.690 0.300 ;
=======
        RECT 1675.410 1700.410 1675.690 1704.000 ;
        RECT 1675.410 1700.270 1676.080 1700.410 ;
        RECT 1675.410 1700.000 1675.690 1700.270 ;
        RECT 1675.940 15.485 1676.080 1700.270 ;
        RECT 1675.870 15.115 1676.150 15.485 ;
        RECT 1947.270 15.115 1947.550 15.485 ;
        RECT 1947.340 2.400 1947.480 15.115 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
      LAYER via2 ;
        RECT 1675.870 15.160 1676.150 15.440 ;
        RECT 1947.270 15.160 1947.550 15.440 ;
      LAYER met3 ;
        RECT 1675.845 15.450 1676.175 15.465 ;
        RECT 1947.245 15.450 1947.575 15.465 ;
        RECT 1675.845 15.150 1947.575 15.450 ;
        RECT 1675.845 15.135 1676.175 15.150 ;
        RECT 1947.245 15.135 1947.575 15.150 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1919.725 1684.785 1919.895 1685.635 ;
      LAYER mcon ;
        RECT 1919.725 1685.465 1919.895 1685.635 ;
      LAYER met1 ;
        RECT 1677.690 1685.620 1678.010 1685.680 ;
        RECT 1919.665 1685.620 1919.955 1685.665 ;
        RECT 1677.690 1685.480 1919.955 1685.620 ;
        RECT 1677.690 1685.420 1678.010 1685.480 ;
        RECT 1919.665 1685.435 1919.955 1685.480 ;
        RECT 1919.665 1684.940 1919.955 1684.985 ;
        RECT 1945.870 1684.940 1946.190 1685.000 ;
        RECT 1919.665 1684.800 1946.190 1684.940 ;
        RECT 1919.665 1684.755 1919.955 1684.800 ;
        RECT 1945.870 1684.740 1946.190 1684.800 ;
      LAYER via ;
        RECT 1677.720 1685.420 1677.980 1685.680 ;
        RECT 1945.900 1684.740 1946.160 1685.000 ;
      LAYER met2 ;
        RECT 1677.710 1700.000 1677.990 1704.000 ;
        RECT 1677.780 1685.710 1677.920 1700.000 ;
        RECT 1677.720 1685.390 1677.980 1685.710 ;
        RECT 1945.900 1684.710 1946.160 1685.030 ;
        RECT 1945.960 3.130 1946.100 1684.710 ;
        RECT 1945.960 2.990 1947.480 3.130 ;
        RECT 1947.340 2.400 1947.480 2.990 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 0.300 ;
=======
      LAYER li1 ;
        RECT 1699.385 14.025 1700.015 14.195 ;
        RECT 1699.845 13.685 1700.015 14.025 ;
      LAYER met1 ;
        RECT 1683.210 14.180 1683.530 14.240 ;
        RECT 1699.325 14.180 1699.615 14.225 ;
        RECT 1965.190 14.180 1965.510 14.240 ;
        RECT 1683.210 14.040 1699.615 14.180 ;
        RECT 1683.210 13.980 1683.530 14.040 ;
        RECT 1699.325 13.995 1699.615 14.040 ;
        RECT 1701.700 14.040 1965.510 14.180 ;
        RECT 1699.785 13.840 1700.075 13.885 ;
        RECT 1701.700 13.840 1701.840 14.040 ;
        RECT 1965.190 13.980 1965.510 14.040 ;
        RECT 1699.785 13.700 1701.840 13.840 ;
        RECT 1699.785 13.655 1700.075 13.700 ;
      LAYER via ;
        RECT 1683.240 13.980 1683.500 14.240 ;
        RECT 1965.220 13.980 1965.480 14.240 ;
      LAYER met2 ;
        RECT 1682.310 1700.410 1682.590 1704.000 ;
        RECT 1682.310 1700.270 1683.440 1700.410 ;
        RECT 1682.310 1700.000 1682.590 1700.270 ;
        RECT 1683.300 14.270 1683.440 1700.270 ;
        RECT 1683.240 13.950 1683.500 14.270 ;
        RECT 1965.220 13.950 1965.480 14.270 ;
        RECT 1965.280 2.400 1965.420 13.950 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1687.350 1685.960 1687.670 1686.020 ;
        RECT 1980.370 1685.960 1980.690 1686.020 ;
        RECT 1687.350 1685.820 1980.690 1685.960 ;
        RECT 1687.350 1685.760 1687.670 1685.820 ;
        RECT 1980.370 1685.760 1980.690 1685.820 ;
        RECT 1980.370 62.120 1980.690 62.180 ;
        RECT 1983.130 62.120 1983.450 62.180 ;
        RECT 1980.370 61.980 1983.450 62.120 ;
        RECT 1980.370 61.920 1980.690 61.980 ;
        RECT 1983.130 61.920 1983.450 61.980 ;
      LAYER via ;
        RECT 1687.380 1685.760 1687.640 1686.020 ;
        RECT 1980.400 1685.760 1980.660 1686.020 ;
        RECT 1980.400 61.920 1980.660 62.180 ;
        RECT 1983.160 61.920 1983.420 62.180 ;
      LAYER met2 ;
        RECT 1687.370 1700.000 1687.650 1704.000 ;
        RECT 1687.440 1686.050 1687.580 1700.000 ;
        RECT 1687.380 1685.730 1687.640 1686.050 ;
        RECT 1980.400 1685.730 1980.660 1686.050 ;
        RECT 1980.460 62.210 1980.600 1685.730 ;
        RECT 1980.400 61.890 1980.660 62.210 ;
        RECT 1983.160 61.890 1983.420 62.210 ;
        RECT 1983.220 2.400 1983.360 61.890 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2000.950 -4.800 2001.510 0.300 ;
=======
        RECT 1690.130 1700.000 1690.410 1704.000 ;
        RECT 1690.200 16.165 1690.340 1700.000 ;
        RECT 1690.130 15.795 1690.410 16.165 ;
        RECT 2001.090 15.795 2001.370 16.165 ;
        RECT 2001.160 2.400 2001.300 15.795 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
      LAYER via2 ;
        RECT 1690.130 15.840 1690.410 16.120 ;
        RECT 2001.090 15.840 2001.370 16.120 ;
      LAYER met3 ;
        RECT 1690.105 16.130 1690.435 16.145 ;
        RECT 2001.065 16.130 2001.395 16.145 ;
        RECT 1690.105 15.830 2001.395 16.130 ;
        RECT 1690.105 15.815 1690.435 15.830 ;
        RECT 2001.065 15.815 2001.395 15.830 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1692.410 1684.260 1692.730 1684.320 ;
        RECT 1697.010 1684.260 1697.330 1684.320 ;
        RECT 1692.410 1684.120 1697.330 1684.260 ;
        RECT 1692.410 1684.060 1692.730 1684.120 ;
        RECT 1697.010 1684.060 1697.330 1684.120 ;
        RECT 1697.010 14.860 1697.330 14.920 ;
        RECT 1697.010 14.720 1698.160 14.860 ;
        RECT 1697.010 14.660 1697.330 14.720 ;
        RECT 1698.020 14.520 1698.160 14.720 ;
        RECT 2001.070 14.520 2001.390 14.580 ;
        RECT 1698.020 14.380 2001.390 14.520 ;
        RECT 2001.070 14.320 2001.390 14.380 ;
      LAYER via ;
        RECT 1692.440 1684.060 1692.700 1684.320 ;
        RECT 1697.040 1684.060 1697.300 1684.320 ;
        RECT 1697.040 14.660 1697.300 14.920 ;
        RECT 2001.100 14.320 2001.360 14.580 ;
      LAYER met2 ;
        RECT 1692.430 1700.000 1692.710 1704.000 ;
        RECT 1692.500 1684.350 1692.640 1700.000 ;
        RECT 1692.440 1684.030 1692.700 1684.350 ;
        RECT 1697.040 1684.030 1697.300 1684.350 ;
        RECT 1697.100 14.950 1697.240 1684.030 ;
        RECT 1697.040 14.630 1697.300 14.950 ;
        RECT 2001.100 14.290 2001.360 14.610 ;
        RECT 2001.160 2.400 2001.300 14.290 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 0.300 ;
=======
      LAYER met1 ;
        RECT 1694.710 1685.960 1695.030 1686.020 ;
        RECT 1697.010 1685.960 1697.330 1686.020 ;
        RECT 1694.710 1685.820 1697.330 1685.960 ;
        RECT 1694.710 1685.760 1695.030 1685.820 ;
        RECT 1697.010 1685.760 1697.330 1685.820 ;
      LAYER via ;
        RECT 1694.740 1685.760 1695.000 1686.020 ;
        RECT 1697.040 1685.760 1697.300 1686.020 ;
      LAYER met2 ;
        RECT 1694.730 1700.000 1695.010 1704.000 ;
        RECT 1694.800 1686.050 1694.940 1700.000 ;
        RECT 1694.740 1685.730 1695.000 1686.050 ;
        RECT 1697.040 1685.730 1697.300 1686.050 ;
        RECT 1697.100 20.245 1697.240 1685.730 ;
        RECT 1697.030 19.875 1697.310 20.245 ;
        RECT 2018.570 19.875 2018.850 20.245 ;
        RECT 2018.640 2.400 2018.780 19.875 ;
=======
      LAYER li1 ;
        RECT 2014.945 1635.485 2015.115 1683.595 ;
        RECT 2014.945 1538.925 2015.115 1587.035 ;
        RECT 2014.945 1442.025 2015.115 1490.475 ;
        RECT 2014.945 766.105 2015.115 814.215 ;
        RECT 2014.945 669.545 2015.115 717.655 ;
        RECT 2014.945 572.645 2015.115 620.755 ;
        RECT 2014.945 476.085 2015.115 524.195 ;
        RECT 2014.945 379.525 2015.115 427.635 ;
        RECT 2014.945 282.965 2015.115 331.075 ;
        RECT 2014.945 186.405 2015.115 234.515 ;
      LAYER mcon ;
        RECT 2014.945 1683.425 2015.115 1683.595 ;
        RECT 2014.945 1586.865 2015.115 1587.035 ;
        RECT 2014.945 1490.305 2015.115 1490.475 ;
        RECT 2014.945 814.045 2015.115 814.215 ;
        RECT 2014.945 717.485 2015.115 717.655 ;
        RECT 2014.945 620.585 2015.115 620.755 ;
        RECT 2014.945 524.025 2015.115 524.195 ;
        RECT 2014.945 427.465 2015.115 427.635 ;
        RECT 2014.945 330.905 2015.115 331.075 ;
        RECT 2014.945 234.345 2015.115 234.515 ;
      LAYER met1 ;
        RECT 1697.010 1686.300 1697.330 1686.360 ;
        RECT 2014.870 1686.300 2015.190 1686.360 ;
        RECT 1697.010 1686.160 2015.190 1686.300 ;
        RECT 1697.010 1686.100 1697.330 1686.160 ;
        RECT 2014.870 1686.100 2015.190 1686.160 ;
        RECT 2014.870 1683.580 2015.190 1683.640 ;
        RECT 2014.675 1683.440 2015.190 1683.580 ;
        RECT 2014.870 1683.380 2015.190 1683.440 ;
        RECT 2014.870 1635.640 2015.190 1635.700 ;
        RECT 2014.675 1635.500 2015.190 1635.640 ;
        RECT 2014.870 1635.440 2015.190 1635.500 ;
        RECT 2014.870 1587.020 2015.190 1587.080 ;
        RECT 2014.675 1586.880 2015.190 1587.020 ;
        RECT 2014.870 1586.820 2015.190 1586.880 ;
        RECT 2014.870 1539.080 2015.190 1539.140 ;
        RECT 2014.675 1538.940 2015.190 1539.080 ;
        RECT 2014.870 1538.880 2015.190 1538.940 ;
        RECT 2014.870 1490.460 2015.190 1490.520 ;
        RECT 2014.675 1490.320 2015.190 1490.460 ;
        RECT 2014.870 1490.260 2015.190 1490.320 ;
        RECT 2014.870 1442.180 2015.190 1442.240 ;
        RECT 2014.675 1442.040 2015.190 1442.180 ;
        RECT 2014.870 1441.980 2015.190 1442.040 ;
        RECT 2014.870 1007.320 2015.190 1007.380 ;
        RECT 2015.790 1007.320 2016.110 1007.380 ;
        RECT 2014.870 1007.180 2016.110 1007.320 ;
        RECT 2014.870 1007.120 2015.190 1007.180 ;
        RECT 2015.790 1007.120 2016.110 1007.180 ;
        RECT 2014.410 821.340 2014.730 821.400 ;
        RECT 2014.870 821.340 2015.190 821.400 ;
        RECT 2014.410 821.200 2015.190 821.340 ;
        RECT 2014.410 821.140 2014.730 821.200 ;
        RECT 2014.870 821.140 2015.190 821.200 ;
        RECT 2014.870 814.200 2015.190 814.260 ;
        RECT 2014.675 814.060 2015.190 814.200 ;
        RECT 2014.870 814.000 2015.190 814.060 ;
        RECT 2014.870 766.260 2015.190 766.320 ;
        RECT 2014.675 766.120 2015.190 766.260 ;
        RECT 2014.870 766.060 2015.190 766.120 ;
        RECT 2014.870 717.640 2015.190 717.700 ;
        RECT 2014.675 717.500 2015.190 717.640 ;
        RECT 2014.870 717.440 2015.190 717.500 ;
        RECT 2014.870 669.700 2015.190 669.760 ;
        RECT 2014.675 669.560 2015.190 669.700 ;
        RECT 2014.870 669.500 2015.190 669.560 ;
        RECT 2014.870 620.740 2015.190 620.800 ;
        RECT 2014.675 620.600 2015.190 620.740 ;
        RECT 2014.870 620.540 2015.190 620.600 ;
        RECT 2014.870 572.800 2015.190 572.860 ;
        RECT 2014.675 572.660 2015.190 572.800 ;
        RECT 2014.870 572.600 2015.190 572.660 ;
        RECT 2014.870 524.180 2015.190 524.240 ;
        RECT 2014.675 524.040 2015.190 524.180 ;
        RECT 2014.870 523.980 2015.190 524.040 ;
        RECT 2014.870 476.240 2015.190 476.300 ;
        RECT 2014.675 476.100 2015.190 476.240 ;
        RECT 2014.870 476.040 2015.190 476.100 ;
        RECT 2014.870 427.620 2015.190 427.680 ;
        RECT 2014.675 427.480 2015.190 427.620 ;
        RECT 2014.870 427.420 2015.190 427.480 ;
        RECT 2014.870 379.680 2015.190 379.740 ;
        RECT 2014.675 379.540 2015.190 379.680 ;
        RECT 2014.870 379.480 2015.190 379.540 ;
        RECT 2014.870 331.060 2015.190 331.120 ;
        RECT 2014.675 330.920 2015.190 331.060 ;
        RECT 2014.870 330.860 2015.190 330.920 ;
        RECT 2014.870 283.120 2015.190 283.180 ;
        RECT 2014.675 282.980 2015.190 283.120 ;
        RECT 2014.870 282.920 2015.190 282.980 ;
        RECT 2014.870 234.500 2015.190 234.560 ;
        RECT 2014.675 234.360 2015.190 234.500 ;
        RECT 2014.870 234.300 2015.190 234.360 ;
        RECT 2014.870 186.560 2015.190 186.620 ;
        RECT 2014.675 186.420 2015.190 186.560 ;
        RECT 2014.870 186.360 2015.190 186.420 ;
        RECT 2014.870 137.940 2015.190 138.000 ;
        RECT 2018.550 137.940 2018.870 138.000 ;
        RECT 2014.870 137.800 2018.870 137.940 ;
        RECT 2014.870 137.740 2015.190 137.800 ;
        RECT 2018.550 137.740 2018.870 137.800 ;
      LAYER via ;
        RECT 1697.040 1686.100 1697.300 1686.360 ;
        RECT 2014.900 1686.100 2015.160 1686.360 ;
        RECT 2014.900 1683.380 2015.160 1683.640 ;
        RECT 2014.900 1635.440 2015.160 1635.700 ;
        RECT 2014.900 1586.820 2015.160 1587.080 ;
        RECT 2014.900 1538.880 2015.160 1539.140 ;
        RECT 2014.900 1490.260 2015.160 1490.520 ;
        RECT 2014.900 1441.980 2015.160 1442.240 ;
        RECT 2014.900 1007.120 2015.160 1007.380 ;
        RECT 2015.820 1007.120 2016.080 1007.380 ;
        RECT 2014.440 821.140 2014.700 821.400 ;
        RECT 2014.900 821.140 2015.160 821.400 ;
        RECT 2014.900 814.000 2015.160 814.260 ;
        RECT 2014.900 766.060 2015.160 766.320 ;
        RECT 2014.900 717.440 2015.160 717.700 ;
        RECT 2014.900 669.500 2015.160 669.760 ;
        RECT 2014.900 620.540 2015.160 620.800 ;
        RECT 2014.900 572.600 2015.160 572.860 ;
        RECT 2014.900 523.980 2015.160 524.240 ;
        RECT 2014.900 476.040 2015.160 476.300 ;
        RECT 2014.900 427.420 2015.160 427.680 ;
        RECT 2014.900 379.480 2015.160 379.740 ;
        RECT 2014.900 330.860 2015.160 331.120 ;
        RECT 2014.900 282.920 2015.160 283.180 ;
        RECT 2014.900 234.300 2015.160 234.560 ;
        RECT 2014.900 186.360 2015.160 186.620 ;
        RECT 2014.900 137.740 2015.160 138.000 ;
        RECT 2018.580 137.740 2018.840 138.000 ;
      LAYER met2 ;
        RECT 1697.030 1700.000 1697.310 1704.000 ;
        RECT 1697.100 1686.390 1697.240 1700.000 ;
        RECT 1697.040 1686.070 1697.300 1686.390 ;
        RECT 2014.900 1686.070 2015.160 1686.390 ;
        RECT 2014.960 1683.670 2015.100 1686.070 ;
        RECT 2014.900 1683.350 2015.160 1683.670 ;
        RECT 2014.900 1635.410 2015.160 1635.730 ;
        RECT 2014.960 1587.110 2015.100 1635.410 ;
        RECT 2014.900 1586.790 2015.160 1587.110 ;
        RECT 2014.900 1538.850 2015.160 1539.170 ;
        RECT 2014.960 1490.550 2015.100 1538.850 ;
        RECT 2014.900 1490.230 2015.160 1490.550 ;
        RECT 2014.900 1441.950 2015.160 1442.270 ;
        RECT 2014.960 1007.410 2015.100 1441.950 ;
        RECT 2014.900 1007.090 2015.160 1007.410 ;
        RECT 2015.820 1007.090 2016.080 1007.410 ;
        RECT 2015.880 959.325 2016.020 1007.090 ;
        RECT 2014.890 958.955 2015.170 959.325 ;
        RECT 2015.810 958.955 2016.090 959.325 ;
        RECT 2014.960 869.450 2015.100 958.955 ;
        RECT 2014.500 869.310 2015.100 869.450 ;
        RECT 2014.500 821.430 2014.640 869.310 ;
        RECT 2014.440 821.110 2014.700 821.430 ;
        RECT 2014.900 821.110 2015.160 821.430 ;
        RECT 2014.960 814.290 2015.100 821.110 ;
        RECT 2014.900 813.970 2015.160 814.290 ;
        RECT 2014.900 766.030 2015.160 766.350 ;
        RECT 2014.960 717.730 2015.100 766.030 ;
        RECT 2014.900 717.410 2015.160 717.730 ;
        RECT 2014.900 669.470 2015.160 669.790 ;
        RECT 2014.960 620.830 2015.100 669.470 ;
        RECT 2014.900 620.510 2015.160 620.830 ;
        RECT 2014.900 572.570 2015.160 572.890 ;
        RECT 2014.960 524.270 2015.100 572.570 ;
        RECT 2014.900 523.950 2015.160 524.270 ;
        RECT 2014.900 476.010 2015.160 476.330 ;
        RECT 2014.960 427.710 2015.100 476.010 ;
        RECT 2014.900 427.390 2015.160 427.710 ;
        RECT 2014.900 379.450 2015.160 379.770 ;
        RECT 2014.960 331.150 2015.100 379.450 ;
        RECT 2014.900 330.830 2015.160 331.150 ;
        RECT 2014.900 282.890 2015.160 283.210 ;
        RECT 2014.960 234.590 2015.100 282.890 ;
        RECT 2014.900 234.270 2015.160 234.590 ;
        RECT 2014.900 186.330 2015.160 186.650 ;
        RECT 2014.960 138.030 2015.100 186.330 ;
        RECT 2014.900 137.710 2015.160 138.030 ;
        RECT 2018.580 137.710 2018.840 138.030 ;
        RECT 2018.640 2.400 2018.780 137.710 ;
>>>>>>> re-updated local openlane
        RECT 2018.430 -4.800 2018.990 2.400 ;
      LAYER via2 ;
        RECT 2014.890 959.000 2015.170 959.280 ;
        RECT 2015.810 959.000 2016.090 959.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1697.005 20.210 1697.335 20.225 ;
        RECT 2018.545 20.210 2018.875 20.225 ;
        RECT 1697.005 19.910 2018.875 20.210 ;
        RECT 1697.005 19.895 1697.335 19.910 ;
        RECT 2018.545 19.895 2018.875 19.910 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 2014.865 959.290 2015.195 959.305 ;
        RECT 2015.785 959.290 2016.115 959.305 ;
        RECT 2014.865 958.990 2016.115 959.290 ;
        RECT 2014.865 958.975 2015.195 958.990 ;
        RECT 2015.785 958.975 2016.115 958.990 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1702.530 14.860 1702.850 14.920 ;
        RECT 2036.490 14.860 2036.810 14.920 ;
        RECT 1702.530 14.720 2036.810 14.860 ;
        RECT 1702.530 14.660 1702.850 14.720 ;
        RECT 2036.490 14.660 2036.810 14.720 ;
      LAYER via ;
        RECT 1702.560 14.660 1702.820 14.920 ;
        RECT 2036.520 14.660 2036.780 14.920 ;
      LAYER met2 ;
        RECT 1702.090 1700.410 1702.370 1704.000 ;
        RECT 1702.090 1700.270 1702.760 1700.410 ;
        RECT 1702.090 1700.000 1702.370 1700.270 ;
        RECT 1702.620 14.950 1702.760 1700.270 ;
        RECT 1702.560 14.630 1702.820 14.950 ;
        RECT 2036.520 14.630 2036.780 14.950 ;
        RECT 2036.580 2.400 2036.720 14.630 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 0.300 ;
=======
      LAYER li1 ;
        RECT 1725.145 14.025 1725.315 18.955 ;
        RECT 1772.985 14.875 1773.155 18.955 ;
        RECT 1773.445 15.725 1773.615 18.955 ;
        RECT 1785.865 15.725 1786.035 16.915 ;
        RECT 1797.365 16.745 1797.535 19.975 ;
        RECT 1824.965 17.425 1825.135 19.975 ;
        RECT 1873.265 17.425 1873.435 18.955 ;
        RECT 1918.345 16.065 1918.515 18.955 ;
        RECT 1966.185 16.065 1966.355 18.955 ;
        RECT 2028.285 18.615 2028.455 18.955 ;
        RECT 2029.205 18.615 2029.375 20.315 ;
        RECT 2028.285 18.445 2029.375 18.615 ;
        RECT 1772.525 14.705 1773.155 14.875 ;
      LAYER mcon ;
        RECT 2029.205 20.145 2029.375 20.315 ;
        RECT 1797.365 19.805 1797.535 19.975 ;
        RECT 1725.145 18.785 1725.315 18.955 ;
        RECT 1772.985 18.785 1773.155 18.955 ;
        RECT 1773.445 18.785 1773.615 18.955 ;
        RECT 1824.965 19.805 1825.135 19.975 ;
        RECT 1873.265 18.785 1873.435 18.955 ;
        RECT 1918.345 18.785 1918.515 18.955 ;
        RECT 1785.865 16.745 1786.035 16.915 ;
        RECT 1966.185 18.785 1966.355 18.955 ;
        RECT 2028.285 18.785 2028.455 18.955 ;
      LAYER met1 ;
        RECT 1704.370 1688.680 1704.690 1688.740 ;
        RECT 1710.350 1688.680 1710.670 1688.740 ;
        RECT 1704.370 1688.540 1710.670 1688.680 ;
        RECT 1704.370 1688.480 1704.690 1688.540 ;
        RECT 1710.350 1688.480 1710.670 1688.540 ;
        RECT 2029.145 20.300 2029.435 20.345 ;
        RECT 2054.430 20.300 2054.750 20.360 ;
        RECT 2029.145 20.160 2054.750 20.300 ;
        RECT 2029.145 20.115 2029.435 20.160 ;
        RECT 2054.430 20.100 2054.750 20.160 ;
        RECT 1797.305 19.960 1797.595 20.005 ;
        RECT 1824.905 19.960 1825.195 20.005 ;
        RECT 1797.305 19.820 1825.195 19.960 ;
        RECT 1797.305 19.775 1797.595 19.820 ;
        RECT 1824.905 19.775 1825.195 19.820 ;
        RECT 1710.350 18.940 1710.670 19.000 ;
        RECT 1725.085 18.940 1725.375 18.985 ;
        RECT 1710.350 18.800 1725.375 18.940 ;
        RECT 1710.350 18.740 1710.670 18.800 ;
        RECT 1725.085 18.755 1725.375 18.800 ;
        RECT 1772.925 18.940 1773.215 18.985 ;
        RECT 1773.385 18.940 1773.675 18.985 ;
        RECT 1772.925 18.800 1773.675 18.940 ;
        RECT 1772.925 18.755 1773.215 18.800 ;
        RECT 1773.385 18.755 1773.675 18.800 ;
        RECT 1873.205 18.940 1873.495 18.985 ;
        RECT 1918.285 18.940 1918.575 18.985 ;
        RECT 1873.205 18.800 1918.575 18.940 ;
        RECT 1873.205 18.755 1873.495 18.800 ;
        RECT 1918.285 18.755 1918.575 18.800 ;
        RECT 1966.125 18.940 1966.415 18.985 ;
        RECT 2028.225 18.940 2028.515 18.985 ;
        RECT 1966.125 18.800 2028.515 18.940 ;
        RECT 1966.125 18.755 1966.415 18.800 ;
        RECT 2028.225 18.755 2028.515 18.800 ;
        RECT 1824.905 17.580 1825.195 17.625 ;
        RECT 1873.205 17.580 1873.495 17.625 ;
        RECT 1824.905 17.440 1873.495 17.580 ;
        RECT 1824.905 17.395 1825.195 17.440 ;
        RECT 1873.205 17.395 1873.495 17.440 ;
        RECT 1785.805 16.900 1786.095 16.945 ;
        RECT 1797.305 16.900 1797.595 16.945 ;
        RECT 1785.805 16.760 1797.595 16.900 ;
        RECT 1785.805 16.715 1786.095 16.760 ;
        RECT 1797.305 16.715 1797.595 16.760 ;
        RECT 1918.285 16.220 1918.575 16.265 ;
        RECT 1966.125 16.220 1966.415 16.265 ;
        RECT 1918.285 16.080 1966.415 16.220 ;
        RECT 1918.285 16.035 1918.575 16.080 ;
        RECT 1966.125 16.035 1966.415 16.080 ;
        RECT 1773.385 15.880 1773.675 15.925 ;
        RECT 1785.805 15.880 1786.095 15.925 ;
        RECT 1773.385 15.740 1786.095 15.880 ;
        RECT 1773.385 15.695 1773.675 15.740 ;
        RECT 1785.805 15.695 1786.095 15.740 ;
        RECT 1772.465 14.860 1772.755 14.905 ;
        RECT 1733.900 14.720 1772.755 14.860 ;
        RECT 1725.085 14.180 1725.375 14.225 ;
        RECT 1733.900 14.180 1734.040 14.720 ;
        RECT 1772.465 14.675 1772.755 14.720 ;
        RECT 1725.085 14.040 1734.040 14.180 ;
        RECT 1725.085 13.995 1725.375 14.040 ;
      LAYER via ;
        RECT 1704.400 1688.480 1704.660 1688.740 ;
        RECT 1710.380 1688.480 1710.640 1688.740 ;
        RECT 2054.460 20.100 2054.720 20.360 ;
        RECT 1710.380 18.740 1710.640 19.000 ;
      LAYER met2 ;
        RECT 1704.390 1700.000 1704.670 1704.000 ;
        RECT 1704.460 1688.770 1704.600 1700.000 ;
        RECT 1704.400 1688.450 1704.660 1688.770 ;
        RECT 1710.380 1688.450 1710.640 1688.770 ;
        RECT 1710.440 19.030 1710.580 1688.450 ;
        RECT 2054.460 20.070 2054.720 20.390 ;
        RECT 1710.380 18.710 1710.640 19.030 ;
        RECT 2054.520 2.400 2054.660 20.070 ;
=======
      LAYER met1 ;
        RECT 1706.670 1686.640 1706.990 1686.700 ;
        RECT 2049.370 1686.640 2049.690 1686.700 ;
        RECT 1706.670 1686.500 2049.690 1686.640 ;
        RECT 1706.670 1686.440 1706.990 1686.500 ;
        RECT 2049.370 1686.440 2049.690 1686.500 ;
        RECT 2049.370 62.120 2049.690 62.180 ;
        RECT 2054.430 62.120 2054.750 62.180 ;
        RECT 2049.370 61.980 2054.750 62.120 ;
        RECT 2049.370 61.920 2049.690 61.980 ;
        RECT 2054.430 61.920 2054.750 61.980 ;
      LAYER via ;
        RECT 1706.700 1686.440 1706.960 1686.700 ;
        RECT 2049.400 1686.440 2049.660 1686.700 ;
        RECT 2049.400 61.920 2049.660 62.180 ;
        RECT 2054.460 61.920 2054.720 62.180 ;
      LAYER met2 ;
        RECT 1706.690 1700.000 1706.970 1704.000 ;
        RECT 1706.760 1686.730 1706.900 1700.000 ;
        RECT 1706.700 1686.410 1706.960 1686.730 ;
        RECT 2049.400 1686.410 2049.660 1686.730 ;
        RECT 2049.460 62.210 2049.600 1686.410 ;
        RECT 2049.400 61.890 2049.660 62.210 ;
        RECT 2054.460 61.890 2054.720 62.210 ;
        RECT 2054.520 2.400 2054.660 61.890 ;
>>>>>>> re-updated local openlane
        RECT 2054.310 -4.800 2054.870 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1352.930 1678.140 1353.250 1678.200 ;
        RECT 1357.070 1678.140 1357.390 1678.200 ;
        RECT 1352.930 1678.000 1357.390 1678.140 ;
        RECT 1352.930 1677.940 1353.250 1678.000 ;
        RECT 1357.070 1677.940 1357.390 1678.000 ;
        RECT 769.650 43.760 769.970 43.820 ;
        RECT 1352.930 43.760 1353.250 43.820 ;
        RECT 769.650 43.620 1353.250 43.760 ;
        RECT 769.650 43.560 769.970 43.620 ;
        RECT 1352.930 43.560 1353.250 43.620 ;
      LAYER via ;
        RECT 1352.960 1677.940 1353.220 1678.200 ;
        RECT 1357.100 1677.940 1357.360 1678.200 ;
        RECT 769.680 43.560 769.940 43.820 ;
        RECT 1352.960 43.560 1353.220 43.820 ;
      LAYER met2 ;
        RECT 1358.470 1700.410 1358.750 1704.000 ;
        RECT 1357.160 1700.270 1358.750 1700.410 ;
        RECT 1357.160 1678.230 1357.300 1700.270 ;
        RECT 1358.470 1700.000 1358.750 1700.270 ;
        RECT 1352.960 1677.910 1353.220 1678.230 ;
        RECT 1357.100 1677.910 1357.360 1678.230 ;
        RECT 1353.020 43.850 1353.160 1677.910 ;
        RECT 769.680 43.530 769.940 43.850 ;
        RECT 1352.960 43.530 1353.220 43.850 ;
        RECT 769.740 2.400 769.880 43.530 ;
        RECT 769.530 -4.800 770.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 0.300 ;
=======
      LAYER li1 ;
        RECT 2038.865 16.405 2039.035 18.615 ;
      LAYER mcon ;
        RECT 2038.865 18.445 2039.035 18.615 ;
      LAYER met1 ;
        RECT 1709.430 1689.360 1709.750 1689.420 ;
        RECT 1710.810 1689.360 1711.130 1689.420 ;
        RECT 1709.430 1689.220 1711.130 1689.360 ;
        RECT 1709.430 1689.160 1709.750 1689.220 ;
        RECT 1710.810 1689.160 1711.130 1689.220 ;
        RECT 1710.810 18.600 1711.130 18.660 ;
        RECT 2038.805 18.600 2039.095 18.645 ;
        RECT 1710.810 18.460 2039.095 18.600 ;
        RECT 1710.810 18.400 1711.130 18.460 ;
        RECT 2038.805 18.415 2039.095 18.460 ;
        RECT 2038.805 16.560 2039.095 16.605 ;
        RECT 2072.370 16.560 2072.690 16.620 ;
        RECT 2038.805 16.420 2072.690 16.560 ;
        RECT 2038.805 16.375 2039.095 16.420 ;
        RECT 2072.370 16.360 2072.690 16.420 ;
      LAYER via ;
        RECT 1709.460 1689.160 1709.720 1689.420 ;
        RECT 1710.840 1689.160 1711.100 1689.420 ;
        RECT 1710.840 18.400 1711.100 18.660 ;
        RECT 2072.400 16.360 2072.660 16.620 ;
      LAYER met2 ;
        RECT 1709.450 1700.000 1709.730 1704.000 ;
        RECT 1709.520 1689.450 1709.660 1700.000 ;
        RECT 1709.460 1689.130 1709.720 1689.450 ;
        RECT 1710.840 1689.130 1711.100 1689.450 ;
        RECT 1710.900 18.690 1711.040 1689.130 ;
        RECT 1710.840 18.370 1711.100 18.690 ;
        RECT 2072.400 16.330 2072.660 16.650 ;
        RECT 2072.460 2.400 2072.600 16.330 ;
=======
      LAYER met1 ;
        RECT 1711.730 1683.920 1712.050 1683.980 ;
        RECT 1716.790 1683.920 1717.110 1683.980 ;
        RECT 1711.730 1683.780 1717.110 1683.920 ;
        RECT 1711.730 1683.720 1712.050 1683.780 ;
        RECT 1716.790 1683.720 1717.110 1683.780 ;
        RECT 1716.790 15.200 1717.110 15.260 ;
        RECT 2072.370 15.200 2072.690 15.260 ;
        RECT 1716.790 15.060 2072.690 15.200 ;
        RECT 1716.790 15.000 1717.110 15.060 ;
        RECT 2072.370 15.000 2072.690 15.060 ;
      LAYER via ;
        RECT 1711.760 1683.720 1712.020 1683.980 ;
        RECT 1716.820 1683.720 1717.080 1683.980 ;
        RECT 1716.820 15.000 1717.080 15.260 ;
        RECT 2072.400 15.000 2072.660 15.260 ;
      LAYER met2 ;
        RECT 1711.750 1700.000 1712.030 1704.000 ;
        RECT 1711.820 1684.010 1711.960 1700.000 ;
        RECT 1711.760 1683.690 1712.020 1684.010 ;
        RECT 1716.820 1683.690 1717.080 1684.010 ;
        RECT 1716.880 15.290 1717.020 1683.690 ;
        RECT 1716.820 14.970 1717.080 15.290 ;
        RECT 2072.400 14.970 2072.660 15.290 ;
        RECT 2072.460 2.400 2072.600 14.970 ;
>>>>>>> re-updated local openlane
        RECT 2072.250 -4.800 2072.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 0.300 ;
=======
      LAYER li1 ;
        RECT 1755.965 1689.545 1756.135 1690.395 ;
        RECT 1779.425 1690.055 1779.595 1690.395 ;
        RECT 1779.425 1689.885 1780.055 1690.055 ;
        RECT 1780.345 1689.885 1780.515 1691.075 ;
        RECT 1828.185 1689.545 1828.355 1691.075 ;
        RECT 1877.405 1689.545 1877.575 1691.075 ;
        RECT 1924.785 1689.545 1924.955 1691.075 ;
        RECT 1925.245 1689.885 1925.875 1690.055 ;
        RECT 1972.625 1689.715 1972.795 1690.055 ;
        RECT 1972.625 1689.545 1973.255 1689.715 ;
      LAYER mcon ;
        RECT 1780.345 1690.905 1780.515 1691.075 ;
        RECT 1755.965 1690.225 1756.135 1690.395 ;
        RECT 1779.425 1690.225 1779.595 1690.395 ;
        RECT 1779.885 1689.885 1780.055 1690.055 ;
        RECT 1828.185 1690.905 1828.355 1691.075 ;
        RECT 1877.405 1690.905 1877.575 1691.075 ;
        RECT 1924.785 1690.905 1924.955 1691.075 ;
        RECT 1925.705 1689.885 1925.875 1690.055 ;
        RECT 1972.625 1689.885 1972.795 1690.055 ;
        RECT 1973.085 1689.545 1973.255 1689.715 ;
      LAYER met1 ;
        RECT 1780.285 1691.060 1780.575 1691.105 ;
        RECT 1828.125 1691.060 1828.415 1691.105 ;
        RECT 1780.285 1690.920 1828.415 1691.060 ;
        RECT 1780.285 1690.875 1780.575 1690.920 ;
        RECT 1828.125 1690.875 1828.415 1690.920 ;
        RECT 1877.345 1691.060 1877.635 1691.105 ;
        RECT 1924.725 1691.060 1925.015 1691.105 ;
        RECT 1877.345 1690.920 1925.015 1691.060 ;
        RECT 1877.345 1690.875 1877.635 1690.920 ;
        RECT 1924.725 1690.875 1925.015 1690.920 ;
        RECT 1755.905 1690.380 1756.195 1690.425 ;
        RECT 1779.365 1690.380 1779.655 1690.425 ;
        RECT 1755.905 1690.240 1779.655 1690.380 ;
        RECT 1755.905 1690.195 1756.195 1690.240 ;
        RECT 1779.365 1690.195 1779.655 1690.240 ;
        RECT 1779.825 1690.040 1780.115 1690.085 ;
        RECT 1780.285 1690.040 1780.575 1690.085 ;
        RECT 1779.825 1689.900 1780.575 1690.040 ;
        RECT 1779.825 1689.855 1780.115 1689.900 ;
        RECT 1780.285 1689.855 1780.575 1689.900 ;
        RECT 1828.570 1689.840 1828.890 1690.100 ;
        RECT 1925.185 1689.855 1925.475 1690.085 ;
        RECT 1925.645 1690.040 1925.935 1690.085 ;
        RECT 1972.565 1690.040 1972.855 1690.085 ;
        RECT 1925.645 1689.900 1972.855 1690.040 ;
        RECT 1925.645 1689.855 1925.935 1689.900 ;
        RECT 1972.565 1689.855 1972.855 1689.900 ;
        RECT 1716.330 1689.700 1716.650 1689.760 ;
        RECT 1755.905 1689.700 1756.195 1689.745 ;
        RECT 1716.330 1689.560 1756.195 1689.700 ;
        RECT 1716.330 1689.500 1716.650 1689.560 ;
        RECT 1755.905 1689.515 1756.195 1689.560 ;
        RECT 1828.125 1689.700 1828.415 1689.745 ;
        RECT 1828.660 1689.700 1828.800 1689.840 ;
        RECT 1828.125 1689.560 1828.800 1689.700 ;
        RECT 1876.410 1689.700 1876.730 1689.760 ;
        RECT 1877.345 1689.700 1877.635 1689.745 ;
        RECT 1876.410 1689.560 1877.635 1689.700 ;
        RECT 1828.125 1689.515 1828.415 1689.560 ;
        RECT 1876.410 1689.500 1876.730 1689.560 ;
        RECT 1877.345 1689.515 1877.635 1689.560 ;
        RECT 1924.725 1689.700 1925.015 1689.745 ;
        RECT 1925.260 1689.700 1925.400 1689.855 ;
        RECT 1924.725 1689.560 1925.400 1689.700 ;
        RECT 1973.025 1689.700 1973.315 1689.745 ;
        RECT 2083.870 1689.700 2084.190 1689.760 ;
        RECT 1973.025 1689.560 2084.190 1689.700 ;
        RECT 1924.725 1689.515 1925.015 1689.560 ;
        RECT 1973.025 1689.515 1973.315 1689.560 ;
        RECT 2083.870 1689.500 2084.190 1689.560 ;
        RECT 2083.870 35.940 2084.190 36.000 ;
        RECT 2089.850 35.940 2090.170 36.000 ;
        RECT 2083.870 35.800 2090.170 35.940 ;
        RECT 2083.870 35.740 2084.190 35.800 ;
        RECT 2089.850 35.740 2090.170 35.800 ;
      LAYER via ;
        RECT 1828.600 1689.840 1828.860 1690.100 ;
        RECT 1716.360 1689.500 1716.620 1689.760 ;
        RECT 1876.440 1689.500 1876.700 1689.760 ;
        RECT 2083.900 1689.500 2084.160 1689.760 ;
        RECT 2083.900 35.740 2084.160 36.000 ;
        RECT 2089.880 35.740 2090.140 36.000 ;
      LAYER met2 ;
        RECT 1716.350 1700.000 1716.630 1704.000 ;
        RECT 1716.420 1689.790 1716.560 1700.000 ;
        RECT 1828.590 1689.955 1828.870 1690.325 ;
        RECT 1876.430 1689.955 1876.710 1690.325 ;
        RECT 1828.600 1689.810 1828.860 1689.955 ;
        RECT 1876.500 1689.790 1876.640 1689.955 ;
        RECT 1716.360 1689.470 1716.620 1689.790 ;
        RECT 1876.440 1689.470 1876.700 1689.790 ;
        RECT 2083.900 1689.470 2084.160 1689.790 ;
        RECT 2083.960 36.030 2084.100 1689.470 ;
        RECT 2083.900 35.710 2084.160 36.030 ;
        RECT 2089.880 35.710 2090.140 36.030 ;
        RECT 2089.940 2.400 2090.080 35.710 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 1828.590 1690.000 1828.870 1690.280 ;
        RECT 1876.430 1690.000 1876.710 1690.280 ;
      LAYER met3 ;
        RECT 1828.565 1690.290 1828.895 1690.305 ;
        RECT 1876.405 1690.290 1876.735 1690.305 ;
        RECT 1828.565 1689.990 1876.735 1690.290 ;
        RECT 1828.565 1689.975 1828.895 1689.990 ;
        RECT 1876.405 1689.975 1876.735 1689.990 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 0.300 ;
=======
      LAYER li1 ;
        RECT 1965.725 16.405 1965.895 20.655 ;
      LAYER mcon ;
        RECT 1965.725 20.485 1965.895 20.655 ;
      LAYER met1 ;
        RECT 1719.090 1686.300 1719.410 1686.360 ;
        RECT 1924.710 1686.300 1925.030 1686.360 ;
        RECT 1942.190 1686.300 1942.510 1686.360 ;
        RECT 1719.090 1686.160 1897.800 1686.300 ;
        RECT 1719.090 1686.100 1719.410 1686.160 ;
        RECT 1897.660 1685.960 1897.800 1686.160 ;
        RECT 1924.710 1686.160 1942.510 1686.300 ;
        RECT 1924.710 1686.100 1925.030 1686.160 ;
        RECT 1942.190 1686.100 1942.510 1686.160 ;
        RECT 1898.490 1685.960 1898.810 1686.020 ;
        RECT 1897.660 1685.820 1898.810 1685.960 ;
        RECT 1898.490 1685.760 1898.810 1685.820 ;
        RECT 1965.665 20.640 1965.955 20.685 ;
        RECT 2107.790 20.640 2108.110 20.700 ;
        RECT 1965.665 20.500 2108.110 20.640 ;
        RECT 1965.665 20.455 1965.955 20.500 ;
        RECT 2107.790 20.440 2108.110 20.500 ;
        RECT 1942.190 16.560 1942.510 16.620 ;
        RECT 1965.665 16.560 1965.955 16.605 ;
        RECT 1942.190 16.420 1965.955 16.560 ;
        RECT 1942.190 16.360 1942.510 16.420 ;
        RECT 1965.665 16.375 1965.955 16.420 ;
      LAYER via ;
        RECT 1719.120 1686.100 1719.380 1686.360 ;
        RECT 1924.740 1686.100 1925.000 1686.360 ;
        RECT 1942.220 1686.100 1942.480 1686.360 ;
        RECT 1898.520 1685.760 1898.780 1686.020 ;
        RECT 2107.820 20.440 2108.080 20.700 ;
        RECT 1942.220 16.360 1942.480 16.620 ;
      LAYER met2 ;
        RECT 1719.110 1700.000 1719.390 1704.000 ;
        RECT 1719.180 1686.390 1719.320 1700.000 ;
        RECT 1719.120 1686.070 1719.380 1686.390 ;
        RECT 1924.740 1686.245 1925.000 1686.390 ;
        RECT 1898.510 1685.875 1898.790 1686.245 ;
        RECT 1924.730 1685.875 1925.010 1686.245 ;
        RECT 1942.220 1686.070 1942.480 1686.390 ;
        RECT 1898.520 1685.730 1898.780 1685.875 ;
        RECT 1942.280 16.650 1942.420 1686.070 ;
        RECT 2107.820 20.410 2108.080 20.730 ;
        RECT 1942.220 16.330 1942.480 16.650 ;
        RECT 2107.880 2.400 2108.020 20.410 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
      LAYER via2 ;
        RECT 1898.510 1685.920 1898.790 1686.200 ;
        RECT 1924.730 1685.920 1925.010 1686.200 ;
      LAYER met3 ;
        RECT 1898.485 1686.210 1898.815 1686.225 ;
        RECT 1924.705 1686.210 1925.035 1686.225 ;
        RECT 1898.485 1685.910 1925.035 1686.210 ;
        RECT 1898.485 1685.895 1898.815 1685.910 ;
        RECT 1924.705 1685.895 1925.035 1685.910 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1721.390 1684.940 1721.710 1685.000 ;
        RECT 1724.610 1684.940 1724.930 1685.000 ;
        RECT 1721.390 1684.800 1724.930 1684.940 ;
        RECT 1721.390 1684.740 1721.710 1684.800 ;
        RECT 1724.610 1684.740 1724.930 1684.800 ;
        RECT 1724.610 15.540 1724.930 15.600 ;
        RECT 1724.610 15.400 2073.060 15.540 ;
        RECT 1724.610 15.340 1724.930 15.400 ;
        RECT 2072.920 15.200 2073.060 15.400 ;
        RECT 2107.790 15.200 2108.110 15.260 ;
        RECT 2072.920 15.060 2108.110 15.200 ;
        RECT 2107.790 15.000 2108.110 15.060 ;
      LAYER via ;
        RECT 1721.420 1684.740 1721.680 1685.000 ;
        RECT 1724.640 1684.740 1724.900 1685.000 ;
        RECT 1724.640 15.340 1724.900 15.600 ;
        RECT 2107.820 15.000 2108.080 15.260 ;
      LAYER met2 ;
        RECT 1721.410 1700.000 1721.690 1704.000 ;
        RECT 1721.480 1685.030 1721.620 1700.000 ;
        RECT 1721.420 1684.710 1721.680 1685.030 ;
        RECT 1724.640 1684.710 1724.900 1685.030 ;
        RECT 1724.700 15.630 1724.840 1684.710 ;
        RECT 1724.640 15.310 1724.900 15.630 ;
        RECT 2107.820 14.970 2108.080 15.290 ;
        RECT 2107.880 2.400 2108.020 14.970 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1723.690 1689.700 1724.010 1689.760 ;
        RECT 2066.390 1689.700 2066.710 1689.760 ;
        RECT 1723.690 1689.560 2066.710 1689.700 ;
        RECT 1723.690 1689.500 1724.010 1689.560 ;
        RECT 2066.390 1689.500 2066.710 1689.560 ;
        RECT 2066.390 19.620 2066.710 19.680 ;
        RECT 2125.730 19.620 2126.050 19.680 ;
        RECT 2066.390 19.480 2126.050 19.620 ;
        RECT 2066.390 19.420 2066.710 19.480 ;
        RECT 2125.730 19.420 2126.050 19.480 ;
      LAYER via ;
        RECT 1723.720 1689.500 1723.980 1689.760 ;
        RECT 2066.420 1689.500 2066.680 1689.760 ;
        RECT 2066.420 19.420 2066.680 19.680 ;
        RECT 2125.760 19.420 2126.020 19.680 ;
      LAYER met2 ;
        RECT 1723.710 1700.000 1723.990 1704.000 ;
        RECT 1723.780 1689.790 1723.920 1700.000 ;
        RECT 1723.720 1689.470 1723.980 1689.790 ;
        RECT 2066.420 1689.470 2066.680 1689.790 ;
        RECT 2066.480 19.710 2066.620 1689.470 ;
        RECT 2066.420 19.390 2066.680 19.710 ;
        RECT 2125.760 19.390 2126.020 19.710 ;
        RECT 2125.820 2.400 2125.960 19.390 ;
=======
      LAYER li1 ;
        RECT 1828.645 1689.205 1829.735 1689.375 ;
        RECT 1876.945 1689.205 1878.035 1689.375 ;
        RECT 1925.245 1689.205 1926.335 1689.375 ;
        RECT 2125.345 48.365 2125.515 96.475 ;
      LAYER mcon ;
        RECT 1829.565 1689.205 1829.735 1689.375 ;
        RECT 1877.865 1689.205 1878.035 1689.375 ;
        RECT 1926.165 1689.205 1926.335 1689.375 ;
        RECT 2125.345 96.305 2125.515 96.475 ;
      LAYER met1 ;
        RECT 1725.990 1690.040 1726.310 1690.100 ;
        RECT 1725.990 1689.900 1777.280 1690.040 ;
        RECT 1725.990 1689.840 1726.310 1689.900 ;
        RECT 1777.140 1689.360 1777.280 1689.900 ;
        RECT 1828.585 1689.360 1828.875 1689.405 ;
        RECT 1777.140 1689.220 1828.875 1689.360 ;
        RECT 1828.585 1689.175 1828.875 1689.220 ;
        RECT 1829.505 1689.360 1829.795 1689.405 ;
        RECT 1876.885 1689.360 1877.175 1689.405 ;
        RECT 1829.505 1689.220 1877.175 1689.360 ;
        RECT 1829.505 1689.175 1829.795 1689.220 ;
        RECT 1876.885 1689.175 1877.175 1689.220 ;
        RECT 1877.805 1689.360 1878.095 1689.405 ;
        RECT 1925.185 1689.360 1925.475 1689.405 ;
        RECT 1877.805 1689.220 1925.475 1689.360 ;
        RECT 1877.805 1689.175 1878.095 1689.220 ;
        RECT 1925.185 1689.175 1925.475 1689.220 ;
        RECT 1926.105 1689.360 1926.395 1689.405 ;
        RECT 2125.270 1689.360 2125.590 1689.420 ;
        RECT 1926.105 1689.220 2125.590 1689.360 ;
        RECT 1926.105 1689.175 1926.395 1689.220 ;
        RECT 2125.270 1689.160 2125.590 1689.220 ;
        RECT 2125.270 96.460 2125.590 96.520 ;
        RECT 2125.270 96.320 2125.785 96.460 ;
        RECT 2125.270 96.260 2125.590 96.320 ;
        RECT 2125.285 48.520 2125.575 48.565 ;
        RECT 2125.730 48.520 2126.050 48.580 ;
        RECT 2125.285 48.380 2126.050 48.520 ;
        RECT 2125.285 48.335 2125.575 48.380 ;
        RECT 2125.730 48.320 2126.050 48.380 ;
      LAYER via ;
        RECT 1726.020 1689.840 1726.280 1690.100 ;
        RECT 2125.300 1689.160 2125.560 1689.420 ;
        RECT 2125.300 96.260 2125.560 96.520 ;
        RECT 2125.760 48.320 2126.020 48.580 ;
      LAYER met2 ;
        RECT 1726.010 1700.000 1726.290 1704.000 ;
        RECT 1726.080 1690.130 1726.220 1700.000 ;
        RECT 1726.020 1689.810 1726.280 1690.130 ;
        RECT 2125.300 1689.130 2125.560 1689.450 ;
        RECT 2125.360 96.550 2125.500 1689.130 ;
        RECT 2125.300 96.230 2125.560 96.550 ;
        RECT 2125.760 48.290 2126.020 48.610 ;
        RECT 2125.820 2.400 2125.960 48.290 ;
>>>>>>> re-updated local openlane
        RECT 2125.610 -4.800 2126.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1731.510 15.880 1731.830 15.940 ;
        RECT 2143.670 15.880 2143.990 15.940 ;
        RECT 1731.510 15.740 2143.990 15.880 ;
        RECT 1731.510 15.680 1731.830 15.740 ;
        RECT 2143.670 15.680 2143.990 15.740 ;
      LAYER via ;
        RECT 1731.540 15.680 1731.800 15.940 ;
        RECT 2143.700 15.680 2143.960 15.940 ;
      LAYER met2 ;
        RECT 1731.070 1700.410 1731.350 1704.000 ;
        RECT 1731.070 1700.270 1731.740 1700.410 ;
        RECT 1731.070 1700.000 1731.350 1700.270 ;
        RECT 1731.600 15.970 1731.740 1700.270 ;
        RECT 1731.540 15.650 1731.800 15.970 ;
        RECT 2143.700 15.650 2143.960 15.970 ;
        RECT 2143.760 2.400 2143.900 15.650 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 0.300 ;
=======
      LAYER li1 ;
        RECT 1771.605 1689.205 1772.695 1689.375 ;
        RECT 1771.605 1687.845 1771.775 1689.205 ;
      LAYER mcon ;
        RECT 1772.525 1689.205 1772.695 1689.375 ;
      LAYER met1 ;
        RECT 2159.770 1689.500 2160.090 1689.760 ;
        RECT 1772.465 1689.360 1772.755 1689.405 ;
        RECT 2159.860 1689.360 2160.000 1689.500 ;
        RECT 1772.465 1689.220 2160.000 1689.360 ;
        RECT 1772.465 1689.175 1772.755 1689.220 ;
        RECT 1733.350 1688.000 1733.670 1688.060 ;
        RECT 1771.545 1688.000 1771.835 1688.045 ;
        RECT 1733.350 1687.860 1771.835 1688.000 ;
        RECT 1733.350 1687.800 1733.670 1687.860 ;
        RECT 1771.545 1687.815 1771.835 1687.860 ;
      LAYER via ;
        RECT 2159.800 1689.500 2160.060 1689.760 ;
        RECT 1733.380 1687.800 1733.640 1688.060 ;
      LAYER met2 ;
        RECT 1733.370 1700.000 1733.650 1704.000 ;
        RECT 1733.440 1688.090 1733.580 1700.000 ;
        RECT 2159.800 1689.470 2160.060 1689.790 ;
        RECT 1733.380 1687.770 1733.640 1688.090 ;
        RECT 2159.860 17.410 2160.000 1689.470 ;
        RECT 2159.860 17.270 2161.840 17.410 ;
        RECT 2161.700 2.400 2161.840 17.270 ;
=======
      LAYER met1 ;
        RECT 1735.650 1689.360 1735.970 1689.420 ;
        RECT 1735.650 1689.220 1757.960 1689.360 ;
        RECT 1735.650 1689.160 1735.970 1689.220 ;
        RECT 1757.820 1689.020 1757.960 1689.220 ;
        RECT 2159.770 1689.020 2160.090 1689.080 ;
        RECT 1757.820 1688.880 2160.090 1689.020 ;
        RECT 2159.770 1688.820 2160.090 1688.880 ;
        RECT 2159.310 48.520 2159.630 48.580 ;
        RECT 2161.610 48.520 2161.930 48.580 ;
        RECT 2159.310 48.380 2161.930 48.520 ;
        RECT 2159.310 48.320 2159.630 48.380 ;
        RECT 2161.610 48.320 2161.930 48.380 ;
      LAYER via ;
        RECT 1735.680 1689.160 1735.940 1689.420 ;
        RECT 2159.800 1688.820 2160.060 1689.080 ;
        RECT 2159.340 48.320 2159.600 48.580 ;
        RECT 2161.640 48.320 2161.900 48.580 ;
      LAYER met2 ;
        RECT 1735.670 1700.000 1735.950 1704.000 ;
        RECT 1735.740 1689.450 1735.880 1700.000 ;
        RECT 1735.680 1689.130 1735.940 1689.450 ;
        RECT 2159.800 1688.790 2160.060 1689.110 ;
        RECT 2159.860 73.170 2160.000 1688.790 ;
        RECT 2159.400 73.030 2160.000 73.170 ;
        RECT 2159.400 48.610 2159.540 73.030 ;
        RECT 2159.340 48.290 2159.600 48.610 ;
        RECT 2161.640 48.290 2161.900 48.610 ;
        RECT 2161.700 2.400 2161.840 48.290 ;
>>>>>>> re-updated local openlane
        RECT 2161.490 -4.800 2162.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 0.300 ;
=======
      LAYER li1 ;
        RECT 2111.545 18.445 2111.715 20.655 ;
      LAYER mcon ;
        RECT 2111.545 20.485 2111.715 20.655 ;
      LAYER met1 ;
        RECT 1738.410 1690.040 1738.730 1690.100 ;
        RECT 2080.190 1690.040 2080.510 1690.100 ;
        RECT 1738.410 1689.900 2080.510 1690.040 ;
        RECT 1738.410 1689.840 1738.730 1689.900 ;
        RECT 2080.190 1689.840 2080.510 1689.900 ;
        RECT 2111.485 20.640 2111.775 20.685 ;
        RECT 2121.130 20.640 2121.450 20.700 ;
        RECT 2111.485 20.500 2121.450 20.640 ;
        RECT 2111.485 20.455 2111.775 20.500 ;
        RECT 2121.130 20.440 2121.450 20.500 ;
        RECT 2091.230 18.600 2091.550 18.660 ;
        RECT 2111.485 18.600 2111.775 18.645 ;
        RECT 2091.230 18.460 2111.775 18.600 ;
        RECT 2091.230 18.400 2091.550 18.460 ;
        RECT 2111.485 18.415 2111.775 18.460 ;
        RECT 2159.310 18.600 2159.630 18.660 ;
        RECT 2179.090 18.600 2179.410 18.660 ;
        RECT 2159.310 18.460 2179.410 18.600 ;
        RECT 2159.310 18.400 2159.630 18.460 ;
        RECT 2179.090 18.400 2179.410 18.460 ;
      LAYER via ;
        RECT 1738.440 1689.840 1738.700 1690.100 ;
        RECT 2080.220 1689.840 2080.480 1690.100 ;
        RECT 2121.160 20.440 2121.420 20.700 ;
        RECT 2091.260 18.400 2091.520 18.660 ;
        RECT 2159.340 18.400 2159.600 18.660 ;
        RECT 2179.120 18.400 2179.380 18.660 ;
      LAYER met2 ;
        RECT 1738.430 1700.000 1738.710 1704.000 ;
        RECT 1738.500 1690.130 1738.640 1700.000 ;
        RECT 1738.440 1689.810 1738.700 1690.130 ;
        RECT 2080.220 1689.810 2080.480 1690.130 ;
        RECT 2080.280 20.925 2080.420 1689.810 ;
        RECT 2080.210 20.555 2080.490 20.925 ;
        RECT 2091.250 20.555 2091.530 20.925 ;
        RECT 2121.150 20.555 2121.430 20.925 ;
        RECT 2159.330 20.555 2159.610 20.925 ;
        RECT 2091.320 18.690 2091.460 20.555 ;
        RECT 2121.160 20.410 2121.420 20.555 ;
        RECT 2159.400 18.690 2159.540 20.555 ;
        RECT 2091.260 18.370 2091.520 18.690 ;
        RECT 2159.340 18.370 2159.600 18.690 ;
        RECT 2179.120 18.370 2179.380 18.690 ;
        RECT 2179.180 2.400 2179.320 18.370 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
      LAYER via2 ;
        RECT 2080.210 20.600 2080.490 20.880 ;
        RECT 2091.250 20.600 2091.530 20.880 ;
        RECT 2121.150 20.600 2121.430 20.880 ;
        RECT 2159.330 20.600 2159.610 20.880 ;
      LAYER met3 ;
        RECT 2080.185 20.890 2080.515 20.905 ;
        RECT 2091.225 20.890 2091.555 20.905 ;
        RECT 2080.185 20.590 2091.555 20.890 ;
        RECT 2080.185 20.575 2080.515 20.590 ;
        RECT 2091.225 20.575 2091.555 20.590 ;
        RECT 2121.125 20.890 2121.455 20.905 ;
        RECT 2159.305 20.890 2159.635 20.905 ;
        RECT 2121.125 20.590 2159.635 20.890 ;
        RECT 2121.125 20.575 2121.455 20.590 ;
        RECT 2159.305 20.575 2159.635 20.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1740.710 1684.940 1741.030 1685.000 ;
        RECT 1745.310 1684.940 1745.630 1685.000 ;
        RECT 1740.710 1684.800 1745.630 1684.940 ;
        RECT 1740.710 1684.740 1741.030 1684.800 ;
        RECT 1745.310 1684.740 1745.630 1684.800 ;
        RECT 1744.850 16.560 1745.170 16.620 ;
        RECT 1744.850 16.420 1746.000 16.560 ;
        RECT 1744.850 16.360 1745.170 16.420 ;
        RECT 1745.860 16.220 1746.000 16.420 ;
        RECT 2179.090 16.220 2179.410 16.280 ;
        RECT 1745.860 16.080 2179.410 16.220 ;
        RECT 2179.090 16.020 2179.410 16.080 ;
      LAYER via ;
        RECT 1740.740 1684.740 1741.000 1685.000 ;
        RECT 1745.340 1684.740 1745.600 1685.000 ;
        RECT 1744.880 16.360 1745.140 16.620 ;
        RECT 2179.120 16.020 2179.380 16.280 ;
      LAYER met2 ;
        RECT 1740.730 1700.000 1741.010 1704.000 ;
        RECT 1740.800 1685.030 1740.940 1700.000 ;
        RECT 1740.740 1684.710 1741.000 1685.030 ;
        RECT 1745.340 1684.710 1745.600 1685.030 ;
        RECT 1745.400 28.290 1745.540 1684.710 ;
        RECT 1744.940 28.150 1745.540 28.290 ;
        RECT 1744.940 16.650 1745.080 28.150 ;
        RECT 1744.880 16.330 1745.140 16.650 ;
        RECT 2179.120 15.990 2179.380 16.310 ;
        RECT 2179.180 2.400 2179.320 15.990 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 0.300 ;
=======
      LAYER li1 ;
        RECT 1800.585 1687.505 1800.755 1688.695 ;
        RECT 2194.345 1587.205 2194.515 1594.175 ;
        RECT 2194.345 766.105 2194.515 814.215 ;
        RECT 2194.345 669.545 2194.515 717.655 ;
        RECT 2194.345 572.645 2194.515 620.755 ;
        RECT 2194.345 476.085 2194.515 524.195 ;
        RECT 2194.345 379.525 2194.515 427.635 ;
        RECT 2194.345 282.965 2194.515 331.075 ;
        RECT 2194.345 186.405 2194.515 234.515 ;
        RECT 2194.345 61.285 2194.515 137.955 ;
      LAYER mcon ;
        RECT 1800.585 1688.525 1800.755 1688.695 ;
        RECT 2194.345 1594.005 2194.515 1594.175 ;
        RECT 2194.345 814.045 2194.515 814.215 ;
        RECT 2194.345 717.485 2194.515 717.655 ;
        RECT 2194.345 620.585 2194.515 620.755 ;
        RECT 2194.345 524.025 2194.515 524.195 ;
        RECT 2194.345 427.465 2194.515 427.635 ;
        RECT 2194.345 330.905 2194.515 331.075 ;
        RECT 2194.345 234.345 2194.515 234.515 ;
        RECT 2194.345 137.785 2194.515 137.955 ;
      LAYER met1 ;
        RECT 1745.310 1689.020 1745.630 1689.080 ;
        RECT 1745.310 1688.880 1752.900 1689.020 ;
        RECT 1745.310 1688.820 1745.630 1688.880 ;
        RECT 1752.760 1687.660 1752.900 1688.880 ;
        RECT 1800.525 1688.680 1800.815 1688.725 ;
        RECT 2194.270 1688.680 2194.590 1688.740 ;
        RECT 1800.525 1688.540 2194.590 1688.680 ;
        RECT 1800.525 1688.495 1800.815 1688.540 ;
        RECT 2194.270 1688.480 2194.590 1688.540 ;
        RECT 1800.525 1687.660 1800.815 1687.705 ;
        RECT 1752.760 1687.520 1800.815 1687.660 ;
        RECT 1800.525 1687.475 1800.815 1687.520 ;
        RECT 2194.270 1594.160 2194.590 1594.220 ;
        RECT 2194.075 1594.020 2194.590 1594.160 ;
        RECT 2194.270 1593.960 2194.590 1594.020 ;
        RECT 2194.270 1587.360 2194.590 1587.420 ;
        RECT 2194.075 1587.220 2194.590 1587.360 ;
        RECT 2194.270 1587.160 2194.590 1587.220 ;
        RECT 2194.270 1208.060 2194.590 1208.320 ;
        RECT 2194.360 1207.640 2194.500 1208.060 ;
        RECT 2194.270 1207.380 2194.590 1207.640 ;
        RECT 2194.270 1152.500 2194.590 1152.560 ;
        RECT 2195.190 1152.500 2195.510 1152.560 ;
        RECT 2194.270 1152.360 2195.510 1152.500 ;
        RECT 2194.270 1152.300 2194.590 1152.360 ;
        RECT 2195.190 1152.300 2195.510 1152.360 ;
        RECT 2194.270 1007.320 2194.590 1007.380 ;
        RECT 2195.190 1007.320 2195.510 1007.380 ;
        RECT 2194.270 1007.180 2195.510 1007.320 ;
        RECT 2194.270 1007.120 2194.590 1007.180 ;
        RECT 2195.190 1007.120 2195.510 1007.180 ;
        RECT 2194.270 910.760 2194.590 910.820 ;
        RECT 2194.730 910.760 2195.050 910.820 ;
        RECT 2194.270 910.620 2195.050 910.760 ;
        RECT 2194.270 910.560 2194.590 910.620 ;
        RECT 2194.730 910.560 2195.050 910.620 ;
        RECT 2194.270 814.200 2194.590 814.260 ;
        RECT 2194.075 814.060 2194.590 814.200 ;
        RECT 2194.270 814.000 2194.590 814.060 ;
        RECT 2194.270 766.260 2194.590 766.320 ;
        RECT 2194.075 766.120 2194.590 766.260 ;
        RECT 2194.270 766.060 2194.590 766.120 ;
        RECT 2194.270 717.640 2194.590 717.700 ;
        RECT 2194.075 717.500 2194.590 717.640 ;
        RECT 2194.270 717.440 2194.590 717.500 ;
        RECT 2194.270 669.700 2194.590 669.760 ;
        RECT 2194.075 669.560 2194.590 669.700 ;
        RECT 2194.270 669.500 2194.590 669.560 ;
        RECT 2194.270 620.740 2194.590 620.800 ;
        RECT 2194.075 620.600 2194.590 620.740 ;
        RECT 2194.270 620.540 2194.590 620.600 ;
        RECT 2194.270 572.800 2194.590 572.860 ;
        RECT 2194.075 572.660 2194.590 572.800 ;
        RECT 2194.270 572.600 2194.590 572.660 ;
        RECT 2194.270 524.180 2194.590 524.240 ;
        RECT 2194.075 524.040 2194.590 524.180 ;
        RECT 2194.270 523.980 2194.590 524.040 ;
        RECT 2194.270 476.240 2194.590 476.300 ;
        RECT 2194.075 476.100 2194.590 476.240 ;
        RECT 2194.270 476.040 2194.590 476.100 ;
        RECT 2194.270 427.620 2194.590 427.680 ;
        RECT 2194.075 427.480 2194.590 427.620 ;
        RECT 2194.270 427.420 2194.590 427.480 ;
        RECT 2194.270 379.680 2194.590 379.740 ;
        RECT 2194.075 379.540 2194.590 379.680 ;
        RECT 2194.270 379.480 2194.590 379.540 ;
        RECT 2194.270 331.060 2194.590 331.120 ;
        RECT 2194.075 330.920 2194.590 331.060 ;
        RECT 2194.270 330.860 2194.590 330.920 ;
        RECT 2194.270 283.120 2194.590 283.180 ;
        RECT 2194.075 282.980 2194.590 283.120 ;
        RECT 2194.270 282.920 2194.590 282.980 ;
        RECT 2194.270 234.500 2194.590 234.560 ;
        RECT 2194.075 234.360 2194.590 234.500 ;
        RECT 2194.270 234.300 2194.590 234.360 ;
        RECT 2194.270 186.560 2194.590 186.620 ;
        RECT 2194.075 186.420 2194.590 186.560 ;
        RECT 2194.270 186.360 2194.590 186.420 ;
        RECT 2194.270 137.940 2194.590 138.000 ;
        RECT 2194.075 137.800 2194.590 137.940 ;
        RECT 2194.270 137.740 2194.590 137.800 ;
        RECT 2194.285 61.440 2194.575 61.485 ;
        RECT 2197.030 61.440 2197.350 61.500 ;
        RECT 2194.285 61.300 2197.350 61.440 ;
        RECT 2194.285 61.255 2194.575 61.300 ;
        RECT 2197.030 61.240 2197.350 61.300 ;
      LAYER via ;
        RECT 1745.340 1688.820 1745.600 1689.080 ;
        RECT 2194.300 1688.480 2194.560 1688.740 ;
        RECT 2194.300 1593.960 2194.560 1594.220 ;
        RECT 2194.300 1587.160 2194.560 1587.420 ;
        RECT 2194.300 1208.060 2194.560 1208.320 ;
        RECT 2194.300 1207.380 2194.560 1207.640 ;
        RECT 2194.300 1152.300 2194.560 1152.560 ;
        RECT 2195.220 1152.300 2195.480 1152.560 ;
        RECT 2194.300 1007.120 2194.560 1007.380 ;
        RECT 2195.220 1007.120 2195.480 1007.380 ;
        RECT 2194.300 910.560 2194.560 910.820 ;
        RECT 2194.760 910.560 2195.020 910.820 ;
        RECT 2194.300 814.000 2194.560 814.260 ;
        RECT 2194.300 766.060 2194.560 766.320 ;
        RECT 2194.300 717.440 2194.560 717.700 ;
        RECT 2194.300 669.500 2194.560 669.760 ;
        RECT 2194.300 620.540 2194.560 620.800 ;
        RECT 2194.300 572.600 2194.560 572.860 ;
        RECT 2194.300 523.980 2194.560 524.240 ;
        RECT 2194.300 476.040 2194.560 476.300 ;
        RECT 2194.300 427.420 2194.560 427.680 ;
        RECT 2194.300 379.480 2194.560 379.740 ;
        RECT 2194.300 330.860 2194.560 331.120 ;
        RECT 2194.300 282.920 2194.560 283.180 ;
        RECT 2194.300 234.300 2194.560 234.560 ;
        RECT 2194.300 186.360 2194.560 186.620 ;
        RECT 2194.300 137.740 2194.560 138.000 ;
        RECT 2197.060 61.240 2197.320 61.500 ;
      LAYER met2 ;
        RECT 1745.330 1700.000 1745.610 1704.000 ;
        RECT 1745.400 1689.110 1745.540 1700.000 ;
        RECT 1745.340 1688.790 1745.600 1689.110 ;
        RECT 2194.300 1688.450 2194.560 1688.770 ;
        RECT 2194.360 1594.250 2194.500 1688.450 ;
        RECT 2194.300 1593.930 2194.560 1594.250 ;
        RECT 2194.300 1587.130 2194.560 1587.450 ;
        RECT 2194.360 1208.350 2194.500 1587.130 ;
        RECT 2194.300 1208.030 2194.560 1208.350 ;
        RECT 2194.300 1207.350 2194.560 1207.670 ;
        RECT 2194.360 1200.725 2194.500 1207.350 ;
        RECT 2194.290 1200.355 2194.570 1200.725 ;
        RECT 2195.210 1200.355 2195.490 1200.725 ;
        RECT 2195.280 1152.590 2195.420 1200.355 ;
        RECT 2194.300 1152.270 2194.560 1152.590 ;
        RECT 2195.220 1152.270 2195.480 1152.590 ;
        RECT 2194.360 1104.165 2194.500 1152.270 ;
        RECT 2194.290 1103.795 2194.570 1104.165 ;
        RECT 2195.210 1103.795 2195.490 1104.165 ;
        RECT 2195.280 1055.885 2195.420 1103.795 ;
        RECT 2194.290 1055.515 2194.570 1055.885 ;
        RECT 2195.210 1055.515 2195.490 1055.885 ;
        RECT 2194.360 1007.410 2194.500 1055.515 ;
        RECT 2194.300 1007.090 2194.560 1007.410 ;
        RECT 2195.220 1007.090 2195.480 1007.410 ;
        RECT 2195.280 959.325 2195.420 1007.090 ;
        RECT 2194.290 958.955 2194.570 959.325 ;
        RECT 2195.210 958.955 2195.490 959.325 ;
        RECT 2194.360 910.850 2194.500 958.955 ;
        RECT 2194.300 910.530 2194.560 910.850 ;
        RECT 2194.760 910.530 2195.020 910.850 ;
        RECT 2194.820 821.170 2194.960 910.530 ;
        RECT 2194.360 821.030 2194.960 821.170 ;
        RECT 2194.360 814.290 2194.500 821.030 ;
        RECT 2194.300 813.970 2194.560 814.290 ;
        RECT 2194.300 766.030 2194.560 766.350 ;
        RECT 2194.360 717.730 2194.500 766.030 ;
        RECT 2194.300 717.410 2194.560 717.730 ;
        RECT 2194.300 669.470 2194.560 669.790 ;
        RECT 2194.360 620.830 2194.500 669.470 ;
        RECT 2194.300 620.510 2194.560 620.830 ;
        RECT 2194.300 572.570 2194.560 572.890 ;
        RECT 2194.360 524.270 2194.500 572.570 ;
        RECT 2194.300 523.950 2194.560 524.270 ;
        RECT 2194.300 476.010 2194.560 476.330 ;
        RECT 2194.360 427.710 2194.500 476.010 ;
        RECT 2194.300 427.390 2194.560 427.710 ;
        RECT 2194.300 379.450 2194.560 379.770 ;
        RECT 2194.360 331.150 2194.500 379.450 ;
        RECT 2194.300 330.830 2194.560 331.150 ;
        RECT 2194.300 282.890 2194.560 283.210 ;
        RECT 2194.360 234.590 2194.500 282.890 ;
        RECT 2194.300 234.270 2194.560 234.590 ;
        RECT 2194.300 186.330 2194.560 186.650 ;
        RECT 2194.360 138.030 2194.500 186.330 ;
        RECT 2194.300 137.710 2194.560 138.030 ;
        RECT 2197.060 61.210 2197.320 61.530 ;
        RECT 2197.120 2.400 2197.260 61.210 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 2194.290 1200.400 2194.570 1200.680 ;
        RECT 2195.210 1200.400 2195.490 1200.680 ;
        RECT 2194.290 1103.840 2194.570 1104.120 ;
        RECT 2195.210 1103.840 2195.490 1104.120 ;
        RECT 2194.290 1055.560 2194.570 1055.840 ;
        RECT 2195.210 1055.560 2195.490 1055.840 ;
        RECT 2194.290 959.000 2194.570 959.280 ;
        RECT 2195.210 959.000 2195.490 959.280 ;
      LAYER met3 ;
        RECT 2194.265 1200.690 2194.595 1200.705 ;
        RECT 2195.185 1200.690 2195.515 1200.705 ;
        RECT 2194.265 1200.390 2195.515 1200.690 ;
        RECT 2194.265 1200.375 2194.595 1200.390 ;
        RECT 2195.185 1200.375 2195.515 1200.390 ;
        RECT 2194.265 1104.130 2194.595 1104.145 ;
        RECT 2195.185 1104.130 2195.515 1104.145 ;
        RECT 2194.265 1103.830 2195.515 1104.130 ;
        RECT 2194.265 1103.815 2194.595 1103.830 ;
        RECT 2195.185 1103.815 2195.515 1103.830 ;
        RECT 2194.265 1055.850 2194.595 1055.865 ;
        RECT 2195.185 1055.850 2195.515 1055.865 ;
        RECT 2194.265 1055.550 2195.515 1055.850 ;
        RECT 2194.265 1055.535 2194.595 1055.550 ;
        RECT 2195.185 1055.535 2195.515 1055.550 ;
        RECT 2194.265 959.290 2194.595 959.305 ;
        RECT 2195.185 959.290 2195.515 959.305 ;
        RECT 2194.265 958.990 2195.515 959.290 ;
        RECT 2194.265 958.975 2194.595 958.990 ;
        RECT 2195.185 958.975 2195.515 958.990 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 0.300 ;
=======
      LAYER met1 ;
        RECT 1750.370 1683.920 1750.690 1683.980 ;
        RECT 1752.210 1683.920 1752.530 1683.980 ;
        RECT 1750.370 1683.780 1752.530 1683.920 ;
        RECT 1750.370 1683.720 1750.690 1683.780 ;
        RECT 1752.210 1683.720 1752.530 1683.780 ;
        RECT 1752.210 16.560 1752.530 16.620 ;
        RECT 2214.970 16.560 2215.290 16.620 ;
        RECT 1752.210 16.420 2215.290 16.560 ;
        RECT 1752.210 16.360 1752.530 16.420 ;
        RECT 2214.970 16.360 2215.290 16.420 ;
      LAYER via ;
        RECT 1750.400 1683.720 1750.660 1683.980 ;
        RECT 1752.240 1683.720 1752.500 1683.980 ;
        RECT 1752.240 16.360 1752.500 16.620 ;
        RECT 2215.000 16.360 2215.260 16.620 ;
      LAYER met2 ;
        RECT 1750.390 1700.000 1750.670 1704.000 ;
        RECT 1750.460 1684.010 1750.600 1700.000 ;
        RECT 1750.400 1683.690 1750.660 1684.010 ;
        RECT 1752.240 1683.690 1752.500 1684.010 ;
        RECT 1752.300 16.650 1752.440 1683.690 ;
        RECT 1752.240 16.330 1752.500 16.650 ;
        RECT 2215.000 16.330 2215.260 16.650 ;
        RECT 2215.060 2.400 2215.200 16.330 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1752.670 1689.020 1752.990 1689.080 ;
        RECT 1752.670 1688.880 1766.240 1689.020 ;
        RECT 1752.670 1688.820 1752.990 1688.880 ;
        RECT 1766.100 1688.680 1766.240 1688.880 ;
        RECT 2228.770 1688.680 2229.090 1688.740 ;
        RECT 1766.100 1688.540 2229.090 1688.680 ;
        RECT 2228.770 1688.480 2229.090 1688.540 ;
      LAYER via ;
        RECT 1752.700 1688.820 1752.960 1689.080 ;
        RECT 2228.800 1688.480 2229.060 1688.740 ;
      LAYER met2 ;
        RECT 1752.690 1700.000 1752.970 1704.000 ;
        RECT 1752.760 1689.110 1752.900 1700.000 ;
        RECT 1752.700 1688.790 1752.960 1689.110 ;
        RECT 2228.800 1688.450 2229.060 1688.770 ;
        RECT 2228.860 17.410 2229.000 1688.450 ;
        RECT 2228.860 17.270 2233.140 17.410 ;
        RECT 2233.000 2.400 2233.140 17.270 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 2230.225 1317.245 2230.395 1393.575 ;
        RECT 2230.225 1220.685 2230.395 1297.015 ;
        RECT 2228.845 1110.865 2229.015 1124.975 ;
        RECT 2229.305 1027.565 2229.475 1038.615 ;
        RECT 2229.765 979.285 2229.935 1007.335 ;
        RECT 2229.765 786.505 2229.935 821.015 ;
        RECT 2229.765 572.645 2229.935 620.755 ;
        RECT 2229.765 350.965 2229.935 386.155 ;
        RECT 2232.065 48.365 2232.235 124.015 ;
      LAYER mcon ;
        RECT 2230.225 1393.405 2230.395 1393.575 ;
        RECT 2230.225 1296.845 2230.395 1297.015 ;
        RECT 2228.845 1124.805 2229.015 1124.975 ;
        RECT 2229.305 1038.445 2229.475 1038.615 ;
        RECT 2229.765 1007.165 2229.935 1007.335 ;
        RECT 2229.765 820.845 2229.935 821.015 ;
        RECT 2229.765 620.585 2229.935 620.755 ;
        RECT 2229.765 385.985 2229.935 386.155 ;
        RECT 2232.065 123.845 2232.235 124.015 ;
      LAYER met1 ;
        RECT 1754.970 1688.340 1755.290 1688.400 ;
        RECT 2228.770 1688.340 2229.090 1688.400 ;
        RECT 1754.970 1688.200 2229.090 1688.340 ;
        RECT 1754.970 1688.140 1755.290 1688.200 ;
        RECT 2228.770 1688.140 2229.090 1688.200 ;
        RECT 2228.770 1684.940 2229.090 1685.000 ;
        RECT 2230.150 1684.940 2230.470 1685.000 ;
        RECT 2228.770 1684.800 2230.470 1684.940 ;
        RECT 2228.770 1684.740 2229.090 1684.800 ;
        RECT 2230.150 1684.740 2230.470 1684.800 ;
        RECT 2229.690 1594.160 2230.010 1594.220 ;
        RECT 2230.150 1594.160 2230.470 1594.220 ;
        RECT 2229.690 1594.020 2230.470 1594.160 ;
        RECT 2229.690 1593.960 2230.010 1594.020 ;
        RECT 2230.150 1593.960 2230.470 1594.020 ;
        RECT 2229.690 1559.820 2230.010 1559.880 ;
        RECT 2230.150 1559.820 2230.470 1559.880 ;
        RECT 2229.690 1559.680 2230.470 1559.820 ;
        RECT 2229.690 1559.620 2230.010 1559.680 ;
        RECT 2230.150 1559.620 2230.470 1559.680 ;
        RECT 2229.230 1511.200 2229.550 1511.260 ;
        RECT 2230.150 1511.200 2230.470 1511.260 ;
        RECT 2229.230 1511.060 2230.470 1511.200 ;
        RECT 2229.230 1511.000 2229.550 1511.060 ;
        RECT 2230.150 1511.000 2230.470 1511.060 ;
        RECT 2228.310 1448.980 2228.630 1449.040 ;
        RECT 2230.150 1448.980 2230.470 1449.040 ;
        RECT 2228.310 1448.840 2230.470 1448.980 ;
        RECT 2228.310 1448.780 2228.630 1448.840 ;
        RECT 2230.150 1448.780 2230.470 1448.840 ;
        RECT 2229.690 1393.560 2230.010 1393.620 ;
        RECT 2230.165 1393.560 2230.455 1393.605 ;
        RECT 2229.690 1393.420 2230.455 1393.560 ;
        RECT 2229.690 1393.360 2230.010 1393.420 ;
        RECT 2230.165 1393.375 2230.455 1393.420 ;
        RECT 2230.150 1317.400 2230.470 1317.460 ;
        RECT 2229.955 1317.260 2230.470 1317.400 ;
        RECT 2230.150 1317.200 2230.470 1317.260 ;
        RECT 2230.150 1297.000 2230.470 1297.060 ;
        RECT 2229.955 1296.860 2230.470 1297.000 ;
        RECT 2230.150 1296.800 2230.470 1296.860 ;
        RECT 2230.150 1220.840 2230.470 1220.900 ;
        RECT 2229.955 1220.700 2230.470 1220.840 ;
        RECT 2230.150 1220.640 2230.470 1220.700 ;
        RECT 2229.230 1173.240 2229.550 1173.300 ;
        RECT 2230.150 1173.240 2230.470 1173.300 ;
        RECT 2229.230 1173.100 2230.470 1173.240 ;
        RECT 2229.230 1173.040 2229.550 1173.100 ;
        RECT 2230.150 1173.040 2230.470 1173.100 ;
        RECT 2228.770 1124.960 2229.090 1125.020 ;
        RECT 2228.575 1124.820 2229.090 1124.960 ;
        RECT 2228.770 1124.760 2229.090 1124.820 ;
        RECT 2228.770 1111.020 2229.090 1111.080 ;
        RECT 2228.575 1110.880 2229.090 1111.020 ;
        RECT 2228.770 1110.820 2229.090 1110.880 ;
        RECT 2228.770 1076.480 2229.090 1076.740 ;
        RECT 2228.860 1076.000 2229.000 1076.480 ;
        RECT 2229.230 1076.000 2229.550 1076.060 ;
        RECT 2228.860 1075.860 2229.550 1076.000 ;
        RECT 2229.230 1075.800 2229.550 1075.860 ;
        RECT 2229.230 1038.600 2229.550 1038.660 ;
        RECT 2229.035 1038.460 2229.550 1038.600 ;
        RECT 2229.230 1038.400 2229.550 1038.460 ;
        RECT 2229.245 1027.720 2229.535 1027.765 ;
        RECT 2230.150 1027.720 2230.470 1027.780 ;
        RECT 2229.245 1027.580 2230.470 1027.720 ;
        RECT 2229.245 1027.535 2229.535 1027.580 ;
        RECT 2230.150 1027.520 2230.470 1027.580 ;
        RECT 2229.705 1007.320 2229.995 1007.365 ;
        RECT 2230.150 1007.320 2230.470 1007.380 ;
        RECT 2229.705 1007.180 2230.470 1007.320 ;
        RECT 2229.705 1007.135 2229.995 1007.180 ;
        RECT 2230.150 1007.120 2230.470 1007.180 ;
        RECT 2229.690 979.440 2230.010 979.500 ;
        RECT 2229.495 979.300 2230.010 979.440 ;
        RECT 2229.690 979.240 2230.010 979.300 ;
        RECT 2229.690 917.900 2230.010 917.960 ;
        RECT 2231.070 917.900 2231.390 917.960 ;
        RECT 2229.690 917.760 2231.390 917.900 ;
        RECT 2229.690 917.700 2230.010 917.760 ;
        RECT 2231.070 917.700 2231.390 917.760 ;
        RECT 2230.150 869.620 2230.470 869.680 ;
        RECT 2231.070 869.620 2231.390 869.680 ;
        RECT 2230.150 869.480 2231.390 869.620 ;
        RECT 2230.150 869.420 2230.470 869.480 ;
        RECT 2231.070 869.420 2231.390 869.480 ;
        RECT 2229.230 835.280 2229.550 835.340 ;
        RECT 2230.150 835.280 2230.470 835.340 ;
        RECT 2229.230 835.140 2230.470 835.280 ;
        RECT 2229.230 835.080 2229.550 835.140 ;
        RECT 2230.150 835.080 2230.470 835.140 ;
        RECT 2229.690 821.000 2230.010 821.060 ;
        RECT 2229.495 820.860 2230.010 821.000 ;
        RECT 2229.690 820.800 2230.010 820.860 ;
        RECT 2229.690 786.660 2230.010 786.720 ;
        RECT 2229.495 786.520 2230.010 786.660 ;
        RECT 2229.690 786.460 2230.010 786.520 ;
        RECT 2229.230 738.380 2229.550 738.440 ;
        RECT 2230.150 738.380 2230.470 738.440 ;
        RECT 2229.230 738.240 2230.470 738.380 ;
        RECT 2229.230 738.180 2229.550 738.240 ;
        RECT 2230.150 738.180 2230.470 738.240 ;
        RECT 2230.150 690.100 2230.470 690.160 ;
        RECT 2229.780 689.960 2230.470 690.100 ;
        RECT 2229.780 689.820 2229.920 689.960 ;
        RECT 2230.150 689.900 2230.470 689.960 ;
        RECT 2229.690 689.560 2230.010 689.820 ;
        RECT 2229.690 641.620 2230.010 641.880 ;
        RECT 2229.780 641.480 2229.920 641.620 ;
        RECT 2230.150 641.480 2230.470 641.540 ;
        RECT 2229.780 641.340 2230.470 641.480 ;
        RECT 2230.150 641.280 2230.470 641.340 ;
        RECT 2229.705 620.740 2229.995 620.785 ;
        RECT 2230.150 620.740 2230.470 620.800 ;
        RECT 2229.705 620.600 2230.470 620.740 ;
        RECT 2229.705 620.555 2229.995 620.600 ;
        RECT 2230.150 620.540 2230.470 620.600 ;
        RECT 2229.690 572.800 2230.010 572.860 ;
        RECT 2229.495 572.660 2230.010 572.800 ;
        RECT 2229.690 572.600 2230.010 572.660 ;
        RECT 2229.690 545.600 2230.010 545.660 ;
        RECT 2229.320 545.460 2230.010 545.600 ;
        RECT 2229.320 544.980 2229.460 545.460 ;
        RECT 2229.690 545.400 2230.010 545.460 ;
        RECT 2229.230 544.720 2229.550 544.980 ;
        RECT 2229.230 496.780 2229.550 497.040 ;
        RECT 2229.320 496.640 2229.460 496.780 ;
        RECT 2230.150 496.640 2230.470 496.700 ;
        RECT 2229.320 496.500 2230.470 496.640 ;
        RECT 2230.150 496.440 2230.470 496.500 ;
        RECT 2229.230 448.700 2229.550 448.760 ;
        RECT 2230.150 448.700 2230.470 448.760 ;
        RECT 2229.230 448.560 2230.470 448.700 ;
        RECT 2229.230 448.500 2229.550 448.560 ;
        RECT 2230.150 448.500 2230.470 448.560 ;
        RECT 2229.690 386.140 2230.010 386.200 ;
        RECT 2229.495 386.000 2230.010 386.140 ;
        RECT 2229.690 385.940 2230.010 386.000 ;
        RECT 2229.690 351.120 2230.010 351.180 ;
        RECT 2229.495 350.980 2230.010 351.120 ;
        RECT 2229.690 350.920 2230.010 350.980 ;
        RECT 2229.690 303.860 2230.010 303.920 ;
        RECT 2229.690 303.720 2230.380 303.860 ;
        RECT 2229.690 303.660 2230.010 303.720 ;
        RECT 2230.240 303.240 2230.380 303.720 ;
        RECT 2230.150 302.980 2230.470 303.240 ;
        RECT 2229.230 159.020 2229.550 159.080 ;
        RECT 2229.230 158.880 2229.920 159.020 ;
        RECT 2229.230 158.820 2229.550 158.880 ;
        RECT 2229.780 158.740 2229.920 158.880 ;
        RECT 2229.690 158.480 2230.010 158.740 ;
        RECT 2229.230 124.000 2229.550 124.060 ;
        RECT 2232.005 124.000 2232.295 124.045 ;
        RECT 2229.230 123.860 2232.295 124.000 ;
        RECT 2229.230 123.800 2229.550 123.860 ;
        RECT 2232.005 123.815 2232.295 123.860 ;
        RECT 2232.005 48.520 2232.295 48.565 ;
        RECT 2232.910 48.520 2233.230 48.580 ;
        RECT 2232.005 48.380 2233.230 48.520 ;
        RECT 2232.005 48.335 2232.295 48.380 ;
        RECT 2232.910 48.320 2233.230 48.380 ;
        RECT 2232.910 2.960 2233.230 3.020 ;
        RECT 2233.370 2.960 2233.690 3.020 ;
        RECT 2232.910 2.820 2233.690 2.960 ;
        RECT 2232.910 2.760 2233.230 2.820 ;
        RECT 2233.370 2.760 2233.690 2.820 ;
      LAYER via ;
        RECT 1755.000 1688.140 1755.260 1688.400 ;
        RECT 2228.800 1688.140 2229.060 1688.400 ;
        RECT 2228.800 1684.740 2229.060 1685.000 ;
        RECT 2230.180 1684.740 2230.440 1685.000 ;
        RECT 2229.720 1593.960 2229.980 1594.220 ;
        RECT 2230.180 1593.960 2230.440 1594.220 ;
        RECT 2229.720 1559.620 2229.980 1559.880 ;
        RECT 2230.180 1559.620 2230.440 1559.880 ;
        RECT 2229.260 1511.000 2229.520 1511.260 ;
        RECT 2230.180 1511.000 2230.440 1511.260 ;
        RECT 2228.340 1448.780 2228.600 1449.040 ;
        RECT 2230.180 1448.780 2230.440 1449.040 ;
        RECT 2229.720 1393.360 2229.980 1393.620 ;
        RECT 2230.180 1317.200 2230.440 1317.460 ;
        RECT 2230.180 1296.800 2230.440 1297.060 ;
        RECT 2230.180 1220.640 2230.440 1220.900 ;
        RECT 2229.260 1173.040 2229.520 1173.300 ;
        RECT 2230.180 1173.040 2230.440 1173.300 ;
        RECT 2228.800 1124.760 2229.060 1125.020 ;
        RECT 2228.800 1110.820 2229.060 1111.080 ;
        RECT 2228.800 1076.480 2229.060 1076.740 ;
        RECT 2229.260 1075.800 2229.520 1076.060 ;
        RECT 2229.260 1038.400 2229.520 1038.660 ;
        RECT 2230.180 1027.520 2230.440 1027.780 ;
        RECT 2230.180 1007.120 2230.440 1007.380 ;
        RECT 2229.720 979.240 2229.980 979.500 ;
        RECT 2229.720 917.700 2229.980 917.960 ;
        RECT 2231.100 917.700 2231.360 917.960 ;
        RECT 2230.180 869.420 2230.440 869.680 ;
        RECT 2231.100 869.420 2231.360 869.680 ;
        RECT 2229.260 835.080 2229.520 835.340 ;
        RECT 2230.180 835.080 2230.440 835.340 ;
        RECT 2229.720 820.800 2229.980 821.060 ;
        RECT 2229.720 786.460 2229.980 786.720 ;
        RECT 2229.260 738.180 2229.520 738.440 ;
        RECT 2230.180 738.180 2230.440 738.440 ;
        RECT 2230.180 689.900 2230.440 690.160 ;
        RECT 2229.720 689.560 2229.980 689.820 ;
        RECT 2229.720 641.620 2229.980 641.880 ;
        RECT 2230.180 641.280 2230.440 641.540 ;
        RECT 2230.180 620.540 2230.440 620.800 ;
        RECT 2229.720 572.600 2229.980 572.860 ;
        RECT 2229.720 545.400 2229.980 545.660 ;
        RECT 2229.260 544.720 2229.520 544.980 ;
        RECT 2229.260 496.780 2229.520 497.040 ;
        RECT 2230.180 496.440 2230.440 496.700 ;
        RECT 2229.260 448.500 2229.520 448.760 ;
        RECT 2230.180 448.500 2230.440 448.760 ;
        RECT 2229.720 385.940 2229.980 386.200 ;
        RECT 2229.720 350.920 2229.980 351.180 ;
        RECT 2229.720 303.660 2229.980 303.920 ;
        RECT 2230.180 302.980 2230.440 303.240 ;
        RECT 2229.260 158.820 2229.520 159.080 ;
        RECT 2229.720 158.480 2229.980 158.740 ;
        RECT 2229.260 123.800 2229.520 124.060 ;
        RECT 2232.940 48.320 2233.200 48.580 ;
        RECT 2232.940 2.760 2233.200 3.020 ;
        RECT 2233.400 2.760 2233.660 3.020 ;
      LAYER met2 ;
        RECT 1754.990 1700.000 1755.270 1704.000 ;
        RECT 1755.060 1688.430 1755.200 1700.000 ;
        RECT 1755.000 1688.110 1755.260 1688.430 ;
        RECT 2228.800 1688.110 2229.060 1688.430 ;
        RECT 2228.860 1685.030 2229.000 1688.110 ;
        RECT 2228.800 1684.710 2229.060 1685.030 ;
        RECT 2230.180 1684.710 2230.440 1685.030 ;
        RECT 2230.240 1594.250 2230.380 1684.710 ;
        RECT 2229.720 1593.930 2229.980 1594.250 ;
        RECT 2230.180 1593.930 2230.440 1594.250 ;
        RECT 2229.780 1559.910 2229.920 1593.930 ;
        RECT 2229.720 1559.590 2229.980 1559.910 ;
        RECT 2230.180 1559.590 2230.440 1559.910 ;
        RECT 2230.240 1511.290 2230.380 1559.590 ;
        RECT 2229.260 1510.970 2229.520 1511.290 ;
        RECT 2230.180 1510.970 2230.440 1511.290 ;
        RECT 2229.320 1510.690 2229.460 1510.970 ;
        RECT 2229.320 1510.550 2229.920 1510.690 ;
        RECT 2229.780 1463.090 2229.920 1510.550 ;
        RECT 2229.780 1462.950 2230.380 1463.090 ;
        RECT 2230.240 1449.070 2230.380 1462.950 ;
        RECT 2228.340 1448.750 2228.600 1449.070 ;
        RECT 2230.180 1448.750 2230.440 1449.070 ;
        RECT 2228.400 1401.325 2228.540 1448.750 ;
        RECT 2228.330 1400.955 2228.610 1401.325 ;
        RECT 2229.250 1401.210 2229.530 1401.325 ;
        RECT 2229.250 1401.070 2229.920 1401.210 ;
        RECT 2229.250 1400.955 2229.530 1401.070 ;
        RECT 2229.780 1393.650 2229.920 1401.070 ;
        RECT 2229.720 1393.330 2229.980 1393.650 ;
        RECT 2230.180 1317.170 2230.440 1317.490 ;
        RECT 2230.240 1297.090 2230.380 1317.170 ;
        RECT 2230.180 1296.770 2230.440 1297.090 ;
        RECT 2230.180 1220.610 2230.440 1220.930 ;
        RECT 2230.240 1173.330 2230.380 1220.610 ;
        RECT 2229.260 1173.010 2229.520 1173.330 ;
        RECT 2230.180 1173.010 2230.440 1173.330 ;
        RECT 2229.320 1159.130 2229.460 1173.010 ;
        RECT 2228.860 1158.990 2229.460 1159.130 ;
        RECT 2228.860 1125.050 2229.000 1158.990 ;
        RECT 2228.800 1124.730 2229.060 1125.050 ;
        RECT 2228.800 1110.790 2229.060 1111.110 ;
        RECT 2228.860 1076.770 2229.000 1110.790 ;
        RECT 2228.800 1076.450 2229.060 1076.770 ;
        RECT 2229.260 1075.770 2229.520 1076.090 ;
        RECT 2229.320 1038.690 2229.460 1075.770 ;
        RECT 2229.260 1038.370 2229.520 1038.690 ;
        RECT 2230.180 1027.490 2230.440 1027.810 ;
        RECT 2230.240 1007.410 2230.380 1027.490 ;
        RECT 2230.180 1007.090 2230.440 1007.410 ;
        RECT 2229.720 979.210 2229.980 979.530 ;
        RECT 2229.780 917.990 2229.920 979.210 ;
        RECT 2229.720 917.670 2229.980 917.990 ;
        RECT 2231.100 917.670 2231.360 917.990 ;
        RECT 2231.160 869.710 2231.300 917.670 ;
        RECT 2230.180 869.390 2230.440 869.710 ;
        RECT 2231.100 869.390 2231.360 869.710 ;
        RECT 2230.240 835.370 2230.380 869.390 ;
        RECT 2229.260 835.050 2229.520 835.370 ;
        RECT 2230.180 835.050 2230.440 835.370 ;
        RECT 2229.320 834.770 2229.460 835.050 ;
        RECT 2229.320 834.630 2229.920 834.770 ;
        RECT 2229.780 821.090 2229.920 834.630 ;
        RECT 2229.720 820.770 2229.980 821.090 ;
        RECT 2229.720 786.430 2229.980 786.750 ;
        RECT 2229.780 772.890 2229.920 786.430 ;
        RECT 2229.780 772.750 2230.380 772.890 ;
        RECT 2230.240 738.470 2230.380 772.750 ;
        RECT 2229.260 738.210 2229.520 738.470 ;
        RECT 2230.180 738.210 2230.440 738.470 ;
        RECT 2229.260 738.150 2230.440 738.210 ;
        RECT 2229.320 738.070 2230.380 738.150 ;
        RECT 2230.240 690.190 2230.380 738.070 ;
        RECT 2230.180 689.870 2230.440 690.190 ;
        RECT 2229.720 689.530 2229.980 689.850 ;
        RECT 2229.780 641.910 2229.920 689.530 ;
        RECT 2229.720 641.590 2229.980 641.910 ;
        RECT 2230.180 641.250 2230.440 641.570 ;
        RECT 2230.240 620.830 2230.380 641.250 ;
        RECT 2230.180 620.510 2230.440 620.830 ;
        RECT 2229.720 572.570 2229.980 572.890 ;
        RECT 2229.780 545.690 2229.920 572.570 ;
        RECT 2229.720 545.370 2229.980 545.690 ;
        RECT 2229.260 544.690 2229.520 545.010 ;
        RECT 2229.320 497.070 2229.460 544.690 ;
        RECT 2229.260 496.750 2229.520 497.070 ;
        RECT 2230.180 496.410 2230.440 496.730 ;
        RECT 2230.240 448.790 2230.380 496.410 ;
        RECT 2229.260 448.530 2229.520 448.790 ;
        RECT 2230.180 448.530 2230.440 448.790 ;
        RECT 2229.260 448.470 2230.440 448.530 ;
        RECT 2229.320 448.390 2230.380 448.470 ;
        RECT 2230.240 401.045 2230.380 448.390 ;
        RECT 2230.170 400.675 2230.450 401.045 ;
        RECT 2229.710 386.395 2229.990 386.765 ;
        RECT 2229.780 386.230 2229.920 386.395 ;
        RECT 2229.720 385.910 2229.980 386.230 ;
        RECT 2229.720 350.890 2229.980 351.210 ;
        RECT 2229.780 303.950 2229.920 350.890 ;
        RECT 2229.720 303.630 2229.980 303.950 ;
        RECT 2230.180 302.950 2230.440 303.270 ;
        RECT 2230.240 255.410 2230.380 302.950 ;
        RECT 2229.320 255.270 2230.380 255.410 ;
        RECT 2229.320 159.110 2229.460 255.270 ;
        RECT 2229.260 158.790 2229.520 159.110 ;
        RECT 2229.720 158.450 2229.980 158.770 ;
        RECT 2229.780 131.650 2229.920 158.450 ;
        RECT 2229.320 131.510 2229.920 131.650 ;
        RECT 2229.320 124.090 2229.460 131.510 ;
        RECT 2229.260 123.770 2229.520 124.090 ;
        RECT 2232.940 48.290 2233.200 48.610 ;
        RECT 2233.000 48.010 2233.140 48.290 ;
        RECT 2233.000 47.870 2233.600 48.010 ;
        RECT 2233.460 3.050 2233.600 47.870 ;
        RECT 2232.940 2.730 2233.200 3.050 ;
        RECT 2233.400 2.730 2233.660 3.050 ;
        RECT 2233.000 2.400 2233.140 2.730 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
      LAYER via2 ;
        RECT 2228.330 1401.000 2228.610 1401.280 ;
        RECT 2229.250 1401.000 2229.530 1401.280 ;
        RECT 2230.170 400.720 2230.450 401.000 ;
        RECT 2229.710 386.440 2229.990 386.720 ;
      LAYER met3 ;
        RECT 2228.305 1401.290 2228.635 1401.305 ;
        RECT 2229.225 1401.290 2229.555 1401.305 ;
        RECT 2228.305 1400.990 2229.555 1401.290 ;
        RECT 2228.305 1400.975 2228.635 1400.990 ;
        RECT 2229.225 1400.975 2229.555 1400.990 ;
        RECT 2229.430 401.010 2229.810 401.020 ;
        RECT 2230.145 401.010 2230.475 401.025 ;
        RECT 2229.430 400.710 2230.475 401.010 ;
        RECT 2229.430 400.700 2229.810 400.710 ;
        RECT 2230.145 400.695 2230.475 400.710 ;
        RECT 2229.685 386.740 2230.015 386.745 ;
        RECT 2229.430 386.730 2230.015 386.740 ;
        RECT 2229.430 386.430 2230.240 386.730 ;
        RECT 2229.430 386.420 2230.015 386.430 ;
        RECT 2229.685 386.415 2230.015 386.420 ;
      LAYER via3 ;
        RECT 2229.460 400.700 2229.780 401.020 ;
        RECT 2229.460 386.420 2229.780 386.740 ;
      LAYER met4 ;
        RECT 2229.455 400.695 2229.785 401.025 ;
        RECT 2229.470 386.745 2229.770 400.695 ;
        RECT 2229.455 386.415 2229.785 386.745 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 0.300 ;
=======
      LAYER met1 ;
        RECT 787.590 44.440 787.910 44.500 ;
        RECT 1360.290 44.440 1360.610 44.500 ;
        RECT 787.590 44.300 1360.610 44.440 ;
        RECT 787.590 44.240 787.910 44.300 ;
        RECT 1360.290 44.240 1360.610 44.300 ;
      LAYER via ;
        RECT 787.620 44.240 787.880 44.500 ;
        RECT 1360.320 44.240 1360.580 44.500 ;
      LAYER met2 ;
        RECT 1362.150 1700.410 1362.430 1704.000 ;
        RECT 1361.300 1700.270 1362.430 1700.410 ;
        RECT 1361.300 1677.970 1361.440 1700.270 ;
        RECT 1362.150 1700.000 1362.430 1700.270 ;
        RECT 1360.380 1677.830 1361.440 1677.970 ;
        RECT 1360.380 44.530 1360.520 1677.830 ;
        RECT 787.620 44.210 787.880 44.530 ;
        RECT 1360.320 44.210 1360.580 44.530 ;
        RECT 787.680 2.400 787.820 44.210 ;
=======
      LAYER li1 ;
        RECT 1361.285 1587.205 1361.455 1635.315 ;
      LAYER mcon ;
        RECT 1361.285 1635.145 1361.455 1635.315 ;
      LAYER met1 ;
        RECT 1361.225 1635.300 1361.515 1635.345 ;
        RECT 1362.130 1635.300 1362.450 1635.360 ;
        RECT 1361.225 1635.160 1362.450 1635.300 ;
        RECT 1361.225 1635.115 1361.515 1635.160 ;
        RECT 1362.130 1635.100 1362.450 1635.160 ;
        RECT 1361.210 1587.360 1361.530 1587.420 ;
        RECT 1361.015 1587.220 1361.530 1587.360 ;
        RECT 1361.210 1587.160 1361.530 1587.220 ;
        RECT 1360.750 96.800 1361.070 96.860 ;
        RECT 1361.210 96.800 1361.530 96.860 ;
        RECT 1360.750 96.660 1361.530 96.800 ;
        RECT 1360.750 96.600 1361.070 96.660 ;
        RECT 1361.210 96.600 1361.530 96.660 ;
        RECT 787.590 43.420 787.910 43.480 ;
        RECT 1360.750 43.420 1361.070 43.480 ;
        RECT 787.590 43.280 1361.070 43.420 ;
        RECT 787.590 43.220 787.910 43.280 ;
        RECT 1360.750 43.220 1361.070 43.280 ;
      LAYER via ;
        RECT 1362.160 1635.100 1362.420 1635.360 ;
        RECT 1361.240 1587.160 1361.500 1587.420 ;
        RECT 1360.780 96.600 1361.040 96.860 ;
        RECT 1361.240 96.600 1361.500 96.860 ;
        RECT 787.620 43.220 787.880 43.480 ;
        RECT 1360.780 43.220 1361.040 43.480 ;
      LAYER met2 ;
        RECT 1363.070 1700.410 1363.350 1704.000 ;
        RECT 1362.220 1700.270 1363.350 1700.410 ;
        RECT 1362.220 1635.390 1362.360 1700.270 ;
        RECT 1363.070 1700.000 1363.350 1700.270 ;
        RECT 1362.160 1635.070 1362.420 1635.390 ;
        RECT 1361.240 1587.130 1361.500 1587.450 ;
        RECT 1361.300 1583.450 1361.440 1587.130 ;
        RECT 1360.840 1583.310 1361.440 1583.450 ;
        RECT 1360.840 1558.970 1360.980 1583.310 ;
        RECT 1360.840 1558.830 1361.440 1558.970 ;
        RECT 1361.300 1125.130 1361.440 1558.830 ;
        RECT 1360.840 1124.990 1361.440 1125.130 ;
        RECT 1360.840 1124.450 1360.980 1124.990 ;
        RECT 1360.840 1124.310 1361.440 1124.450 ;
        RECT 1361.300 932.010 1361.440 1124.310 ;
        RECT 1360.840 931.870 1361.440 932.010 ;
        RECT 1360.840 931.330 1360.980 931.870 ;
        RECT 1360.840 931.190 1361.440 931.330 ;
        RECT 1361.300 835.450 1361.440 931.190 ;
        RECT 1360.840 835.310 1361.440 835.450 ;
        RECT 1360.840 834.770 1360.980 835.310 ;
        RECT 1360.840 834.630 1361.440 834.770 ;
        RECT 1361.300 642.330 1361.440 834.630 ;
        RECT 1360.840 642.190 1361.440 642.330 ;
        RECT 1360.840 641.650 1360.980 642.190 ;
        RECT 1360.840 641.510 1361.440 641.650 ;
        RECT 1361.300 96.890 1361.440 641.510 ;
        RECT 1360.780 96.570 1361.040 96.890 ;
        RECT 1361.240 96.570 1361.500 96.890 ;
        RECT 1360.840 43.510 1360.980 96.570 ;
        RECT 787.620 43.190 787.880 43.510 ;
        RECT 1360.780 43.190 1361.040 43.510 ;
        RECT 787.680 2.400 787.820 43.190 ;
>>>>>>> re-updated local openlane
        RECT 787.470 -4.800 788.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 0.300 ;
=======
      LAYER met1 ;
        RECT 1760.030 1684.600 1760.350 1684.660 ;
        RECT 1766.010 1684.600 1766.330 1684.660 ;
        RECT 1760.030 1684.460 1766.330 1684.600 ;
        RECT 1760.030 1684.400 1760.350 1684.460 ;
        RECT 1766.010 1684.400 1766.330 1684.460 ;
        RECT 1766.010 16.900 1766.330 16.960 ;
        RECT 2250.850 16.900 2251.170 16.960 ;
        RECT 1766.010 16.760 2251.170 16.900 ;
        RECT 1766.010 16.700 1766.330 16.760 ;
        RECT 2250.850 16.700 2251.170 16.760 ;
      LAYER via ;
        RECT 1760.060 1684.400 1760.320 1684.660 ;
        RECT 1766.040 1684.400 1766.300 1684.660 ;
        RECT 1766.040 16.700 1766.300 16.960 ;
        RECT 2250.880 16.700 2251.140 16.960 ;
      LAYER met2 ;
        RECT 1760.050 1700.000 1760.330 1704.000 ;
        RECT 1760.120 1684.690 1760.260 1700.000 ;
        RECT 1760.060 1684.370 1760.320 1684.690 ;
        RECT 1766.040 1684.370 1766.300 1684.690 ;
        RECT 1766.100 16.990 1766.240 1684.370 ;
        RECT 1766.040 16.670 1766.300 16.990 ;
        RECT 2250.880 16.670 2251.140 16.990 ;
        RECT 2250.940 2.400 2251.080 16.670 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 0.300 ;
=======
      LAYER met1 ;
        RECT 1764.630 1688.000 1764.950 1688.060 ;
        RECT 2263.270 1688.000 2263.590 1688.060 ;
        RECT 1764.630 1687.860 2263.590 1688.000 ;
        RECT 1764.630 1687.800 1764.950 1687.860 ;
        RECT 2263.270 1687.800 2263.590 1687.860 ;
        RECT 2263.270 62.120 2263.590 62.180 ;
        RECT 2268.330 62.120 2268.650 62.180 ;
        RECT 2263.270 61.980 2268.650 62.120 ;
        RECT 2263.270 61.920 2263.590 61.980 ;
        RECT 2268.330 61.920 2268.650 61.980 ;
      LAYER via ;
        RECT 1764.660 1687.800 1764.920 1688.060 ;
        RECT 2263.300 1687.800 2263.560 1688.060 ;
        RECT 2263.300 61.920 2263.560 62.180 ;
        RECT 2268.360 61.920 2268.620 62.180 ;
      LAYER met2 ;
        RECT 1764.650 1700.000 1764.930 1704.000 ;
        RECT 1764.720 1688.090 1764.860 1700.000 ;
        RECT 1764.660 1687.770 1764.920 1688.090 ;
        RECT 2263.300 1687.770 2263.560 1688.090 ;
        RECT 2263.360 62.210 2263.500 1687.770 ;
        RECT 2263.300 61.890 2263.560 62.210 ;
        RECT 2268.360 61.890 2268.620 62.210 ;
        RECT 2268.420 2.400 2268.560 61.890 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 0.300 ;
=======
      LAYER met1 ;
        RECT 1771.070 20.640 1771.390 20.700 ;
        RECT 2286.270 20.640 2286.590 20.700 ;
        RECT 1771.070 20.500 2286.590 20.640 ;
        RECT 1771.070 20.440 1771.390 20.500 ;
        RECT 2286.270 20.440 2286.590 20.500 ;
      LAYER via ;
        RECT 1771.100 20.440 1771.360 20.700 ;
        RECT 2286.300 20.440 2286.560 20.700 ;
      LAYER met2 ;
        RECT 1769.710 1700.410 1769.990 1704.000 ;
        RECT 1769.710 1700.270 1770.380 1700.410 ;
        RECT 1769.710 1700.000 1769.990 1700.270 ;
        RECT 1770.240 1656.210 1770.380 1700.270 ;
        RECT 1770.240 1656.070 1771.300 1656.210 ;
        RECT 1771.160 20.730 1771.300 1656.070 ;
        RECT 1771.100 20.410 1771.360 20.730 ;
        RECT 2286.300 20.410 2286.560 20.730 ;
        RECT 2286.360 2.400 2286.500 20.410 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 0.300 ;
=======
      LAYER met1 ;
        RECT 1772.450 1688.000 1772.770 1688.060 ;
        RECT 2266.490 1688.000 2266.810 1688.060 ;
        RECT 1772.450 1687.860 2266.810 1688.000 ;
        RECT 1772.450 1687.800 1772.770 1687.860 ;
        RECT 2266.490 1687.800 2266.810 1687.860 ;
        RECT 2268.880 14.040 2300.300 14.180 ;
        RECT 2266.490 13.840 2266.810 13.900 ;
        RECT 2268.880 13.840 2269.020 14.040 ;
        RECT 2266.490 13.700 2269.020 13.840 ;
        RECT 2266.490 13.640 2266.810 13.700 ;
        RECT 2300.160 13.500 2300.300 14.040 ;
        RECT 2304.210 13.500 2304.530 13.560 ;
        RECT 2300.160 13.360 2304.530 13.500 ;
        RECT 2304.210 13.300 2304.530 13.360 ;
      LAYER via ;
        RECT 1772.480 1687.800 1772.740 1688.060 ;
        RECT 2266.520 1687.800 2266.780 1688.060 ;
        RECT 2266.520 13.640 2266.780 13.900 ;
        RECT 2304.240 13.300 2304.500 13.560 ;
      LAYER met2 ;
        RECT 1772.010 1700.410 1772.290 1704.000 ;
        RECT 1772.010 1700.270 1772.680 1700.410 ;
        RECT 1772.010 1700.000 1772.290 1700.270 ;
        RECT 1772.540 1688.090 1772.680 1700.270 ;
        RECT 1772.480 1687.770 1772.740 1688.090 ;
        RECT 2266.520 1687.770 2266.780 1688.090 ;
        RECT 2266.580 13.930 2266.720 1687.770 ;
        RECT 2266.520 13.610 2266.780 13.930 ;
        RECT 2304.240 13.270 2304.500 13.590 ;
        RECT 2304.300 2.400 2304.440 13.270 ;
=======
      LAYER li1 ;
        RECT 1779.885 1690.565 1780.055 1695.495 ;
        RECT 1824.965 1687.505 1825.135 1690.395 ;
      LAYER mcon ;
        RECT 1779.885 1695.325 1780.055 1695.495 ;
        RECT 1824.965 1690.225 1825.135 1690.395 ;
      LAYER met1 ;
        RECT 1774.290 1695.480 1774.610 1695.540 ;
        RECT 1779.825 1695.480 1780.115 1695.525 ;
        RECT 1774.290 1695.340 1780.115 1695.480 ;
        RECT 1774.290 1695.280 1774.610 1695.340 ;
        RECT 1779.825 1695.295 1780.115 1695.340 ;
        RECT 1779.825 1690.535 1780.115 1690.765 ;
        RECT 1779.900 1690.380 1780.040 1690.535 ;
        RECT 1824.905 1690.380 1825.195 1690.425 ;
        RECT 1779.900 1690.240 1825.195 1690.380 ;
        RECT 1824.905 1690.195 1825.195 1690.240 ;
        RECT 1824.905 1687.660 1825.195 1687.705 ;
        RECT 2297.770 1687.660 2298.090 1687.720 ;
        RECT 1824.905 1687.520 2298.090 1687.660 ;
        RECT 1824.905 1687.475 1825.195 1687.520 ;
        RECT 2297.770 1687.460 2298.090 1687.520 ;
        RECT 2297.770 35.940 2298.090 36.000 ;
        RECT 2304.210 35.940 2304.530 36.000 ;
        RECT 2297.770 35.800 2304.530 35.940 ;
        RECT 2297.770 35.740 2298.090 35.800 ;
        RECT 2304.210 35.740 2304.530 35.800 ;
      LAYER via ;
        RECT 1774.320 1695.280 1774.580 1695.540 ;
        RECT 2297.800 1687.460 2298.060 1687.720 ;
        RECT 2297.800 35.740 2298.060 36.000 ;
        RECT 2304.240 35.740 2304.500 36.000 ;
      LAYER met2 ;
        RECT 1774.310 1700.000 1774.590 1704.000 ;
        RECT 1774.380 1695.570 1774.520 1700.000 ;
        RECT 1774.320 1695.250 1774.580 1695.570 ;
        RECT 2297.800 1687.430 2298.060 1687.750 ;
        RECT 2297.860 36.030 2298.000 1687.430 ;
        RECT 2297.800 35.710 2298.060 36.030 ;
        RECT 2304.240 35.710 2304.500 36.030 ;
        RECT 2304.300 2.400 2304.440 35.710 ;
>>>>>>> re-updated local openlane
        RECT 2304.090 -4.800 2304.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1779.810 20.300 1780.130 20.360 ;
        RECT 2322.150 20.300 2322.470 20.360 ;
        RECT 1779.810 20.160 2322.470 20.300 ;
        RECT 1779.810 20.100 1780.130 20.160 ;
        RECT 2322.150 20.100 2322.470 20.160 ;
      LAYER via ;
        RECT 1779.840 20.100 1780.100 20.360 ;
        RECT 2322.180 20.100 2322.440 20.360 ;
      LAYER met2 ;
        RECT 1779.370 1700.410 1779.650 1704.000 ;
        RECT 1779.370 1700.270 1780.040 1700.410 ;
        RECT 1779.370 1700.000 1779.650 1700.270 ;
        RECT 1779.900 20.390 1780.040 1700.270 ;
        RECT 1779.840 20.070 1780.100 20.390 ;
        RECT 2322.180 20.070 2322.440 20.390 ;
        RECT 2322.240 2.400 2322.380 20.070 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 0.300 ;
=======
      LAYER li1 ;
        RECT 2339.245 48.365 2339.415 96.475 ;
      LAYER mcon ;
        RECT 2339.245 96.305 2339.415 96.475 ;
      LAYER met1 ;
        RECT 1783.950 1687.320 1784.270 1687.380 ;
        RECT 2339.170 1687.320 2339.490 1687.380 ;
        RECT 1783.950 1687.180 2339.490 1687.320 ;
        RECT 1783.950 1687.120 1784.270 1687.180 ;
        RECT 2339.170 1687.120 2339.490 1687.180 ;
        RECT 2339.170 96.460 2339.490 96.520 ;
        RECT 2338.975 96.320 2339.490 96.460 ;
        RECT 2339.170 96.260 2339.490 96.320 ;
        RECT 2339.185 48.520 2339.475 48.565 ;
        RECT 2339.630 48.520 2339.950 48.580 ;
        RECT 2339.185 48.380 2339.950 48.520 ;
        RECT 2339.185 48.335 2339.475 48.380 ;
        RECT 2339.630 48.320 2339.950 48.380 ;
      LAYER via ;
        RECT 1783.980 1687.120 1784.240 1687.380 ;
        RECT 2339.200 1687.120 2339.460 1687.380 ;
        RECT 2339.200 96.260 2339.460 96.520 ;
        RECT 2339.660 48.320 2339.920 48.580 ;
      LAYER met2 ;
        RECT 1783.970 1700.000 1784.250 1704.000 ;
        RECT 1784.040 1687.410 1784.180 1700.000 ;
        RECT 1783.980 1687.090 1784.240 1687.410 ;
        RECT 2339.200 1687.090 2339.460 1687.410 ;
        RECT 2339.260 96.550 2339.400 1687.090 ;
        RECT 2339.200 96.230 2339.460 96.550 ;
        RECT 2339.660 48.290 2339.920 48.610 ;
        RECT 2339.720 2.400 2339.860 48.290 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 0.300 ;
=======
      LAYER met1 ;
        RECT 1789.010 1684.940 1789.330 1685.000 ;
        RECT 1793.610 1684.940 1793.930 1685.000 ;
        RECT 1789.010 1684.800 1793.930 1684.940 ;
        RECT 1789.010 1684.740 1789.330 1684.800 ;
        RECT 1793.610 1684.740 1793.930 1684.800 ;
        RECT 1793.610 19.960 1793.930 20.020 ;
        RECT 2357.570 19.960 2357.890 20.020 ;
        RECT 1793.610 19.820 2357.890 19.960 ;
        RECT 1793.610 19.760 1793.930 19.820 ;
        RECT 2357.570 19.760 2357.890 19.820 ;
      LAYER via ;
        RECT 1789.040 1684.740 1789.300 1685.000 ;
        RECT 1793.640 1684.740 1793.900 1685.000 ;
        RECT 1793.640 19.760 1793.900 20.020 ;
        RECT 2357.600 19.760 2357.860 20.020 ;
      LAYER met2 ;
        RECT 1789.030 1700.000 1789.310 1704.000 ;
        RECT 1789.100 1685.030 1789.240 1700.000 ;
        RECT 1789.040 1684.710 1789.300 1685.030 ;
        RECT 1793.640 1684.710 1793.900 1685.030 ;
        RECT 1793.700 20.050 1793.840 1684.710 ;
        RECT 1793.640 19.730 1793.900 20.050 ;
        RECT 2357.600 19.730 2357.860 20.050 ;
        RECT 2357.660 2.400 2357.800 19.730 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 0.300 ;
=======
      LAYER li1 ;
        RECT 2373.745 1635.485 2373.915 1683.595 ;
        RECT 2373.745 1538.925 2373.915 1587.035 ;
        RECT 2373.745 1442.025 2373.915 1490.475 ;
        RECT 2373.745 766.105 2373.915 814.215 ;
        RECT 2373.745 669.545 2373.915 717.655 ;
        RECT 2373.745 572.645 2373.915 620.755 ;
        RECT 2373.745 476.085 2373.915 524.195 ;
        RECT 2373.745 379.525 2373.915 427.635 ;
        RECT 2373.745 282.965 2373.915 331.075 ;
        RECT 2373.745 186.405 2373.915 234.515 ;
        RECT 2373.745 89.845 2373.915 137.955 ;
      LAYER mcon ;
        RECT 2373.745 1683.425 2373.915 1683.595 ;
        RECT 2373.745 1586.865 2373.915 1587.035 ;
        RECT 2373.745 1490.305 2373.915 1490.475 ;
        RECT 2373.745 814.045 2373.915 814.215 ;
        RECT 2373.745 717.485 2373.915 717.655 ;
        RECT 2373.745 620.585 2373.915 620.755 ;
        RECT 2373.745 524.025 2373.915 524.195 ;
        RECT 2373.745 427.465 2373.915 427.635 ;
        RECT 2373.745 330.905 2373.915 331.075 ;
        RECT 2373.745 234.345 2373.915 234.515 ;
        RECT 2373.745 137.785 2373.915 137.955 ;
      LAYER met1 ;
        RECT 1793.610 1686.980 1793.930 1687.040 ;
        RECT 2373.670 1686.980 2373.990 1687.040 ;
        RECT 1793.610 1686.840 2373.990 1686.980 ;
        RECT 1793.610 1686.780 1793.930 1686.840 ;
        RECT 2373.670 1686.780 2373.990 1686.840 ;
        RECT 2373.670 1683.580 2373.990 1683.640 ;
        RECT 2373.475 1683.440 2373.990 1683.580 ;
        RECT 2373.670 1683.380 2373.990 1683.440 ;
        RECT 2373.670 1635.640 2373.990 1635.700 ;
        RECT 2373.475 1635.500 2373.990 1635.640 ;
        RECT 2373.670 1635.440 2373.990 1635.500 ;
        RECT 2373.670 1587.020 2373.990 1587.080 ;
        RECT 2373.475 1586.880 2373.990 1587.020 ;
        RECT 2373.670 1586.820 2373.990 1586.880 ;
        RECT 2373.670 1539.080 2373.990 1539.140 ;
        RECT 2373.475 1538.940 2373.990 1539.080 ;
        RECT 2373.670 1538.880 2373.990 1538.940 ;
        RECT 2373.670 1490.460 2373.990 1490.520 ;
        RECT 2373.475 1490.320 2373.990 1490.460 ;
        RECT 2373.670 1490.260 2373.990 1490.320 ;
        RECT 2373.670 1442.180 2373.990 1442.240 ;
        RECT 2373.475 1442.040 2373.990 1442.180 ;
        RECT 2373.670 1441.980 2373.990 1442.040 ;
        RECT 2373.670 1345.620 2373.990 1345.680 ;
        RECT 2374.590 1345.620 2374.910 1345.680 ;
        RECT 2373.670 1345.480 2374.910 1345.620 ;
        RECT 2373.670 1345.420 2373.990 1345.480 ;
        RECT 2374.590 1345.420 2374.910 1345.480 ;
        RECT 2373.670 1249.060 2373.990 1249.120 ;
        RECT 2374.590 1249.060 2374.910 1249.120 ;
        RECT 2373.670 1248.920 2374.910 1249.060 ;
        RECT 2373.670 1248.860 2373.990 1248.920 ;
        RECT 2374.590 1248.860 2374.910 1248.920 ;
        RECT 2373.670 1152.500 2373.990 1152.560 ;
        RECT 2374.590 1152.500 2374.910 1152.560 ;
        RECT 2373.670 1152.360 2374.910 1152.500 ;
        RECT 2373.670 1152.300 2373.990 1152.360 ;
        RECT 2374.590 1152.300 2374.910 1152.360 ;
        RECT 2373.670 1007.320 2373.990 1007.380 ;
        RECT 2374.590 1007.320 2374.910 1007.380 ;
        RECT 2373.670 1007.180 2374.910 1007.320 ;
        RECT 2373.670 1007.120 2373.990 1007.180 ;
        RECT 2374.590 1007.120 2374.910 1007.180 ;
        RECT 2373.670 910.760 2373.990 910.820 ;
        RECT 2374.590 910.760 2374.910 910.820 ;
        RECT 2373.670 910.620 2374.910 910.760 ;
        RECT 2373.670 910.560 2373.990 910.620 ;
        RECT 2374.590 910.560 2374.910 910.620 ;
        RECT 2373.670 814.200 2373.990 814.260 ;
        RECT 2373.475 814.060 2373.990 814.200 ;
        RECT 2373.670 814.000 2373.990 814.060 ;
        RECT 2373.670 766.260 2373.990 766.320 ;
        RECT 2373.475 766.120 2373.990 766.260 ;
        RECT 2373.670 766.060 2373.990 766.120 ;
        RECT 2373.670 717.640 2373.990 717.700 ;
        RECT 2373.475 717.500 2373.990 717.640 ;
        RECT 2373.670 717.440 2373.990 717.500 ;
        RECT 2373.670 669.700 2373.990 669.760 ;
        RECT 2373.475 669.560 2373.990 669.700 ;
        RECT 2373.670 669.500 2373.990 669.560 ;
        RECT 2373.670 620.740 2373.990 620.800 ;
        RECT 2373.475 620.600 2373.990 620.740 ;
        RECT 2373.670 620.540 2373.990 620.600 ;
        RECT 2373.670 572.800 2373.990 572.860 ;
        RECT 2373.475 572.660 2373.990 572.800 ;
        RECT 2373.670 572.600 2373.990 572.660 ;
        RECT 2373.670 524.180 2373.990 524.240 ;
        RECT 2373.475 524.040 2373.990 524.180 ;
        RECT 2373.670 523.980 2373.990 524.040 ;
        RECT 2373.670 476.240 2373.990 476.300 ;
        RECT 2373.475 476.100 2373.990 476.240 ;
        RECT 2373.670 476.040 2373.990 476.100 ;
        RECT 2373.670 427.620 2373.990 427.680 ;
        RECT 2373.475 427.480 2373.990 427.620 ;
        RECT 2373.670 427.420 2373.990 427.480 ;
        RECT 2373.670 379.680 2373.990 379.740 ;
        RECT 2373.475 379.540 2373.990 379.680 ;
        RECT 2373.670 379.480 2373.990 379.540 ;
        RECT 2373.670 331.060 2373.990 331.120 ;
        RECT 2373.475 330.920 2373.990 331.060 ;
        RECT 2373.670 330.860 2373.990 330.920 ;
        RECT 2373.670 283.120 2373.990 283.180 ;
        RECT 2373.475 282.980 2373.990 283.120 ;
        RECT 2373.670 282.920 2373.990 282.980 ;
        RECT 2373.670 234.500 2373.990 234.560 ;
        RECT 2373.475 234.360 2373.990 234.500 ;
        RECT 2373.670 234.300 2373.990 234.360 ;
        RECT 2373.670 186.560 2373.990 186.620 ;
        RECT 2373.475 186.420 2373.990 186.560 ;
        RECT 2373.670 186.360 2373.990 186.420 ;
        RECT 2373.670 137.940 2373.990 138.000 ;
        RECT 2373.475 137.800 2373.990 137.940 ;
        RECT 2373.670 137.740 2373.990 137.800 ;
        RECT 2373.670 90.000 2373.990 90.060 ;
        RECT 2373.475 89.860 2373.990 90.000 ;
        RECT 2373.670 89.800 2373.990 89.860 ;
        RECT 2373.210 48.520 2373.530 48.580 ;
        RECT 2374.590 48.520 2374.910 48.580 ;
        RECT 2373.210 48.380 2374.910 48.520 ;
        RECT 2373.210 48.320 2373.530 48.380 ;
        RECT 2374.590 48.320 2374.910 48.380 ;
      LAYER via ;
        RECT 1793.640 1686.780 1793.900 1687.040 ;
        RECT 2373.700 1686.780 2373.960 1687.040 ;
        RECT 2373.700 1683.380 2373.960 1683.640 ;
        RECT 2373.700 1635.440 2373.960 1635.700 ;
        RECT 2373.700 1586.820 2373.960 1587.080 ;
        RECT 2373.700 1538.880 2373.960 1539.140 ;
        RECT 2373.700 1490.260 2373.960 1490.520 ;
        RECT 2373.700 1441.980 2373.960 1442.240 ;
        RECT 2373.700 1345.420 2373.960 1345.680 ;
        RECT 2374.620 1345.420 2374.880 1345.680 ;
        RECT 2373.700 1248.860 2373.960 1249.120 ;
        RECT 2374.620 1248.860 2374.880 1249.120 ;
        RECT 2373.700 1152.300 2373.960 1152.560 ;
        RECT 2374.620 1152.300 2374.880 1152.560 ;
        RECT 2373.700 1007.120 2373.960 1007.380 ;
        RECT 2374.620 1007.120 2374.880 1007.380 ;
        RECT 2373.700 910.560 2373.960 910.820 ;
        RECT 2374.620 910.560 2374.880 910.820 ;
        RECT 2373.700 814.000 2373.960 814.260 ;
        RECT 2373.700 766.060 2373.960 766.320 ;
        RECT 2373.700 717.440 2373.960 717.700 ;
        RECT 2373.700 669.500 2373.960 669.760 ;
        RECT 2373.700 620.540 2373.960 620.800 ;
        RECT 2373.700 572.600 2373.960 572.860 ;
        RECT 2373.700 523.980 2373.960 524.240 ;
        RECT 2373.700 476.040 2373.960 476.300 ;
        RECT 2373.700 427.420 2373.960 427.680 ;
        RECT 2373.700 379.480 2373.960 379.740 ;
        RECT 2373.700 330.860 2373.960 331.120 ;
        RECT 2373.700 282.920 2373.960 283.180 ;
        RECT 2373.700 234.300 2373.960 234.560 ;
        RECT 2373.700 186.360 2373.960 186.620 ;
        RECT 2373.700 137.740 2373.960 138.000 ;
        RECT 2373.700 89.800 2373.960 90.060 ;
        RECT 2373.240 48.320 2373.500 48.580 ;
        RECT 2374.620 48.320 2374.880 48.580 ;
      LAYER met2 ;
        RECT 1793.630 1700.000 1793.910 1704.000 ;
        RECT 1793.700 1687.070 1793.840 1700.000 ;
        RECT 1793.640 1686.750 1793.900 1687.070 ;
        RECT 2373.700 1686.750 2373.960 1687.070 ;
        RECT 2373.760 1683.670 2373.900 1686.750 ;
        RECT 2373.700 1683.350 2373.960 1683.670 ;
        RECT 2373.700 1635.410 2373.960 1635.730 ;
        RECT 2373.760 1587.110 2373.900 1635.410 ;
        RECT 2373.700 1586.790 2373.960 1587.110 ;
        RECT 2373.700 1538.850 2373.960 1539.170 ;
        RECT 2373.760 1490.550 2373.900 1538.850 ;
        RECT 2373.700 1490.230 2373.960 1490.550 ;
        RECT 2373.700 1441.950 2373.960 1442.270 ;
        RECT 2373.760 1393.845 2373.900 1441.950 ;
        RECT 2373.690 1393.475 2373.970 1393.845 ;
        RECT 2374.610 1393.475 2374.890 1393.845 ;
        RECT 2374.680 1345.710 2374.820 1393.475 ;
        RECT 2373.700 1345.390 2373.960 1345.710 ;
        RECT 2374.620 1345.390 2374.880 1345.710 ;
        RECT 2373.760 1297.285 2373.900 1345.390 ;
        RECT 2373.690 1296.915 2373.970 1297.285 ;
        RECT 2374.610 1296.915 2374.890 1297.285 ;
        RECT 2374.680 1249.150 2374.820 1296.915 ;
        RECT 2373.700 1248.830 2373.960 1249.150 ;
        RECT 2374.620 1248.830 2374.880 1249.150 ;
        RECT 2373.760 1200.725 2373.900 1248.830 ;
        RECT 2373.690 1200.355 2373.970 1200.725 ;
        RECT 2374.610 1200.355 2374.890 1200.725 ;
        RECT 2374.680 1152.590 2374.820 1200.355 ;
        RECT 2373.700 1152.270 2373.960 1152.590 ;
        RECT 2374.620 1152.270 2374.880 1152.590 ;
        RECT 2373.760 1104.165 2373.900 1152.270 ;
        RECT 2373.690 1103.795 2373.970 1104.165 ;
        RECT 2374.610 1103.795 2374.890 1104.165 ;
        RECT 2374.680 1055.885 2374.820 1103.795 ;
        RECT 2373.690 1055.515 2373.970 1055.885 ;
        RECT 2374.610 1055.515 2374.890 1055.885 ;
        RECT 2373.760 1007.410 2373.900 1055.515 ;
        RECT 2373.700 1007.090 2373.960 1007.410 ;
        RECT 2374.620 1007.090 2374.880 1007.410 ;
        RECT 2374.680 959.325 2374.820 1007.090 ;
        RECT 2373.690 958.955 2373.970 959.325 ;
        RECT 2374.610 958.955 2374.890 959.325 ;
        RECT 2373.760 910.850 2373.900 958.955 ;
        RECT 2373.700 910.530 2373.960 910.850 ;
        RECT 2374.620 910.530 2374.880 910.850 ;
        RECT 2374.680 862.765 2374.820 910.530 ;
        RECT 2373.690 862.395 2373.970 862.765 ;
        RECT 2374.610 862.395 2374.890 862.765 ;
        RECT 2373.760 814.290 2373.900 862.395 ;
        RECT 2373.700 813.970 2373.960 814.290 ;
        RECT 2373.700 766.030 2373.960 766.350 ;
        RECT 2373.760 717.730 2373.900 766.030 ;
        RECT 2373.700 717.410 2373.960 717.730 ;
        RECT 2373.700 669.470 2373.960 669.790 ;
        RECT 2373.760 620.830 2373.900 669.470 ;
        RECT 2373.700 620.510 2373.960 620.830 ;
        RECT 2373.700 572.570 2373.960 572.890 ;
        RECT 2373.760 524.270 2373.900 572.570 ;
        RECT 2373.700 523.950 2373.960 524.270 ;
        RECT 2373.700 476.010 2373.960 476.330 ;
        RECT 2373.760 427.710 2373.900 476.010 ;
        RECT 2373.700 427.390 2373.960 427.710 ;
        RECT 2373.700 379.450 2373.960 379.770 ;
        RECT 2373.760 331.150 2373.900 379.450 ;
        RECT 2373.700 330.830 2373.960 331.150 ;
        RECT 2373.700 282.890 2373.960 283.210 ;
        RECT 2373.760 234.590 2373.900 282.890 ;
        RECT 2373.700 234.270 2373.960 234.590 ;
        RECT 2373.700 186.330 2373.960 186.650 ;
        RECT 2373.760 138.030 2373.900 186.330 ;
        RECT 2373.700 137.710 2373.960 138.030 ;
        RECT 2373.700 89.770 2373.960 90.090 ;
        RECT 2373.760 72.490 2373.900 89.770 ;
        RECT 2373.300 72.350 2373.900 72.490 ;
        RECT 2373.300 48.610 2373.440 72.350 ;
        RECT 2373.240 48.290 2373.500 48.610 ;
        RECT 2374.620 48.290 2374.880 48.610 ;
        RECT 2374.680 24.210 2374.820 48.290 ;
        RECT 2374.680 24.070 2375.740 24.210 ;
        RECT 2375.600 2.400 2375.740 24.070 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
<<<<<<< HEAD
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER via2 ;
        RECT 2373.690 1393.520 2373.970 1393.800 ;
        RECT 2374.610 1393.520 2374.890 1393.800 ;
        RECT 2373.690 1296.960 2373.970 1297.240 ;
        RECT 2374.610 1296.960 2374.890 1297.240 ;
        RECT 2373.690 1200.400 2373.970 1200.680 ;
        RECT 2374.610 1200.400 2374.890 1200.680 ;
        RECT 2373.690 1103.840 2373.970 1104.120 ;
        RECT 2374.610 1103.840 2374.890 1104.120 ;
        RECT 2373.690 1055.560 2373.970 1055.840 ;
        RECT 2374.610 1055.560 2374.890 1055.840 ;
        RECT 2373.690 959.000 2373.970 959.280 ;
        RECT 2374.610 959.000 2374.890 959.280 ;
        RECT 2373.690 862.440 2373.970 862.720 ;
        RECT 2374.610 862.440 2374.890 862.720 ;
      LAYER met3 ;
        RECT 2373.665 1393.810 2373.995 1393.825 ;
        RECT 2374.585 1393.810 2374.915 1393.825 ;
        RECT 2373.665 1393.510 2374.915 1393.810 ;
        RECT 2373.665 1393.495 2373.995 1393.510 ;
        RECT 2374.585 1393.495 2374.915 1393.510 ;
        RECT 2373.665 1297.250 2373.995 1297.265 ;
        RECT 2374.585 1297.250 2374.915 1297.265 ;
        RECT 2373.665 1296.950 2374.915 1297.250 ;
        RECT 2373.665 1296.935 2373.995 1296.950 ;
        RECT 2374.585 1296.935 2374.915 1296.950 ;
        RECT 2373.665 1200.690 2373.995 1200.705 ;
        RECT 2374.585 1200.690 2374.915 1200.705 ;
        RECT 2373.665 1200.390 2374.915 1200.690 ;
        RECT 2373.665 1200.375 2373.995 1200.390 ;
        RECT 2374.585 1200.375 2374.915 1200.390 ;
        RECT 2373.665 1104.130 2373.995 1104.145 ;
        RECT 2374.585 1104.130 2374.915 1104.145 ;
        RECT 2373.665 1103.830 2374.915 1104.130 ;
        RECT 2373.665 1103.815 2373.995 1103.830 ;
        RECT 2374.585 1103.815 2374.915 1103.830 ;
        RECT 2373.665 1055.850 2373.995 1055.865 ;
        RECT 2374.585 1055.850 2374.915 1055.865 ;
        RECT 2373.665 1055.550 2374.915 1055.850 ;
        RECT 2373.665 1055.535 2373.995 1055.550 ;
        RECT 2374.585 1055.535 2374.915 1055.550 ;
        RECT 2373.665 959.290 2373.995 959.305 ;
        RECT 2374.585 959.290 2374.915 959.305 ;
        RECT 2373.665 958.990 2374.915 959.290 ;
        RECT 2373.665 958.975 2373.995 958.990 ;
        RECT 2374.585 958.975 2374.915 958.990 ;
        RECT 2373.665 862.730 2373.995 862.745 ;
        RECT 2374.585 862.730 2374.915 862.745 ;
        RECT 2373.665 862.430 2374.915 862.730 ;
        RECT 2373.665 862.415 2373.995 862.430 ;
        RECT 2374.585 862.415 2374.915 862.430 ;
>>>>>>> re-updated local openlane
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 0.300 ;
=======
      LAYER met1 ;
        RECT 1798.670 1683.920 1798.990 1683.980 ;
        RECT 1800.510 1683.920 1800.830 1683.980 ;
        RECT 1798.670 1683.780 1800.830 1683.920 ;
        RECT 1798.670 1683.720 1798.990 1683.780 ;
        RECT 1800.510 1683.720 1800.830 1683.780 ;
        RECT 1800.510 19.620 1800.830 19.680 ;
        RECT 2393.450 19.620 2393.770 19.680 ;
        RECT 1800.510 19.480 2393.770 19.620 ;
        RECT 1800.510 19.420 1800.830 19.480 ;
        RECT 2393.450 19.420 2393.770 19.480 ;
      LAYER via ;
        RECT 1798.700 1683.720 1798.960 1683.980 ;
        RECT 1800.540 1683.720 1800.800 1683.980 ;
        RECT 1800.540 19.420 1800.800 19.680 ;
        RECT 2393.480 19.420 2393.740 19.680 ;
      LAYER met2 ;
        RECT 1798.690 1700.000 1798.970 1704.000 ;
        RECT 1798.760 1684.010 1798.900 1700.000 ;
        RECT 1798.700 1683.690 1798.960 1684.010 ;
        RECT 1800.540 1683.690 1800.800 1684.010 ;
        RECT 1800.600 19.710 1800.740 1683.690 ;
        RECT 1800.540 19.390 1800.800 19.710 ;
        RECT 2393.480 19.390 2393.740 19.710 ;
        RECT 2393.540 2.400 2393.680 19.390 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 0.300 ;
=======
      LAYER met1 ;
        RECT 1803.270 1683.920 1803.590 1683.980 ;
        RECT 1806.030 1683.920 1806.350 1683.980 ;
        RECT 1803.270 1683.780 1806.350 1683.920 ;
        RECT 1803.270 1683.720 1803.590 1683.780 ;
        RECT 1806.030 1683.720 1806.350 1683.780 ;
        RECT 1806.030 19.280 1806.350 19.340 ;
        RECT 2411.390 19.280 2411.710 19.340 ;
        RECT 1806.030 19.140 2411.710 19.280 ;
        RECT 1806.030 19.080 1806.350 19.140 ;
        RECT 2411.390 19.080 2411.710 19.140 ;
      LAYER via ;
        RECT 1803.300 1683.720 1803.560 1683.980 ;
        RECT 1806.060 1683.720 1806.320 1683.980 ;
        RECT 1806.060 19.080 1806.320 19.340 ;
        RECT 2411.420 19.080 2411.680 19.340 ;
      LAYER met2 ;
        RECT 1803.290 1700.000 1803.570 1704.000 ;
        RECT 1803.360 1684.010 1803.500 1700.000 ;
        RECT 1803.300 1683.690 1803.560 1684.010 ;
        RECT 1806.060 1683.690 1806.320 1684.010 ;
        RECT 1806.120 19.370 1806.260 1683.690 ;
        RECT 1806.060 19.050 1806.320 19.370 ;
        RECT 2411.420 19.050 2411.680 19.370 ;
        RECT 2411.480 2.400 2411.620 19.050 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 0.300 ;
=======
      LAYER met1 ;
        RECT 805.530 43.080 805.850 43.140 ;
        RECT 1367.650 43.080 1367.970 43.140 ;
        RECT 805.530 42.940 1367.970 43.080 ;
        RECT 805.530 42.880 805.850 42.940 ;
        RECT 1367.650 42.880 1367.970 42.940 ;
      LAYER via ;
        RECT 805.560 42.880 805.820 43.140 ;
        RECT 1367.680 42.880 1367.940 43.140 ;
      LAYER met2 ;
        RECT 1368.130 1700.410 1368.410 1704.000 ;
        RECT 1367.740 1700.270 1368.410 1700.410 ;
        RECT 1367.740 43.170 1367.880 1700.270 ;
        RECT 1368.130 1700.000 1368.410 1700.270 ;
        RECT 805.560 42.850 805.820 43.170 ;
        RECT 1367.680 42.850 1367.940 43.170 ;
        RECT 805.620 2.400 805.760 42.850 ;
        RECT 805.410 -4.800 805.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 0.300 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 0.300 ;
=======
      LAYER met1 ;
        RECT 2.830 24.040 3.150 24.100 ;
        RECT 1145.930 24.040 1146.250 24.100 ;
        RECT 2.830 23.900 1146.250 24.040 ;
        RECT 2.830 23.840 3.150 23.900 ;
        RECT 1145.930 23.840 1146.250 23.900 ;
      LAYER via ;
        RECT 2.860 23.840 3.120 24.100 ;
        RECT 1145.960 23.840 1146.220 24.100 ;
      LAYER met2 ;
        RECT 1150.550 1700.410 1150.830 1704.000 ;
        RECT 1146.020 1700.270 1150.830 1700.410 ;
        RECT 1146.020 24.130 1146.160 1700.270 ;
        RECT 1150.550 1700.000 1150.830 1700.270 ;
        RECT 2.860 23.810 3.120 24.130 ;
        RECT 1145.960 23.810 1146.220 24.130 ;
        RECT 2.920 2.400 3.060 23.810 ;
        RECT 2.710 -4.800 3.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 0.300 ;
=======
      LAYER li1 ;
        RECT 1147.385 1510.365 1147.555 1579.895 ;
        RECT 1146.465 1400.885 1146.635 1463.615 ;
        RECT 1147.385 1352.605 1147.555 1376.915 ;
        RECT 1146.925 1268.965 1147.095 1304.155 ;
        RECT 1146.465 917.745 1146.635 961.775 ;
        RECT 1146.465 531.505 1146.635 579.615 ;
        RECT 1146.465 434.945 1146.635 483.055 ;
        RECT 1146.465 338.045 1146.635 386.155 ;
        RECT 1146.465 241.485 1146.635 289.255 ;
        RECT 1146.925 193.205 1147.095 207.655 ;
        RECT 1146.005 138.125 1146.175 162.095 ;
      LAYER mcon ;
        RECT 1147.385 1579.725 1147.555 1579.895 ;
        RECT 1146.465 1463.445 1146.635 1463.615 ;
        RECT 1147.385 1376.745 1147.555 1376.915 ;
        RECT 1146.925 1303.985 1147.095 1304.155 ;
        RECT 1146.465 961.605 1146.635 961.775 ;
        RECT 1146.465 579.445 1146.635 579.615 ;
        RECT 1146.465 482.885 1146.635 483.055 ;
        RECT 1146.465 385.985 1146.635 386.155 ;
        RECT 1146.465 289.085 1146.635 289.255 ;
        RECT 1146.925 207.485 1147.095 207.655 ;
        RECT 1146.005 161.925 1146.175 162.095 ;
      LAYER met1 ;
        RECT 1147.310 1676.780 1147.630 1676.840 ;
        RECT 1151.910 1676.780 1152.230 1676.840 ;
        RECT 1147.310 1676.640 1152.230 1676.780 ;
        RECT 1147.310 1676.580 1147.630 1676.640 ;
        RECT 1151.910 1676.580 1152.230 1676.640 ;
        RECT 1146.390 1580.560 1146.710 1580.620 ;
        RECT 1147.310 1580.560 1147.630 1580.620 ;
        RECT 1146.390 1580.420 1147.630 1580.560 ;
        RECT 1146.390 1580.360 1146.710 1580.420 ;
        RECT 1147.310 1580.360 1147.630 1580.420 ;
        RECT 1147.310 1579.880 1147.630 1579.940 ;
        RECT 1147.115 1579.740 1147.630 1579.880 ;
        RECT 1147.310 1579.680 1147.630 1579.740 ;
        RECT 1147.310 1510.520 1147.630 1510.580 ;
        RECT 1147.115 1510.380 1147.630 1510.520 ;
        RECT 1147.310 1510.320 1147.630 1510.380 ;
        RECT 1146.405 1463.600 1146.695 1463.645 ;
        RECT 1147.310 1463.600 1147.630 1463.660 ;
        RECT 1146.405 1463.460 1147.630 1463.600 ;
        RECT 1146.405 1463.415 1146.695 1463.460 ;
        RECT 1147.310 1463.400 1147.630 1463.460 ;
        RECT 1146.405 1401.040 1146.695 1401.085 ;
        RECT 1147.310 1401.040 1147.630 1401.100 ;
        RECT 1146.405 1400.900 1147.630 1401.040 ;
        RECT 1146.405 1400.855 1146.695 1400.900 ;
        RECT 1147.310 1400.840 1147.630 1400.900 ;
        RECT 1147.310 1376.900 1147.630 1376.960 ;
        RECT 1147.115 1376.760 1147.630 1376.900 ;
        RECT 1147.310 1376.700 1147.630 1376.760 ;
        RECT 1146.390 1352.760 1146.710 1352.820 ;
        RECT 1147.325 1352.760 1147.615 1352.805 ;
        RECT 1146.390 1352.620 1147.615 1352.760 ;
        RECT 1146.390 1352.560 1146.710 1352.620 ;
        RECT 1147.325 1352.575 1147.615 1352.620 ;
        RECT 1146.390 1317.880 1146.710 1318.140 ;
        RECT 1146.480 1317.740 1146.620 1317.880 ;
        RECT 1146.850 1317.740 1147.170 1317.800 ;
        RECT 1146.480 1317.600 1147.170 1317.740 ;
        RECT 1146.850 1317.540 1147.170 1317.600 ;
        RECT 1146.850 1304.140 1147.170 1304.200 ;
        RECT 1146.655 1304.000 1147.170 1304.140 ;
        RECT 1146.850 1303.940 1147.170 1304.000 ;
        RECT 1146.850 1269.120 1147.170 1269.180 ;
        RECT 1146.655 1268.980 1147.170 1269.120 ;
        RECT 1146.850 1268.920 1147.170 1268.980 ;
        RECT 1146.850 1221.860 1147.170 1221.920 ;
        RECT 1146.480 1221.720 1147.170 1221.860 ;
        RECT 1146.480 1221.240 1146.620 1221.720 ;
        RECT 1146.850 1221.660 1147.170 1221.720 ;
        RECT 1146.390 1220.980 1146.710 1221.240 ;
        RECT 1146.850 1152.500 1147.170 1152.560 ;
        RECT 1147.770 1152.500 1148.090 1152.560 ;
        RECT 1146.850 1152.360 1148.090 1152.500 ;
        RECT 1146.850 1152.300 1147.170 1152.360 ;
        RECT 1147.770 1152.300 1148.090 1152.360 ;
        RECT 1146.850 1125.300 1147.170 1125.360 ;
        RECT 1146.480 1125.160 1147.170 1125.300 ;
        RECT 1146.480 1124.680 1146.620 1125.160 ;
        RECT 1146.850 1125.100 1147.170 1125.160 ;
        RECT 1146.390 1124.420 1146.710 1124.680 ;
        RECT 1147.310 1027.720 1147.630 1027.780 ;
        RECT 1148.230 1027.720 1148.550 1027.780 ;
        RECT 1147.310 1027.580 1148.550 1027.720 ;
        RECT 1147.310 1027.520 1147.630 1027.580 ;
        RECT 1148.230 1027.520 1148.550 1027.580 ;
        RECT 1146.390 980.120 1146.710 980.180 ;
        RECT 1147.310 980.120 1147.630 980.180 ;
        RECT 1146.390 979.980 1147.630 980.120 ;
        RECT 1146.390 979.920 1146.710 979.980 ;
        RECT 1147.310 979.920 1147.630 979.980 ;
        RECT 1146.390 961.760 1146.710 961.820 ;
        RECT 1146.195 961.620 1146.710 961.760 ;
        RECT 1146.390 961.560 1146.710 961.620 ;
        RECT 1146.405 917.900 1146.695 917.945 ;
        RECT 1146.850 917.900 1147.170 917.960 ;
        RECT 1146.405 917.760 1147.170 917.900 ;
        RECT 1146.405 917.715 1146.695 917.760 ;
        RECT 1146.850 917.700 1147.170 917.760 ;
        RECT 1146.850 883.700 1147.170 883.960 ;
        RECT 1146.940 882.940 1147.080 883.700 ;
        RECT 1146.850 882.680 1147.170 882.940 ;
        RECT 1146.390 786.800 1146.710 787.060 ;
        RECT 1146.480 786.660 1146.620 786.800 ;
        RECT 1146.850 786.660 1147.170 786.720 ;
        RECT 1146.480 786.520 1147.170 786.660 ;
        RECT 1146.850 786.460 1147.170 786.520 ;
        RECT 1146.850 772.720 1147.170 772.780 ;
        RECT 1147.770 772.720 1148.090 772.780 ;
        RECT 1146.850 772.580 1148.090 772.720 ;
        RECT 1146.850 772.520 1147.170 772.580 ;
        RECT 1147.770 772.520 1148.090 772.580 ;
        RECT 1146.390 689.900 1146.710 690.160 ;
        RECT 1146.480 689.760 1146.620 689.900 ;
        RECT 1146.850 689.760 1147.170 689.820 ;
        RECT 1146.480 689.620 1147.170 689.760 ;
        RECT 1146.850 689.560 1147.170 689.620 ;
        RECT 1146.850 676.160 1147.170 676.220 ;
        RECT 1147.770 676.160 1148.090 676.220 ;
        RECT 1146.850 676.020 1148.090 676.160 ;
        RECT 1146.850 675.960 1147.170 676.020 ;
        RECT 1147.770 675.960 1148.090 676.020 ;
        RECT 1146.390 593.340 1146.710 593.600 ;
        RECT 1146.480 593.200 1146.620 593.340 ;
        RECT 1146.850 593.200 1147.170 593.260 ;
        RECT 1146.480 593.060 1147.170 593.200 ;
        RECT 1146.850 593.000 1147.170 593.060 ;
        RECT 1146.405 579.600 1146.695 579.645 ;
        RECT 1146.850 579.600 1147.170 579.660 ;
        RECT 1146.405 579.460 1147.170 579.600 ;
        RECT 1146.405 579.415 1146.695 579.460 ;
        RECT 1146.850 579.400 1147.170 579.460 ;
        RECT 1146.390 531.660 1146.710 531.720 ;
        RECT 1146.195 531.520 1146.710 531.660 ;
        RECT 1146.390 531.460 1146.710 531.520 ;
        RECT 1146.390 496.780 1146.710 497.040 ;
        RECT 1146.480 496.640 1146.620 496.780 ;
        RECT 1146.850 496.640 1147.170 496.700 ;
        RECT 1146.480 496.500 1147.170 496.640 ;
        RECT 1146.850 496.440 1147.170 496.500 ;
        RECT 1146.405 483.040 1146.695 483.085 ;
        RECT 1146.850 483.040 1147.170 483.100 ;
        RECT 1146.405 482.900 1147.170 483.040 ;
        RECT 1146.405 482.855 1146.695 482.900 ;
        RECT 1146.850 482.840 1147.170 482.900 ;
        RECT 1146.390 435.100 1146.710 435.160 ;
        RECT 1146.195 434.960 1146.710 435.100 ;
        RECT 1146.390 434.900 1146.710 434.960 ;
        RECT 1146.390 400.220 1146.710 400.480 ;
        RECT 1146.480 399.740 1146.620 400.220 ;
        RECT 1146.850 399.740 1147.170 399.800 ;
        RECT 1146.480 399.600 1147.170 399.740 ;
        RECT 1146.850 399.540 1147.170 399.600 ;
        RECT 1146.405 386.140 1146.695 386.185 ;
        RECT 1146.850 386.140 1147.170 386.200 ;
        RECT 1146.405 386.000 1147.170 386.140 ;
        RECT 1146.405 385.955 1146.695 386.000 ;
        RECT 1146.850 385.940 1147.170 386.000 ;
        RECT 1146.390 338.200 1146.710 338.260 ;
        RECT 1146.195 338.060 1146.710 338.200 ;
        RECT 1146.390 338.000 1146.710 338.060 ;
        RECT 1146.390 289.920 1146.710 289.980 ;
        RECT 1146.850 289.920 1147.170 289.980 ;
        RECT 1146.390 289.780 1147.170 289.920 ;
        RECT 1146.390 289.720 1146.710 289.780 ;
        RECT 1146.850 289.720 1147.170 289.780 ;
        RECT 1146.390 289.240 1146.710 289.300 ;
        RECT 1146.195 289.100 1146.710 289.240 ;
        RECT 1146.390 289.040 1146.710 289.100 ;
        RECT 1146.405 241.640 1146.695 241.685 ;
        RECT 1146.850 241.640 1147.170 241.700 ;
        RECT 1146.405 241.500 1147.170 241.640 ;
        RECT 1146.405 241.455 1146.695 241.500 ;
        RECT 1146.850 241.440 1147.170 241.500 ;
        RECT 1146.850 207.640 1147.170 207.700 ;
        RECT 1146.655 207.500 1147.170 207.640 ;
        RECT 1146.850 207.440 1147.170 207.500 ;
        RECT 1145.930 193.360 1146.250 193.420 ;
        RECT 1146.865 193.360 1147.155 193.405 ;
        RECT 1145.930 193.220 1147.155 193.360 ;
        RECT 1145.930 193.160 1146.250 193.220 ;
        RECT 1146.865 193.175 1147.155 193.220 ;
        RECT 1145.930 162.080 1146.250 162.140 ;
        RECT 1145.735 161.940 1146.250 162.080 ;
        RECT 1145.930 161.880 1146.250 161.940 ;
        RECT 1145.945 138.280 1146.235 138.325 ;
        RECT 1146.850 138.280 1147.170 138.340 ;
        RECT 1145.945 138.140 1147.170 138.280 ;
        RECT 1145.945 138.095 1146.235 138.140 ;
        RECT 1146.850 138.080 1147.170 138.140 ;
        RECT 1146.850 110.740 1147.170 110.800 ;
        RECT 1146.480 110.600 1147.170 110.740 ;
        RECT 1146.480 110.460 1146.620 110.600 ;
        RECT 1146.850 110.540 1147.170 110.600 ;
        RECT 1146.390 110.200 1146.710 110.460 ;
=======
      LAYER met1 ;
        RECT 1145.470 1678.140 1145.790 1678.200 ;
        RECT 1150.990 1678.140 1151.310 1678.200 ;
        RECT 1145.470 1678.000 1151.310 1678.140 ;
        RECT 1145.470 1677.940 1145.790 1678.000 ;
        RECT 1150.990 1677.940 1151.310 1678.000 ;
>>>>>>> re-updated local openlane
        RECT 8.350 24.720 8.670 24.780 ;
        RECT 1145.470 24.720 1145.790 24.780 ;
        RECT 8.350 24.580 1145.790 24.720 ;
        RECT 8.350 24.520 8.670 24.580 ;
        RECT 1145.470 24.520 1145.790 24.580 ;
      LAYER via ;
        RECT 1145.500 1677.940 1145.760 1678.200 ;
        RECT 1151.020 1677.940 1151.280 1678.200 ;
        RECT 8.380 24.520 8.640 24.780 ;
        RECT 1145.500 24.520 1145.760 24.780 ;
      LAYER met2 ;
        RECT 1151.930 1700.410 1152.210 1704.000 ;
        RECT 1151.080 1700.270 1152.210 1700.410 ;
        RECT 1151.080 1678.230 1151.220 1700.270 ;
        RECT 1151.930 1700.000 1152.210 1700.270 ;
        RECT 1145.500 1677.910 1145.760 1678.230 ;
        RECT 1151.020 1677.910 1151.280 1678.230 ;
        RECT 1145.560 24.810 1145.700 1677.910 ;
        RECT 8.380 24.490 8.640 24.810 ;
        RECT 1145.500 24.490 1145.760 24.810 ;
        RECT 8.440 2.400 8.580 24.490 ;
        RECT 8.230 -4.800 8.790 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1146.410 1628.120 1146.690 1628.400 ;
        RECT 1147.330 1628.120 1147.610 1628.400 ;
        RECT 1146.410 1200.400 1146.690 1200.680 ;
        RECT 1147.790 1200.400 1148.070 1200.680 ;
        RECT 1146.410 1103.840 1146.690 1104.120 ;
        RECT 1148.250 1103.840 1148.530 1104.120 ;
        RECT 1146.410 724.400 1146.690 724.680 ;
        RECT 1147.790 724.400 1148.070 724.680 ;
        RECT 1146.410 627.840 1146.690 628.120 ;
        RECT 1147.790 627.840 1148.070 628.120 ;
      LAYER met3 ;
        RECT 1146.385 1628.410 1146.715 1628.425 ;
        RECT 1147.305 1628.410 1147.635 1628.425 ;
        RECT 1146.385 1628.110 1147.635 1628.410 ;
        RECT 1146.385 1628.095 1146.715 1628.110 ;
        RECT 1147.305 1628.095 1147.635 1628.110 ;
        RECT 1146.385 1200.690 1146.715 1200.705 ;
        RECT 1147.765 1200.690 1148.095 1200.705 ;
        RECT 1146.385 1200.390 1148.095 1200.690 ;
        RECT 1146.385 1200.375 1146.715 1200.390 ;
        RECT 1147.765 1200.375 1148.095 1200.390 ;
        RECT 1146.385 1104.130 1146.715 1104.145 ;
        RECT 1148.225 1104.130 1148.555 1104.145 ;
        RECT 1146.385 1103.830 1148.555 1104.130 ;
        RECT 1146.385 1103.815 1146.715 1103.830 ;
        RECT 1148.225 1103.815 1148.555 1103.830 ;
        RECT 1146.385 724.690 1146.715 724.705 ;
        RECT 1147.765 724.690 1148.095 724.705 ;
        RECT 1146.385 724.390 1148.095 724.690 ;
        RECT 1146.385 724.375 1146.715 724.390 ;
        RECT 1147.765 724.375 1148.095 724.390 ;
        RECT 1146.385 628.130 1146.715 628.145 ;
        RECT 1147.765 628.130 1148.095 628.145 ;
        RECT 1146.385 627.830 1148.095 628.130 ;
        RECT 1146.385 627.815 1146.715 627.830 ;
        RECT 1147.765 627.815 1148.095 627.830 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 0.300 ;
=======
=======
      LAYER li1 ;
        RECT 1097.245 20.825 1097.415 24.395 ;
        RECT 1132.205 20.825 1132.375 24.395 ;
      LAYER mcon ;
        RECT 1097.245 24.225 1097.415 24.395 ;
        RECT 1132.205 24.225 1132.375 24.395 ;
>>>>>>> re-updated local openlane
      LAYER met1 ;
        RECT 14.330 24.380 14.650 24.440 ;
        RECT 1097.185 24.380 1097.475 24.425 ;
        RECT 14.330 24.240 1097.475 24.380 ;
        RECT 14.330 24.180 14.650 24.240 ;
        RECT 1097.185 24.195 1097.475 24.240 ;
        RECT 1132.145 24.380 1132.435 24.425 ;
        RECT 1152.830 24.380 1153.150 24.440 ;
        RECT 1132.145 24.240 1153.150 24.380 ;
        RECT 1132.145 24.195 1132.435 24.240 ;
        RECT 1152.830 24.180 1153.150 24.240 ;
        RECT 1097.185 20.980 1097.475 21.025 ;
        RECT 1132.145 20.980 1132.435 21.025 ;
        RECT 1097.185 20.840 1132.435 20.980 ;
        RECT 1097.185 20.795 1097.475 20.840 ;
        RECT 1132.145 20.795 1132.435 20.840 ;
      LAYER via ;
        RECT 14.360 24.180 14.620 24.440 ;
        RECT 1152.860 24.180 1153.120 24.440 ;
      LAYER met2 ;
        RECT 1153.770 1700.410 1154.050 1704.000 ;
        RECT 1152.920 1700.270 1154.050 1700.410 ;
        RECT 1152.920 24.470 1153.060 1700.270 ;
        RECT 1153.770 1700.000 1154.050 1700.270 ;
        RECT 14.360 24.150 14.620 24.470 ;
        RECT 1152.860 24.150 1153.120 24.470 ;
        RECT 14.420 2.400 14.560 24.150 ;
        RECT 14.210 -4.800 14.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 0.300 ;
=======
      LAYER met1 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 1160.190 25.060 1160.510 25.120 ;
        RECT 38.250 24.920 1160.510 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 1160.190 24.860 1160.510 24.920 ;
      LAYER via ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 1160.220 24.860 1160.480 25.120 ;
      LAYER met2 ;
        RECT 1160.210 1700.000 1160.490 1704.000 ;
        RECT 1160.280 25.150 1160.420 1700.000 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 1160.220 24.830 1160.480 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 38.130 -4.800 38.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 240.650 25.400 240.970 25.460 ;
        RECT 1215.390 25.400 1215.710 25.460 ;
        RECT 240.650 25.260 1215.710 25.400 ;
        RECT 240.650 25.200 240.970 25.260 ;
        RECT 1215.390 25.200 1215.710 25.260 ;
      LAYER via ;
        RECT 240.680 25.200 240.940 25.460 ;
        RECT 1215.420 25.200 1215.680 25.460 ;
      LAYER met2 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 240.530 -4.800 241.090 0.300 ;
=======
        RECT 1214.490 1700.000 1214.770 1704.000 ;
        RECT 1214.560 24.325 1214.700 1700.000 ;
        RECT 240.670 23.955 240.950 24.325 ;
        RECT 1214.490 23.955 1214.770 24.325 ;
        RECT 240.740 2.400 240.880 23.955 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 240.670 24.000 240.950 24.280 ;
        RECT 1214.490 24.000 1214.770 24.280 ;
      LAYER met3 ;
        RECT 240.645 24.290 240.975 24.305 ;
        RECT 1214.465 24.290 1214.795 24.305 ;
        RECT 240.645 23.990 1214.795 24.290 ;
        RECT 240.645 23.975 240.975 23.990 ;
        RECT 1214.465 23.975 1214.795 23.990 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1214.950 1700.410 1215.230 1704.000 ;
        RECT 1214.950 1700.270 1215.620 1700.410 ;
        RECT 1214.950 1700.000 1215.230 1700.270 ;
        RECT 1215.480 25.490 1215.620 1700.270 ;
        RECT 240.680 25.170 240.940 25.490 ;
        RECT 1215.420 25.170 1215.680 25.490 ;
        RECT 240.740 2.400 240.880 25.170 ;
        RECT 240.530 -4.800 241.090 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 0.300 ;
=======
      LAYER met1 ;
        RECT 1214.930 1678.140 1215.250 1678.200 ;
        RECT 1218.150 1678.140 1218.470 1678.200 ;
        RECT 1214.930 1678.000 1218.470 1678.140 ;
        RECT 1214.930 1677.940 1215.250 1678.000 ;
        RECT 1218.150 1677.940 1218.470 1678.000 ;
      LAYER via ;
        RECT 1214.960 1677.940 1215.220 1678.200 ;
        RECT 1218.180 1677.940 1218.440 1678.200 ;
=======
      LAYER li1 ;
        RECT 1216.845 745.365 1217.015 793.475 ;
        RECT 1216.845 524.365 1217.015 572.475 ;
        RECT 1216.385 469.285 1216.555 476.595 ;
      LAYER mcon ;
        RECT 1216.845 793.305 1217.015 793.475 ;
        RECT 1216.845 572.305 1217.015 572.475 ;
        RECT 1216.385 476.425 1216.555 476.595 ;
      LAYER met1 ;
        RECT 1216.310 1510.860 1216.630 1510.920 ;
        RECT 1217.230 1510.860 1217.550 1510.920 ;
        RECT 1216.310 1510.720 1217.550 1510.860 ;
        RECT 1216.310 1510.660 1216.630 1510.720 ;
        RECT 1217.230 1510.660 1217.550 1510.720 ;
        RECT 1216.770 1449.320 1217.090 1449.380 ;
        RECT 1217.230 1449.320 1217.550 1449.380 ;
        RECT 1216.770 1449.180 1217.550 1449.320 ;
        RECT 1216.770 1449.120 1217.090 1449.180 ;
        RECT 1217.230 1449.120 1217.550 1449.180 ;
        RECT 1216.770 1028.200 1217.090 1028.460 ;
        RECT 1216.860 1027.780 1217.000 1028.200 ;
        RECT 1216.770 1027.520 1217.090 1027.780 ;
        RECT 1216.310 848.880 1216.630 848.940 ;
        RECT 1216.770 848.880 1217.090 848.940 ;
        RECT 1216.310 848.740 1217.090 848.880 ;
        RECT 1216.310 848.680 1216.630 848.740 ;
        RECT 1216.770 848.680 1217.090 848.740 ;
        RECT 1216.770 793.460 1217.090 793.520 ;
        RECT 1216.575 793.320 1217.090 793.460 ;
        RECT 1216.770 793.260 1217.090 793.320 ;
        RECT 1216.785 745.520 1217.075 745.565 ;
        RECT 1217.690 745.520 1218.010 745.580 ;
        RECT 1216.785 745.380 1218.010 745.520 ;
        RECT 1216.785 745.335 1217.075 745.380 ;
        RECT 1217.690 745.320 1218.010 745.380 ;
        RECT 1216.770 704.040 1217.090 704.100 ;
        RECT 1217.690 704.040 1218.010 704.100 ;
        RECT 1216.770 703.900 1218.010 704.040 ;
        RECT 1216.770 703.840 1217.090 703.900 ;
        RECT 1217.690 703.840 1218.010 703.900 ;
        RECT 1216.310 641.620 1216.630 641.880 ;
        RECT 1216.400 641.480 1216.540 641.620 ;
        RECT 1216.770 641.480 1217.090 641.540 ;
        RECT 1216.400 641.340 1217.090 641.480 ;
        RECT 1216.770 641.280 1217.090 641.340 ;
        RECT 1216.770 572.460 1217.090 572.520 ;
        RECT 1216.575 572.320 1217.090 572.460 ;
        RECT 1216.770 572.260 1217.090 572.320 ;
        RECT 1216.770 524.520 1217.090 524.580 ;
        RECT 1216.575 524.380 1217.090 524.520 ;
        RECT 1216.770 524.320 1217.090 524.380 ;
        RECT 1216.325 476.580 1216.615 476.625 ;
        RECT 1216.770 476.580 1217.090 476.640 ;
        RECT 1216.325 476.440 1217.090 476.580 ;
        RECT 1216.325 476.395 1216.615 476.440 ;
        RECT 1216.770 476.380 1217.090 476.440 ;
        RECT 1216.310 469.440 1216.630 469.500 ;
        RECT 1216.115 469.300 1216.630 469.440 ;
        RECT 1216.310 469.240 1216.630 469.300 ;
        RECT 1216.770 338.200 1217.090 338.260 ;
        RECT 1217.230 338.200 1217.550 338.260 ;
        RECT 1216.770 338.060 1217.550 338.200 ;
        RECT 1216.770 338.000 1217.090 338.060 ;
        RECT 1217.230 338.000 1217.550 338.060 ;
        RECT 1216.310 144.740 1216.630 144.800 ;
        RECT 1216.770 144.740 1217.090 144.800 ;
        RECT 1216.310 144.600 1217.090 144.740 ;
        RECT 1216.310 144.540 1216.630 144.600 ;
        RECT 1216.770 144.540 1217.090 144.600 ;
        RECT 258.130 25.740 258.450 25.800 ;
        RECT 1216.310 25.740 1216.630 25.800 ;
        RECT 258.130 25.600 1216.630 25.740 ;
        RECT 258.130 25.540 258.450 25.600 ;
        RECT 1216.310 25.540 1216.630 25.600 ;
      LAYER via ;
        RECT 1216.340 1510.660 1216.600 1510.920 ;
        RECT 1217.260 1510.660 1217.520 1510.920 ;
        RECT 1216.800 1449.120 1217.060 1449.380 ;
        RECT 1217.260 1449.120 1217.520 1449.380 ;
        RECT 1216.800 1028.200 1217.060 1028.460 ;
        RECT 1216.800 1027.520 1217.060 1027.780 ;
        RECT 1216.340 848.680 1216.600 848.940 ;
        RECT 1216.800 848.680 1217.060 848.940 ;
        RECT 1216.800 793.260 1217.060 793.520 ;
        RECT 1217.720 745.320 1217.980 745.580 ;
        RECT 1216.800 703.840 1217.060 704.100 ;
        RECT 1217.720 703.840 1217.980 704.100 ;
        RECT 1216.340 641.620 1216.600 641.880 ;
        RECT 1216.800 641.280 1217.060 641.540 ;
        RECT 1216.800 572.260 1217.060 572.520 ;
        RECT 1216.800 524.320 1217.060 524.580 ;
        RECT 1216.800 476.380 1217.060 476.640 ;
        RECT 1216.340 469.240 1216.600 469.500 ;
        RECT 1216.800 338.000 1217.060 338.260 ;
        RECT 1217.260 338.000 1217.520 338.260 ;
        RECT 1216.340 144.540 1216.600 144.800 ;
        RECT 1216.800 144.540 1217.060 144.800 ;
        RECT 258.160 25.540 258.420 25.800 ;
        RECT 1216.340 25.540 1216.600 25.800 ;
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1219.550 1700.410 1219.830 1704.000 ;
        RECT 1219.160 1700.270 1219.830 1700.410 ;
        RECT 1219.160 1677.290 1219.300 1700.270 ;
        RECT 1219.550 1700.000 1219.830 1700.270 ;
        RECT 1216.400 1677.150 1219.300 1677.290 ;
        RECT 1216.400 1655.530 1216.540 1677.150 ;
        RECT 1216.400 1655.390 1217.000 1655.530 ;
        RECT 1216.860 1511.370 1217.000 1655.390 ;
        RECT 1216.400 1511.230 1217.000 1511.370 ;
        RECT 1216.400 1510.950 1216.540 1511.230 ;
        RECT 1216.340 1510.630 1216.600 1510.950 ;
        RECT 1217.260 1510.630 1217.520 1510.950 ;
        RECT 1217.320 1449.410 1217.460 1510.630 ;
        RECT 1216.800 1449.090 1217.060 1449.410 ;
        RECT 1217.260 1449.090 1217.520 1449.410 ;
        RECT 1216.860 1414.810 1217.000 1449.090 ;
        RECT 1216.400 1414.670 1217.000 1414.810 ;
        RECT 1216.400 1414.130 1216.540 1414.670 ;
        RECT 1216.400 1413.990 1217.000 1414.130 ;
        RECT 1216.860 1318.250 1217.000 1413.990 ;
        RECT 1216.400 1318.110 1217.000 1318.250 ;
        RECT 1216.400 1317.570 1216.540 1318.110 ;
        RECT 1216.400 1317.430 1217.000 1317.570 ;
        RECT 1216.860 1221.690 1217.000 1317.430 ;
        RECT 1216.400 1221.550 1217.000 1221.690 ;
        RECT 1216.400 1221.010 1216.540 1221.550 ;
        RECT 1216.400 1220.870 1217.000 1221.010 ;
        RECT 1216.860 1125.130 1217.000 1220.870 ;
        RECT 1216.400 1124.990 1217.000 1125.130 ;
        RECT 1216.400 1124.450 1216.540 1124.990 ;
        RECT 1216.400 1124.310 1217.000 1124.450 ;
        RECT 1216.860 1028.490 1217.000 1124.310 ;
        RECT 1216.800 1028.170 1217.060 1028.490 ;
        RECT 1216.800 1027.490 1217.060 1027.810 ;
        RECT 1216.860 976.890 1217.000 1027.490 ;
        RECT 1216.860 976.750 1217.460 976.890 ;
        RECT 1217.320 904.925 1217.460 976.750 ;
        RECT 1217.250 904.555 1217.530 904.925 ;
        RECT 1216.330 903.875 1216.610 904.245 ;
        RECT 1216.400 848.970 1216.540 903.875 ;
        RECT 1216.340 848.650 1216.600 848.970 ;
        RECT 1216.800 848.650 1217.060 848.970 ;
        RECT 1216.860 848.370 1217.000 848.650 ;
        RECT 1216.400 848.230 1217.000 848.370 ;
        RECT 1216.400 801.565 1216.540 848.230 ;
        RECT 1216.330 801.195 1216.610 801.565 ;
        RECT 1216.790 800.515 1217.070 800.885 ;
        RECT 1216.860 793.550 1217.000 800.515 ;
        RECT 1216.800 793.230 1217.060 793.550 ;
        RECT 1217.720 745.290 1217.980 745.610 ;
        RECT 1217.780 704.130 1217.920 745.290 ;
        RECT 1216.800 703.810 1217.060 704.130 ;
        RECT 1217.720 703.810 1217.980 704.130 ;
        RECT 1216.860 690.610 1217.000 703.810 ;
        RECT 1216.400 690.470 1217.000 690.610 ;
        RECT 1216.400 641.910 1216.540 690.470 ;
        RECT 1216.340 641.590 1216.600 641.910 ;
        RECT 1216.800 641.250 1217.060 641.570 ;
        RECT 1216.860 572.550 1217.000 641.250 ;
        RECT 1216.800 572.230 1217.060 572.550 ;
        RECT 1216.800 524.290 1217.060 524.610 ;
        RECT 1216.860 476.670 1217.000 524.290 ;
        RECT 1216.800 476.350 1217.060 476.670 ;
        RECT 1216.340 469.210 1216.600 469.530 ;
        RECT 1216.400 451.930 1216.540 469.210 ;
        RECT 1216.400 451.790 1217.000 451.930 ;
        RECT 1216.860 420.650 1217.000 451.790 ;
        RECT 1216.400 420.510 1217.000 420.650 ;
        RECT 1216.400 385.970 1216.540 420.510 ;
        RECT 1216.400 385.830 1217.460 385.970 ;
        RECT 1217.320 338.290 1217.460 385.830 ;
        RECT 1216.800 337.970 1217.060 338.290 ;
        RECT 1217.260 337.970 1217.520 338.290 ;
        RECT 1216.860 169.050 1217.000 337.970 ;
        RECT 1216.400 168.910 1217.000 169.050 ;
        RECT 1216.400 144.830 1216.540 168.910 ;
        RECT 1216.340 144.510 1216.600 144.830 ;
        RECT 1216.800 144.510 1217.060 144.830 ;
        RECT 1216.860 62.290 1217.000 144.510 ;
        RECT 1216.400 62.150 1217.000 62.290 ;
        RECT 1216.400 25.830 1216.540 62.150 ;
        RECT 258.160 25.510 258.420 25.830 ;
        RECT 1216.340 25.510 1216.600 25.830 ;
        RECT 258.220 2.400 258.360 25.510 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 1217.250 904.600 1217.530 904.880 ;
        RECT 1216.330 903.920 1216.610 904.200 ;
        RECT 1216.330 801.240 1216.610 801.520 ;
        RECT 1216.790 800.560 1217.070 800.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 258.125 24.970 258.455 24.985 ;
        RECT 1214.925 24.970 1215.255 24.985 ;
        RECT 258.125 24.670 1215.255 24.970 ;
        RECT 258.125 24.655 258.455 24.670 ;
        RECT 1214.925 24.655 1215.255 24.670 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1217.225 904.890 1217.555 904.905 ;
        RECT 1215.630 904.590 1217.555 904.890 ;
        RECT 1215.630 904.210 1215.930 904.590 ;
        RECT 1217.225 904.575 1217.555 904.590 ;
        RECT 1216.305 904.210 1216.635 904.225 ;
        RECT 1215.630 903.910 1216.635 904.210 ;
        RECT 1216.305 903.895 1216.635 903.910 ;
        RECT 1216.305 801.530 1216.635 801.545 ;
        RECT 1216.305 801.230 1217.770 801.530 ;
        RECT 1216.305 801.215 1216.635 801.230 ;
        RECT 1216.765 800.850 1217.095 800.865 ;
        RECT 1217.470 800.850 1217.770 801.230 ;
        RECT 1216.765 800.550 1217.770 800.850 ;
        RECT 1216.765 800.535 1217.095 800.550 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 0.300 ;
=======
      LAYER met1 ;
        RECT 1222.290 1678.140 1222.610 1678.200 ;
        RECT 1223.670 1678.140 1223.990 1678.200 ;
        RECT 1222.290 1678.000 1223.990 1678.140 ;
        RECT 1222.290 1677.940 1222.610 1678.000 ;
        RECT 1223.670 1677.940 1223.990 1678.000 ;
        RECT 276.070 26.080 276.390 26.140 ;
        RECT 1222.290 26.080 1222.610 26.140 ;
        RECT 276.070 25.940 1222.610 26.080 ;
        RECT 276.070 25.880 276.390 25.940 ;
        RECT 1222.290 25.880 1222.610 25.940 ;
      LAYER via ;
        RECT 1222.320 1677.940 1222.580 1678.200 ;
        RECT 1223.700 1677.940 1223.960 1678.200 ;
        RECT 276.100 25.880 276.360 26.140 ;
        RECT 1222.320 25.880 1222.580 26.140 ;
      LAYER met2 ;
        RECT 1224.610 1700.410 1224.890 1704.000 ;
        RECT 1223.760 1700.270 1224.890 1700.410 ;
        RECT 1223.760 1678.230 1223.900 1700.270 ;
        RECT 1224.610 1700.000 1224.890 1700.270 ;
        RECT 1222.320 1677.910 1222.580 1678.230 ;
        RECT 1223.700 1677.910 1223.960 1678.230 ;
        RECT 1222.380 26.170 1222.520 1677.910 ;
        RECT 276.100 25.850 276.360 26.170 ;
        RECT 1222.320 25.850 1222.580 26.170 ;
        RECT 276.160 2.400 276.300 25.850 ;
        RECT 275.950 -4.800 276.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 294.010 30.840 294.330 30.900 ;
        RECT 1228.730 30.840 1229.050 30.900 ;
        RECT 294.010 30.700 1229.050 30.840 ;
        RECT 294.010 30.640 294.330 30.700 ;
        RECT 1228.730 30.640 1229.050 30.700 ;
      LAYER via ;
        RECT 294.040 30.640 294.300 30.900 ;
        RECT 1228.760 30.640 1229.020 30.900 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 293.890 -4.800 294.450 0.300 ;
=======
        RECT 1229.210 1700.410 1229.490 1704.000 ;
        RECT 1228.820 1700.270 1229.490 1700.410 ;
        RECT 1228.820 30.930 1228.960 1700.270 ;
        RECT 1229.210 1700.000 1229.490 1700.270 ;
        RECT 294.040 30.610 294.300 30.930 ;
        RECT 1228.760 30.610 1229.020 30.930 ;
        RECT 294.100 2.400 294.240 30.610 ;
        RECT 293.890 -4.800 294.450 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 294.030 30.800 294.310 31.080 ;
        RECT 1229.670 30.800 1229.950 31.080 ;
      LAYER met3 ;
        RECT 294.005 31.090 294.335 31.105 ;
        RECT 1229.645 31.090 1229.975 31.105 ;
        RECT 294.005 30.790 1229.975 31.090 ;
        RECT 294.005 30.775 294.335 30.790 ;
        RECT 1229.645 30.775 1229.975 30.790 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 0.300 ;
=======
      LAYER met1 ;
        RECT 1228.730 1678.140 1229.050 1678.200 ;
        RECT 1232.870 1678.140 1233.190 1678.200 ;
        RECT 1228.730 1678.000 1233.190 1678.140 ;
        RECT 1228.730 1677.940 1229.050 1678.000 ;
        RECT 1232.870 1677.940 1233.190 1678.000 ;
      LAYER via ;
        RECT 1228.760 1677.940 1229.020 1678.200 ;
        RECT 1232.900 1677.940 1233.160 1678.200 ;
      LAYER met2 ;
        RECT 1233.810 1700.410 1234.090 1704.000 ;
        RECT 1232.960 1700.270 1234.090 1700.410 ;
        RECT 1232.960 1678.230 1233.100 1700.270 ;
        RECT 1233.810 1700.000 1234.090 1700.270 ;
        RECT 1228.760 1677.910 1229.020 1678.230 ;
        RECT 1232.900 1677.910 1233.160 1678.230 ;
        RECT 1228.820 31.805 1228.960 1677.910 ;
        RECT 311.970 31.435 312.250 31.805 ;
        RECT 1228.750 31.435 1229.030 31.805 ;
        RECT 312.040 2.400 312.180 31.435 ;
=======
      LAYER li1 ;
        RECT 1230.645 1538.925 1230.815 1587.035 ;
        RECT 1230.185 1490.645 1230.355 1522.435 ;
        RECT 1230.645 948.685 1230.815 993.395 ;
        RECT 1230.645 758.965 1230.815 807.075 ;
        RECT 1230.185 565.845 1230.355 613.275 ;
        RECT 1230.185 469.285 1230.355 476.595 ;
        RECT 1230.645 331.245 1230.815 379.355 ;
        RECT 1230.645 89.845 1230.815 137.955 ;
      LAYER mcon ;
        RECT 1230.645 1586.865 1230.815 1587.035 ;
        RECT 1230.185 1522.265 1230.355 1522.435 ;
        RECT 1230.645 993.225 1230.815 993.395 ;
        RECT 1230.645 806.905 1230.815 807.075 ;
        RECT 1230.185 613.105 1230.355 613.275 ;
        RECT 1230.185 476.425 1230.355 476.595 ;
        RECT 1230.645 379.185 1230.815 379.355 ;
        RECT 1230.645 137.785 1230.815 137.955 ;
      LAYER met1 ;
        RECT 1230.110 1628.500 1230.430 1628.560 ;
        RECT 1232.870 1628.500 1233.190 1628.560 ;
        RECT 1230.110 1628.360 1233.190 1628.500 ;
        RECT 1230.110 1628.300 1230.430 1628.360 ;
        RECT 1232.870 1628.300 1233.190 1628.360 ;
        RECT 1230.570 1587.020 1230.890 1587.080 ;
        RECT 1230.375 1586.880 1230.890 1587.020 ;
        RECT 1230.570 1586.820 1230.890 1586.880 ;
        RECT 1230.570 1539.080 1230.890 1539.140 ;
        RECT 1230.375 1538.940 1230.890 1539.080 ;
        RECT 1230.570 1538.880 1230.890 1538.940 ;
        RECT 1230.125 1522.420 1230.415 1522.465 ;
        RECT 1230.570 1522.420 1230.890 1522.480 ;
        RECT 1230.125 1522.280 1230.890 1522.420 ;
        RECT 1230.125 1522.235 1230.415 1522.280 ;
        RECT 1230.570 1522.220 1230.890 1522.280 ;
        RECT 1230.110 1490.800 1230.430 1490.860 ;
        RECT 1229.915 1490.660 1230.430 1490.800 ;
        RECT 1230.110 1490.600 1230.430 1490.660 ;
        RECT 1230.110 1462.720 1230.430 1462.980 ;
        RECT 1230.200 1462.580 1230.340 1462.720 ;
        RECT 1230.570 1462.580 1230.890 1462.640 ;
        RECT 1230.200 1462.440 1230.890 1462.580 ;
        RECT 1230.570 1462.380 1230.890 1462.440 ;
        RECT 1230.570 1401.180 1230.890 1401.440 ;
        RECT 1230.660 1400.420 1230.800 1401.180 ;
        RECT 1230.570 1400.160 1230.890 1400.420 ;
        RECT 1229.190 1338.820 1229.510 1338.880 ;
        RECT 1230.110 1338.820 1230.430 1338.880 ;
        RECT 1229.190 1338.680 1230.430 1338.820 ;
        RECT 1229.190 1338.620 1229.510 1338.680 ;
        RECT 1230.110 1338.620 1230.430 1338.680 ;
        RECT 1230.110 1249.060 1230.430 1249.120 ;
        RECT 1231.030 1249.060 1231.350 1249.120 ;
        RECT 1230.110 1248.920 1231.350 1249.060 ;
        RECT 1230.110 1248.860 1230.430 1248.920 ;
        RECT 1231.030 1248.860 1231.350 1248.920 ;
        RECT 1230.110 1076.480 1230.430 1076.740 ;
        RECT 1230.200 1076.340 1230.340 1076.480 ;
        RECT 1230.570 1076.340 1230.890 1076.400 ;
        RECT 1230.200 1076.200 1230.890 1076.340 ;
        RECT 1230.570 1076.140 1230.890 1076.200 ;
        RECT 1230.110 1000.520 1230.430 1000.580 ;
        RECT 1230.570 1000.520 1230.890 1000.580 ;
        RECT 1230.110 1000.380 1230.890 1000.520 ;
        RECT 1230.110 1000.320 1230.430 1000.380 ;
        RECT 1230.570 1000.320 1230.890 1000.380 ;
        RECT 1230.570 993.380 1230.890 993.440 ;
        RECT 1230.375 993.240 1230.890 993.380 ;
        RECT 1230.570 993.180 1230.890 993.240 ;
        RECT 1230.570 948.840 1230.890 948.900 ;
        RECT 1230.375 948.700 1230.890 948.840 ;
        RECT 1230.570 948.640 1230.890 948.700 ;
        RECT 1230.110 904.300 1230.430 904.360 ;
        RECT 1230.570 904.300 1230.890 904.360 ;
        RECT 1230.110 904.160 1230.890 904.300 ;
        RECT 1230.110 904.100 1230.430 904.160 ;
        RECT 1230.570 904.100 1230.890 904.160 ;
        RECT 1230.570 807.060 1230.890 807.120 ;
        RECT 1230.375 806.920 1230.890 807.060 ;
        RECT 1230.570 806.860 1230.890 806.920 ;
        RECT 1230.570 759.120 1230.890 759.180 ;
        RECT 1230.375 758.980 1230.890 759.120 ;
        RECT 1230.570 758.920 1230.890 758.980 ;
        RECT 1229.190 738.720 1229.510 738.780 ;
        RECT 1230.570 738.720 1230.890 738.780 ;
        RECT 1229.190 738.580 1230.890 738.720 ;
        RECT 1229.190 738.520 1229.510 738.580 ;
        RECT 1230.570 738.520 1230.890 738.580 ;
        RECT 1229.190 662.560 1229.510 662.620 ;
        RECT 1230.110 662.560 1230.430 662.620 ;
        RECT 1229.190 662.420 1230.430 662.560 ;
        RECT 1229.190 662.360 1229.510 662.420 ;
        RECT 1230.110 662.360 1230.430 662.420 ;
        RECT 1230.110 613.740 1230.430 614.000 ;
        RECT 1230.200 613.305 1230.340 613.740 ;
        RECT 1230.125 613.075 1230.415 613.305 ;
        RECT 1230.110 566.000 1230.430 566.060 ;
        RECT 1229.915 565.860 1230.430 566.000 ;
        RECT 1230.110 565.800 1230.430 565.860 ;
        RECT 1230.125 476.580 1230.415 476.625 ;
        RECT 1230.570 476.580 1230.890 476.640 ;
        RECT 1230.125 476.440 1230.890 476.580 ;
        RECT 1230.125 476.395 1230.415 476.440 ;
        RECT 1230.570 476.380 1230.890 476.440 ;
        RECT 1230.110 469.440 1230.430 469.500 ;
        RECT 1229.915 469.300 1230.430 469.440 ;
        RECT 1230.110 469.240 1230.430 469.300 ;
        RECT 1230.570 379.340 1230.890 379.400 ;
        RECT 1230.375 379.200 1230.890 379.340 ;
        RECT 1230.570 379.140 1230.890 379.200 ;
        RECT 1230.570 331.400 1230.890 331.460 ;
        RECT 1230.375 331.260 1230.890 331.400 ;
        RECT 1230.570 331.200 1230.890 331.260 ;
        RECT 1230.110 207.100 1230.430 207.360 ;
        RECT 1230.200 206.680 1230.340 207.100 ;
        RECT 1230.110 206.420 1230.430 206.680 ;
        RECT 1230.110 144.740 1230.430 144.800 ;
        RECT 1230.570 144.740 1230.890 144.800 ;
        RECT 1230.110 144.600 1230.890 144.740 ;
        RECT 1230.110 144.540 1230.430 144.600 ;
        RECT 1230.570 144.540 1230.890 144.600 ;
        RECT 1230.570 137.940 1230.890 138.000 ;
        RECT 1230.375 137.800 1230.890 137.940 ;
        RECT 1230.570 137.740 1230.890 137.800 ;
        RECT 1230.570 90.000 1230.890 90.060 ;
        RECT 1230.375 89.860 1230.890 90.000 ;
        RECT 1230.570 89.800 1230.890 89.860 ;
        RECT 311.950 31.180 312.270 31.240 ;
        RECT 1211.710 31.180 1212.030 31.240 ;
        RECT 311.950 31.040 1212.030 31.180 ;
        RECT 311.950 30.980 312.270 31.040 ;
        RECT 1211.710 30.980 1212.030 31.040 ;
      LAYER via ;
        RECT 1230.140 1628.300 1230.400 1628.560 ;
        RECT 1232.900 1628.300 1233.160 1628.560 ;
        RECT 1230.600 1586.820 1230.860 1587.080 ;
        RECT 1230.600 1538.880 1230.860 1539.140 ;
        RECT 1230.600 1522.220 1230.860 1522.480 ;
        RECT 1230.140 1490.600 1230.400 1490.860 ;
        RECT 1230.140 1462.720 1230.400 1462.980 ;
        RECT 1230.600 1462.380 1230.860 1462.640 ;
        RECT 1230.600 1401.180 1230.860 1401.440 ;
        RECT 1230.600 1400.160 1230.860 1400.420 ;
        RECT 1229.220 1338.620 1229.480 1338.880 ;
        RECT 1230.140 1338.620 1230.400 1338.880 ;
        RECT 1230.140 1248.860 1230.400 1249.120 ;
        RECT 1231.060 1248.860 1231.320 1249.120 ;
        RECT 1230.140 1076.480 1230.400 1076.740 ;
        RECT 1230.600 1076.140 1230.860 1076.400 ;
        RECT 1230.140 1000.320 1230.400 1000.580 ;
        RECT 1230.600 1000.320 1230.860 1000.580 ;
        RECT 1230.600 993.180 1230.860 993.440 ;
        RECT 1230.600 948.640 1230.860 948.900 ;
        RECT 1230.140 904.100 1230.400 904.360 ;
        RECT 1230.600 904.100 1230.860 904.360 ;
        RECT 1230.600 806.860 1230.860 807.120 ;
        RECT 1230.600 758.920 1230.860 759.180 ;
        RECT 1229.220 738.520 1229.480 738.780 ;
        RECT 1230.600 738.520 1230.860 738.780 ;
        RECT 1229.220 662.360 1229.480 662.620 ;
        RECT 1230.140 662.360 1230.400 662.620 ;
        RECT 1230.140 613.740 1230.400 614.000 ;
        RECT 1230.140 565.800 1230.400 566.060 ;
        RECT 1230.600 476.380 1230.860 476.640 ;
        RECT 1230.140 469.240 1230.400 469.500 ;
        RECT 1230.600 379.140 1230.860 379.400 ;
        RECT 1230.600 331.200 1230.860 331.460 ;
        RECT 1230.140 207.100 1230.400 207.360 ;
        RECT 1230.140 206.420 1230.400 206.680 ;
        RECT 1230.140 144.540 1230.400 144.800 ;
        RECT 1230.600 144.540 1230.860 144.800 ;
        RECT 1230.600 137.740 1230.860 138.000 ;
        RECT 1230.600 89.800 1230.860 90.060 ;
        RECT 311.980 30.980 312.240 31.240 ;
        RECT 1211.740 30.980 1212.000 31.240 ;
      LAYER met2 ;
        RECT 1234.270 1700.410 1234.550 1704.000 ;
        RECT 1232.960 1700.270 1234.550 1700.410 ;
        RECT 1232.960 1628.590 1233.100 1700.270 ;
        RECT 1234.270 1700.000 1234.550 1700.270 ;
        RECT 1230.140 1628.270 1230.400 1628.590 ;
        RECT 1232.900 1628.270 1233.160 1628.590 ;
        RECT 1230.200 1611.330 1230.340 1628.270 ;
        RECT 1230.200 1611.190 1230.800 1611.330 ;
        RECT 1230.660 1587.110 1230.800 1611.190 ;
        RECT 1230.600 1586.790 1230.860 1587.110 ;
        RECT 1230.600 1538.850 1230.860 1539.170 ;
        RECT 1230.660 1522.510 1230.800 1538.850 ;
        RECT 1230.600 1522.190 1230.860 1522.510 ;
        RECT 1230.140 1490.570 1230.400 1490.890 ;
        RECT 1230.200 1463.010 1230.340 1490.570 ;
        RECT 1230.140 1462.690 1230.400 1463.010 ;
        RECT 1230.600 1462.350 1230.860 1462.670 ;
        RECT 1230.660 1401.470 1230.800 1462.350 ;
        RECT 1230.600 1401.150 1230.860 1401.470 ;
        RECT 1230.600 1400.130 1230.860 1400.450 ;
        RECT 1230.660 1387.045 1230.800 1400.130 ;
        RECT 1229.210 1386.675 1229.490 1387.045 ;
        RECT 1230.590 1386.675 1230.870 1387.045 ;
        RECT 1229.280 1338.910 1229.420 1386.675 ;
        RECT 1229.220 1338.590 1229.480 1338.910 ;
        RECT 1230.140 1338.590 1230.400 1338.910 ;
        RECT 1230.200 1297.285 1230.340 1338.590 ;
        RECT 1230.130 1296.915 1230.410 1297.285 ;
        RECT 1231.050 1296.915 1231.330 1297.285 ;
        RECT 1231.120 1249.150 1231.260 1296.915 ;
        RECT 1230.140 1248.830 1230.400 1249.150 ;
        RECT 1231.060 1248.830 1231.320 1249.150 ;
        RECT 1230.200 1199.930 1230.340 1248.830 ;
        RECT 1230.200 1199.790 1230.800 1199.930 ;
        RECT 1230.660 1128.530 1230.800 1199.790 ;
        RECT 1230.200 1128.390 1230.800 1128.530 ;
        RECT 1230.200 1076.770 1230.340 1128.390 ;
        RECT 1230.140 1076.450 1230.400 1076.770 ;
        RECT 1230.600 1076.110 1230.860 1076.430 ;
        RECT 1230.660 1001.485 1230.800 1076.110 ;
        RECT 1230.590 1001.115 1230.870 1001.485 ;
        RECT 1230.130 1000.435 1230.410 1000.805 ;
        RECT 1230.140 1000.290 1230.400 1000.435 ;
        RECT 1230.600 1000.290 1230.860 1000.610 ;
        RECT 1230.660 993.470 1230.800 1000.290 ;
        RECT 1230.600 993.150 1230.860 993.470 ;
        RECT 1230.600 948.610 1230.860 948.930 ;
        RECT 1230.660 904.390 1230.800 948.610 ;
        RECT 1230.140 904.070 1230.400 904.390 ;
        RECT 1230.600 904.070 1230.860 904.390 ;
        RECT 1230.200 831.370 1230.340 904.070 ;
        RECT 1230.200 831.230 1231.260 831.370 ;
        RECT 1231.120 820.490 1231.260 831.230 ;
        RECT 1230.660 820.350 1231.260 820.490 ;
        RECT 1230.660 807.150 1230.800 820.350 ;
        RECT 1230.600 806.830 1230.860 807.150 ;
        RECT 1230.600 758.890 1230.860 759.210 ;
        RECT 1230.660 738.810 1230.800 758.890 ;
        RECT 1229.220 738.490 1229.480 738.810 ;
        RECT 1230.600 738.490 1230.860 738.810 ;
        RECT 1229.280 662.650 1229.420 738.490 ;
        RECT 1229.220 662.330 1229.480 662.650 ;
        RECT 1230.140 662.330 1230.400 662.650 ;
        RECT 1230.200 614.030 1230.340 662.330 ;
        RECT 1230.140 613.710 1230.400 614.030 ;
        RECT 1230.140 565.770 1230.400 566.090 ;
        RECT 1230.200 548.490 1230.340 565.770 ;
        RECT 1230.200 548.350 1230.800 548.490 ;
        RECT 1230.660 476.670 1230.800 548.350 ;
        RECT 1230.600 476.350 1230.860 476.670 ;
        RECT 1230.140 469.210 1230.400 469.530 ;
        RECT 1230.200 451.930 1230.340 469.210 ;
        RECT 1230.200 451.790 1230.800 451.930 ;
        RECT 1230.660 379.430 1230.800 451.790 ;
        RECT 1230.600 379.110 1230.860 379.430 ;
        RECT 1230.600 331.170 1230.860 331.490 ;
        RECT 1230.660 282.610 1230.800 331.170 ;
        RECT 1230.200 282.470 1230.800 282.610 ;
        RECT 1230.200 207.390 1230.340 282.470 ;
        RECT 1230.140 207.070 1230.400 207.390 ;
        RECT 1230.140 206.390 1230.400 206.710 ;
        RECT 1230.200 144.830 1230.340 206.390 ;
        RECT 1230.140 144.510 1230.400 144.830 ;
        RECT 1230.600 144.510 1230.860 144.830 ;
        RECT 1230.660 138.030 1230.800 144.510 ;
        RECT 1230.600 137.710 1230.860 138.030 ;
        RECT 1230.600 89.770 1230.860 90.090 ;
        RECT 1230.660 49.485 1230.800 89.770 ;
        RECT 1230.590 49.115 1230.870 49.485 ;
        RECT 1211.730 47.075 1212.010 47.445 ;
        RECT 1211.800 31.270 1211.940 47.075 ;
        RECT 311.980 30.950 312.240 31.270 ;
        RECT 1211.740 30.950 1212.000 31.270 ;
        RECT 312.040 2.400 312.180 30.950 ;
>>>>>>> re-updated local openlane
        RECT 311.830 -4.800 312.390 2.400 ;
      LAYER via2 ;
        RECT 1229.210 1386.720 1229.490 1387.000 ;
        RECT 1230.590 1386.720 1230.870 1387.000 ;
        RECT 1230.130 1296.960 1230.410 1297.240 ;
        RECT 1231.050 1296.960 1231.330 1297.240 ;
        RECT 1230.590 1001.160 1230.870 1001.440 ;
        RECT 1230.130 1000.480 1230.410 1000.760 ;
        RECT 1230.590 49.160 1230.870 49.440 ;
        RECT 1211.730 47.120 1212.010 47.400 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 311.945 31.770 312.275 31.785 ;
        RECT 1228.725 31.770 1229.055 31.785 ;
        RECT 311.945 31.470 1229.055 31.770 ;
        RECT 311.945 31.455 312.275 31.470 ;
        RECT 1228.725 31.455 1229.055 31.470 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1229.185 1387.010 1229.515 1387.025 ;
        RECT 1230.565 1387.010 1230.895 1387.025 ;
        RECT 1229.185 1386.710 1230.895 1387.010 ;
        RECT 1229.185 1386.695 1229.515 1386.710 ;
        RECT 1230.565 1386.695 1230.895 1386.710 ;
        RECT 1230.105 1297.250 1230.435 1297.265 ;
        RECT 1231.025 1297.250 1231.355 1297.265 ;
        RECT 1230.105 1296.950 1231.355 1297.250 ;
        RECT 1230.105 1296.935 1230.435 1296.950 ;
        RECT 1231.025 1296.935 1231.355 1296.950 ;
        RECT 1230.565 1001.450 1230.895 1001.465 ;
        RECT 1230.350 1001.135 1230.895 1001.450 ;
        RECT 1230.350 1000.785 1230.650 1001.135 ;
        RECT 1230.105 1000.470 1230.650 1000.785 ;
        RECT 1230.105 1000.455 1230.435 1000.470 ;
        RECT 1230.565 49.450 1230.895 49.465 ;
        RECT 1230.350 49.135 1230.895 49.450 ;
        RECT 1211.705 47.410 1212.035 47.425 ;
        RECT 1230.350 47.410 1230.650 49.135 ;
        RECT 1211.705 47.110 1230.650 47.410 ;
        RECT 1211.705 47.095 1212.035 47.110 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 329.770 -4.800 330.330 0.300 ;
=======
        RECT 1238.870 1700.410 1239.150 1704.000 ;
        RECT 1238.020 1700.270 1239.150 1700.410 ;
        RECT 1238.020 1678.650 1238.160 1700.270 ;
        RECT 1238.870 1700.000 1239.150 1700.270 ;
        RECT 1236.640 1678.510 1238.160 1678.650 ;
        RECT 1236.640 32.485 1236.780 1678.510 ;
        RECT 329.910 32.115 330.190 32.485 ;
        RECT 1236.570 32.115 1236.850 32.485 ;
        RECT 329.980 2.400 330.120 32.115 ;
=======
      LAYER li1 ;
        RECT 1237.085 1496.765 1237.255 1535.015 ;
        RECT 1237.085 565.845 1237.255 613.275 ;
        RECT 1237.545 469.285 1237.715 517.395 ;
        RECT 1237.545 427.805 1237.715 435.115 ;
        RECT 1236.625 186.405 1236.795 234.515 ;
      LAYER mcon ;
        RECT 1237.085 1534.845 1237.255 1535.015 ;
        RECT 1237.085 613.105 1237.255 613.275 ;
        RECT 1237.545 517.225 1237.715 517.395 ;
        RECT 1237.545 434.945 1237.715 435.115 ;
        RECT 1236.625 234.345 1236.795 234.515 ;
      LAYER met1 ;
        RECT 1237.930 1684.260 1238.250 1684.320 ;
        RECT 1238.850 1684.260 1239.170 1684.320 ;
        RECT 1237.930 1684.120 1239.170 1684.260 ;
        RECT 1237.930 1684.060 1238.250 1684.120 ;
        RECT 1238.850 1684.060 1239.170 1684.120 ;
        RECT 1237.930 1676.440 1238.250 1676.500 ;
        RECT 1238.390 1676.440 1238.710 1676.500 ;
        RECT 1237.930 1676.300 1238.710 1676.440 ;
        RECT 1237.930 1676.240 1238.250 1676.300 ;
        RECT 1238.390 1676.240 1238.710 1676.300 ;
        RECT 1237.025 1535.000 1237.315 1535.045 ;
        RECT 1238.390 1535.000 1238.710 1535.060 ;
        RECT 1237.025 1534.860 1238.710 1535.000 ;
        RECT 1237.025 1534.815 1237.315 1534.860 ;
        RECT 1238.390 1534.800 1238.710 1534.860 ;
        RECT 1237.025 1496.920 1237.315 1496.965 ;
        RECT 1237.470 1496.920 1237.790 1496.980 ;
        RECT 1237.025 1496.780 1237.790 1496.920 ;
        RECT 1237.025 1496.735 1237.315 1496.780 ;
        RECT 1237.470 1496.720 1237.790 1496.780 ;
        RECT 1236.550 1435.380 1236.870 1435.440 ;
        RECT 1238.390 1435.380 1238.710 1435.440 ;
        RECT 1236.550 1435.240 1238.710 1435.380 ;
        RECT 1236.550 1435.180 1236.870 1435.240 ;
        RECT 1238.390 1435.180 1238.710 1435.240 ;
        RECT 1236.550 1338.820 1236.870 1338.880 ;
        RECT 1237.010 1338.820 1237.330 1338.880 ;
        RECT 1236.550 1338.680 1237.330 1338.820 ;
        RECT 1236.550 1338.620 1236.870 1338.680 ;
        RECT 1237.010 1338.620 1237.330 1338.680 ;
        RECT 1236.550 1269.600 1236.870 1269.860 ;
        RECT 1236.640 1269.120 1236.780 1269.600 ;
        RECT 1237.010 1269.120 1237.330 1269.180 ;
        RECT 1236.640 1268.980 1237.330 1269.120 ;
        RECT 1237.010 1268.920 1237.330 1268.980 ;
        RECT 1237.010 1207.920 1237.330 1207.980 ;
        RECT 1236.640 1207.780 1237.330 1207.920 ;
        RECT 1236.640 1207.640 1236.780 1207.780 ;
        RECT 1237.010 1207.720 1237.330 1207.780 ;
        RECT 1236.550 1207.380 1236.870 1207.640 ;
        RECT 1235.630 1151.820 1235.950 1151.880 ;
        RECT 1237.470 1151.820 1237.790 1151.880 ;
        RECT 1235.630 1151.680 1237.790 1151.820 ;
        RECT 1235.630 1151.620 1235.950 1151.680 ;
        RECT 1237.470 1151.620 1237.790 1151.680 ;
        RECT 1237.470 1145.360 1237.790 1145.420 ;
        RECT 1238.390 1145.360 1238.710 1145.420 ;
        RECT 1237.470 1145.220 1238.710 1145.360 ;
        RECT 1237.470 1145.160 1237.790 1145.220 ;
        RECT 1238.390 1145.160 1238.710 1145.220 ;
        RECT 1236.550 855.340 1236.870 855.400 ;
        RECT 1237.010 855.340 1237.330 855.400 ;
        RECT 1236.550 855.200 1237.330 855.340 ;
        RECT 1236.550 855.140 1236.870 855.200 ;
        RECT 1237.010 855.140 1237.330 855.200 ;
        RECT 1237.010 613.740 1237.330 614.000 ;
        RECT 1237.100 613.305 1237.240 613.740 ;
        RECT 1237.025 613.075 1237.315 613.305 ;
        RECT 1237.010 566.000 1237.330 566.060 ;
        RECT 1236.815 565.860 1237.330 566.000 ;
        RECT 1237.010 565.800 1237.330 565.860 ;
        RECT 1237.470 517.380 1237.790 517.440 ;
        RECT 1237.275 517.240 1237.790 517.380 ;
        RECT 1237.470 517.180 1237.790 517.240 ;
        RECT 1237.470 469.440 1237.790 469.500 ;
        RECT 1237.275 469.300 1237.790 469.440 ;
        RECT 1237.470 469.240 1237.790 469.300 ;
        RECT 1237.470 435.100 1237.790 435.160 ;
        RECT 1237.275 434.960 1237.790 435.100 ;
        RECT 1237.470 434.900 1237.790 434.960 ;
        RECT 1237.470 427.960 1237.790 428.020 ;
        RECT 1237.275 427.820 1237.790 427.960 ;
        RECT 1237.470 427.760 1237.790 427.820 ;
        RECT 1236.550 379.340 1236.870 379.400 ;
        RECT 1237.470 379.340 1237.790 379.400 ;
        RECT 1236.550 379.200 1237.790 379.340 ;
        RECT 1236.550 379.140 1236.870 379.200 ;
        RECT 1237.470 379.140 1237.790 379.200 ;
        RECT 1236.550 241.640 1236.870 241.700 ;
        RECT 1237.930 241.640 1238.250 241.700 ;
        RECT 1236.550 241.500 1238.250 241.640 ;
        RECT 1236.550 241.440 1236.870 241.500 ;
        RECT 1237.930 241.440 1238.250 241.500 ;
        RECT 1236.550 234.500 1236.870 234.560 ;
        RECT 1236.355 234.360 1236.870 234.500 ;
        RECT 1236.550 234.300 1236.870 234.360 ;
        RECT 1236.550 186.560 1236.870 186.620 ;
        RECT 1236.355 186.420 1236.870 186.560 ;
        RECT 1236.550 186.360 1236.870 186.420 ;
        RECT 1236.550 137.940 1236.870 138.000 ;
        RECT 1237.010 137.940 1237.330 138.000 ;
        RECT 1236.550 137.800 1237.330 137.940 ;
        RECT 1236.550 137.740 1236.870 137.800 ;
        RECT 1237.010 137.740 1237.330 137.800 ;
        RECT 329.890 31.520 330.210 31.580 ;
        RECT 1237.010 31.520 1237.330 31.580 ;
        RECT 329.890 31.380 1237.330 31.520 ;
        RECT 329.890 31.320 330.210 31.380 ;
        RECT 1237.010 31.320 1237.330 31.380 ;
      LAYER via ;
        RECT 1237.960 1684.060 1238.220 1684.320 ;
        RECT 1238.880 1684.060 1239.140 1684.320 ;
        RECT 1237.960 1676.240 1238.220 1676.500 ;
        RECT 1238.420 1676.240 1238.680 1676.500 ;
        RECT 1238.420 1534.800 1238.680 1535.060 ;
        RECT 1237.500 1496.720 1237.760 1496.980 ;
        RECT 1236.580 1435.180 1236.840 1435.440 ;
        RECT 1238.420 1435.180 1238.680 1435.440 ;
        RECT 1236.580 1338.620 1236.840 1338.880 ;
        RECT 1237.040 1338.620 1237.300 1338.880 ;
        RECT 1236.580 1269.600 1236.840 1269.860 ;
        RECT 1237.040 1268.920 1237.300 1269.180 ;
        RECT 1237.040 1207.720 1237.300 1207.980 ;
        RECT 1236.580 1207.380 1236.840 1207.640 ;
        RECT 1235.660 1151.620 1235.920 1151.880 ;
        RECT 1237.500 1151.620 1237.760 1151.880 ;
        RECT 1237.500 1145.160 1237.760 1145.420 ;
        RECT 1238.420 1145.160 1238.680 1145.420 ;
        RECT 1236.580 855.140 1236.840 855.400 ;
        RECT 1237.040 855.140 1237.300 855.400 ;
        RECT 1237.040 613.740 1237.300 614.000 ;
        RECT 1237.040 565.800 1237.300 566.060 ;
        RECT 1237.500 517.180 1237.760 517.440 ;
        RECT 1237.500 469.240 1237.760 469.500 ;
        RECT 1237.500 434.900 1237.760 435.160 ;
        RECT 1237.500 427.760 1237.760 428.020 ;
        RECT 1236.580 379.140 1236.840 379.400 ;
        RECT 1237.500 379.140 1237.760 379.400 ;
        RECT 1236.580 241.440 1236.840 241.700 ;
        RECT 1237.960 241.440 1238.220 241.700 ;
        RECT 1236.580 234.300 1236.840 234.560 ;
        RECT 1236.580 186.360 1236.840 186.620 ;
        RECT 1236.580 137.740 1236.840 138.000 ;
        RECT 1237.040 137.740 1237.300 138.000 ;
        RECT 329.920 31.320 330.180 31.580 ;
        RECT 1237.040 31.320 1237.300 31.580 ;
      LAYER met2 ;
        RECT 1238.870 1700.000 1239.150 1704.000 ;
        RECT 1238.940 1684.350 1239.080 1700.000 ;
        RECT 1237.960 1684.030 1238.220 1684.350 ;
        RECT 1238.880 1684.030 1239.140 1684.350 ;
        RECT 1238.020 1676.530 1238.160 1684.030 ;
        RECT 1237.960 1676.210 1238.220 1676.530 ;
        RECT 1238.420 1676.210 1238.680 1676.530 ;
        RECT 1238.480 1535.090 1238.620 1676.210 ;
        RECT 1238.420 1534.770 1238.680 1535.090 ;
        RECT 1237.500 1496.690 1237.760 1497.010 ;
        RECT 1237.560 1483.605 1237.700 1496.690 ;
        RECT 1237.490 1483.235 1237.770 1483.605 ;
        RECT 1238.410 1483.235 1238.690 1483.605 ;
        RECT 1238.480 1435.470 1238.620 1483.235 ;
        RECT 1236.580 1435.150 1236.840 1435.470 ;
        RECT 1238.420 1435.150 1238.680 1435.470 ;
        RECT 1236.640 1386.930 1236.780 1435.150 ;
        RECT 1236.640 1386.790 1237.240 1386.930 ;
        RECT 1237.100 1338.910 1237.240 1386.790 ;
        RECT 1236.580 1338.590 1236.840 1338.910 ;
        RECT 1237.040 1338.590 1237.300 1338.910 ;
        RECT 1236.640 1269.890 1236.780 1338.590 ;
        RECT 1236.580 1269.570 1236.840 1269.890 ;
        RECT 1237.040 1268.890 1237.300 1269.210 ;
        RECT 1237.100 1208.010 1237.240 1268.890 ;
        RECT 1237.040 1207.690 1237.300 1208.010 ;
        RECT 1236.580 1207.350 1236.840 1207.670 ;
        RECT 1236.640 1200.725 1236.780 1207.350 ;
        RECT 1235.650 1200.355 1235.930 1200.725 ;
        RECT 1236.570 1200.355 1236.850 1200.725 ;
        RECT 1235.720 1151.910 1235.860 1200.355 ;
        RECT 1235.660 1151.590 1235.920 1151.910 ;
        RECT 1237.500 1151.590 1237.760 1151.910 ;
        RECT 1237.560 1145.450 1237.700 1151.590 ;
        RECT 1237.500 1145.130 1237.760 1145.450 ;
        RECT 1238.420 1145.130 1238.680 1145.450 ;
        RECT 1238.480 1097.365 1238.620 1145.130 ;
        RECT 1237.030 1096.995 1237.310 1097.365 ;
        RECT 1238.410 1096.995 1238.690 1097.365 ;
        RECT 1237.100 855.430 1237.240 1096.995 ;
        RECT 1236.580 855.110 1236.840 855.430 ;
        RECT 1237.040 855.110 1237.300 855.430 ;
        RECT 1236.640 783.090 1236.780 855.110 ;
        RECT 1236.640 782.950 1237.240 783.090 ;
        RECT 1237.100 614.030 1237.240 782.950 ;
        RECT 1237.040 613.710 1237.300 614.030 ;
        RECT 1237.040 565.770 1237.300 566.090 ;
        RECT 1237.100 565.605 1237.240 565.770 ;
        RECT 1237.030 565.235 1237.310 565.605 ;
        RECT 1237.490 517.635 1237.770 518.005 ;
        RECT 1237.560 517.470 1237.700 517.635 ;
        RECT 1237.500 517.150 1237.760 517.470 ;
        RECT 1237.500 469.210 1237.760 469.530 ;
        RECT 1237.560 435.190 1237.700 469.210 ;
        RECT 1237.500 434.870 1237.760 435.190 ;
        RECT 1237.500 427.730 1237.760 428.050 ;
        RECT 1237.560 379.430 1237.700 427.730 ;
        RECT 1236.580 379.110 1236.840 379.430 ;
        RECT 1237.500 379.110 1237.760 379.430 ;
        RECT 1236.640 307.090 1236.780 379.110 ;
        RECT 1236.640 306.950 1237.700 307.090 ;
        RECT 1237.560 288.730 1237.700 306.950 ;
        RECT 1237.560 288.590 1238.160 288.730 ;
        RECT 1238.020 241.730 1238.160 288.590 ;
        RECT 1236.580 241.410 1236.840 241.730 ;
        RECT 1237.960 241.410 1238.220 241.730 ;
        RECT 1236.640 234.590 1236.780 241.410 ;
        RECT 1236.580 234.270 1236.840 234.590 ;
        RECT 1236.580 186.330 1236.840 186.650 ;
        RECT 1236.640 138.030 1236.780 186.330 ;
        RECT 1236.580 137.710 1236.840 138.030 ;
        RECT 1237.040 137.710 1237.300 138.030 ;
        RECT 1237.100 31.610 1237.240 137.710 ;
        RECT 329.920 31.290 330.180 31.610 ;
        RECT 1237.040 31.290 1237.300 31.610 ;
        RECT 329.980 2.400 330.120 31.290 ;
>>>>>>> re-updated local openlane
        RECT 329.770 -4.800 330.330 2.400 ;
      LAYER via2 ;
        RECT 1237.490 1483.280 1237.770 1483.560 ;
        RECT 1238.410 1483.280 1238.690 1483.560 ;
        RECT 1235.650 1200.400 1235.930 1200.680 ;
        RECT 1236.570 1200.400 1236.850 1200.680 ;
        RECT 1237.030 1097.040 1237.310 1097.320 ;
        RECT 1238.410 1097.040 1238.690 1097.320 ;
        RECT 1237.030 565.280 1237.310 565.560 ;
        RECT 1237.490 517.680 1237.770 517.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 329.885 32.450 330.215 32.465 ;
        RECT 1236.545 32.450 1236.875 32.465 ;
        RECT 329.885 32.150 1236.875 32.450 ;
        RECT 329.885 32.135 330.215 32.150 ;
        RECT 1236.545 32.135 1236.875 32.150 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1237.465 1483.570 1237.795 1483.585 ;
        RECT 1238.385 1483.570 1238.715 1483.585 ;
        RECT 1237.465 1483.270 1238.715 1483.570 ;
        RECT 1237.465 1483.255 1237.795 1483.270 ;
        RECT 1238.385 1483.255 1238.715 1483.270 ;
        RECT 1235.625 1200.690 1235.955 1200.705 ;
        RECT 1236.545 1200.690 1236.875 1200.705 ;
        RECT 1235.625 1200.390 1236.875 1200.690 ;
        RECT 1235.625 1200.375 1235.955 1200.390 ;
        RECT 1236.545 1200.375 1236.875 1200.390 ;
        RECT 1237.005 1097.330 1237.335 1097.345 ;
        RECT 1238.385 1097.330 1238.715 1097.345 ;
        RECT 1237.005 1097.030 1238.715 1097.330 ;
        RECT 1237.005 1097.015 1237.335 1097.030 ;
        RECT 1238.385 1097.015 1238.715 1097.030 ;
        RECT 1237.005 565.570 1237.335 565.585 ;
        RECT 1237.005 565.270 1238.010 565.570 ;
        RECT 1237.005 565.255 1237.335 565.270 ;
        RECT 1236.750 564.890 1237.130 564.900 ;
        RECT 1237.710 564.890 1238.010 565.270 ;
        RECT 1236.750 564.590 1238.010 564.890 ;
        RECT 1236.750 564.580 1237.130 564.590 ;
        RECT 1236.750 517.970 1237.130 517.980 ;
        RECT 1237.465 517.970 1237.795 517.985 ;
        RECT 1236.750 517.670 1237.795 517.970 ;
        RECT 1236.750 517.660 1237.130 517.670 ;
        RECT 1237.465 517.655 1237.795 517.670 ;
      LAYER via3 ;
        RECT 1236.780 564.580 1237.100 564.900 ;
        RECT 1236.780 517.660 1237.100 517.980 ;
      LAYER met4 ;
        RECT 1236.775 564.575 1237.105 564.905 ;
        RECT 1236.790 517.985 1237.090 564.575 ;
        RECT 1236.775 517.655 1237.105 517.985 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 0.300 ;
=======
      LAYER met1 ;
        RECT 347.370 39.680 347.690 39.740 ;
        RECT 1242.990 39.680 1243.310 39.740 ;
        RECT 347.370 39.540 1243.310 39.680 ;
        RECT 347.370 39.480 347.690 39.540 ;
        RECT 1242.990 39.480 1243.310 39.540 ;
      LAYER via ;
        RECT 347.400 39.480 347.660 39.740 ;
        RECT 1243.020 39.480 1243.280 39.740 ;
      LAYER met2 ;
        RECT 1243.930 1700.410 1244.210 1704.000 ;
        RECT 1243.080 1700.270 1244.210 1700.410 ;
        RECT 1243.080 39.770 1243.220 1700.270 ;
        RECT 1243.930 1700.000 1244.210 1700.270 ;
        RECT 347.400 39.450 347.660 39.770 ;
        RECT 1243.020 39.450 1243.280 39.770 ;
        RECT 347.460 2.400 347.600 39.450 ;
        RECT 347.250 -4.800 347.810 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 0.300 ;
=======
      LAYER met1 ;
        RECT 1243.450 1664.880 1243.770 1664.940 ;
        RECT 1247.590 1664.880 1247.910 1664.940 ;
        RECT 1243.450 1664.740 1247.910 1664.880 ;
        RECT 1243.450 1664.680 1243.770 1664.740 ;
        RECT 1247.590 1664.680 1247.910 1664.740 ;
        RECT 365.310 40.020 365.630 40.080 ;
        RECT 1243.450 40.020 1243.770 40.080 ;
        RECT 365.310 39.880 1243.770 40.020 ;
        RECT 365.310 39.820 365.630 39.880 ;
        RECT 1243.450 39.820 1243.770 39.880 ;
      LAYER via ;
        RECT 1243.480 1664.680 1243.740 1664.940 ;
        RECT 1247.620 1664.680 1247.880 1664.940 ;
        RECT 365.340 39.820 365.600 40.080 ;
        RECT 1243.480 39.820 1243.740 40.080 ;
      LAYER met2 ;
        RECT 1248.530 1700.410 1248.810 1704.000 ;
        RECT 1247.680 1700.270 1248.810 1700.410 ;
        RECT 1247.680 1664.970 1247.820 1700.270 ;
        RECT 1248.530 1700.000 1248.810 1700.270 ;
        RECT 1243.480 1664.650 1243.740 1664.970 ;
        RECT 1247.620 1664.650 1247.880 1664.970 ;
        RECT 1243.540 40.110 1243.680 1664.650 ;
        RECT 365.340 39.790 365.600 40.110 ;
        RECT 1243.480 39.790 1243.740 40.110 ;
        RECT 365.400 2.400 365.540 39.790 ;
        RECT 365.190 -4.800 365.750 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 0.300 ;
=======
      LAYER met1 ;
        RECT 1249.430 1677.800 1249.750 1677.860 ;
        RECT 1252.190 1677.800 1252.510 1677.860 ;
        RECT 1249.430 1677.660 1252.510 1677.800 ;
        RECT 1249.430 1677.600 1249.750 1677.660 ;
        RECT 1252.190 1677.600 1252.510 1677.660 ;
        RECT 383.250 40.360 383.570 40.420 ;
        RECT 1249.430 40.360 1249.750 40.420 ;
        RECT 383.250 40.220 1249.750 40.360 ;
        RECT 383.250 40.160 383.570 40.220 ;
        RECT 1249.430 40.160 1249.750 40.220 ;
      LAYER via ;
        RECT 1249.460 1677.600 1249.720 1677.860 ;
        RECT 1252.220 1677.600 1252.480 1677.860 ;
        RECT 383.280 40.160 383.540 40.420 ;
        RECT 1249.460 40.160 1249.720 40.420 ;
      LAYER met2 ;
        RECT 1253.590 1700.410 1253.870 1704.000 ;
        RECT 1252.280 1700.270 1253.870 1700.410 ;
        RECT 1252.280 1677.890 1252.420 1700.270 ;
        RECT 1253.590 1700.000 1253.870 1700.270 ;
        RECT 1249.460 1677.570 1249.720 1677.890 ;
        RECT 1252.220 1677.570 1252.480 1677.890 ;
        RECT 1249.520 40.450 1249.660 1677.570 ;
        RECT 383.280 40.130 383.540 40.450 ;
        RECT 1249.460 40.130 1249.720 40.450 ;
        RECT 383.340 2.400 383.480 40.130 ;
        RECT 383.130 -4.800 383.690 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 0.300 ;
=======
      LAYER li1 ;
        RECT 1258.245 1635.485 1258.415 1683.595 ;
        RECT 1257.785 1497.785 1257.955 1563.235 ;
        RECT 1257.785 1048.985 1257.955 1103.895 ;
        RECT 1258.245 421.345 1258.415 510.595 ;
        RECT 1258.245 228.225 1258.415 275.995 ;
        RECT 1257.785 89.845 1257.955 137.955 ;
      LAYER mcon ;
        RECT 1258.245 1683.425 1258.415 1683.595 ;
        RECT 1257.785 1563.065 1257.955 1563.235 ;
        RECT 1257.785 1103.725 1257.955 1103.895 ;
        RECT 1258.245 510.425 1258.415 510.595 ;
        RECT 1258.245 275.825 1258.415 275.995 ;
        RECT 1257.785 137.785 1257.955 137.955 ;
      LAYER met1 ;
        RECT 1258.170 1683.580 1258.490 1683.640 ;
        RECT 1257.975 1683.440 1258.490 1683.580 ;
        RECT 1258.170 1683.380 1258.490 1683.440 ;
        RECT 1258.170 1635.640 1258.490 1635.700 ;
        RECT 1257.975 1635.500 1258.490 1635.640 ;
        RECT 1258.170 1635.440 1258.490 1635.500 ;
        RECT 1257.250 1563.220 1257.570 1563.280 ;
        RECT 1257.725 1563.220 1258.015 1563.265 ;
        RECT 1257.250 1563.080 1258.015 1563.220 ;
        RECT 1257.250 1563.020 1257.570 1563.080 ;
        RECT 1257.725 1563.035 1258.015 1563.080 ;
        RECT 1257.710 1497.940 1258.030 1498.000 ;
        RECT 1257.515 1497.800 1258.030 1497.940 ;
        RECT 1257.710 1497.740 1258.030 1497.800 ;
        RECT 1257.710 1448.640 1258.030 1448.700 ;
        RECT 1259.090 1448.640 1259.410 1448.700 ;
        RECT 1257.710 1448.500 1259.410 1448.640 ;
        RECT 1257.710 1448.440 1258.030 1448.500 ;
        RECT 1259.090 1448.440 1259.410 1448.500 ;
        RECT 1257.250 1352.760 1257.570 1352.820 ;
        RECT 1258.170 1352.760 1258.490 1352.820 ;
        RECT 1257.250 1352.620 1258.490 1352.760 ;
        RECT 1257.250 1352.560 1257.570 1352.620 ;
        RECT 1258.170 1352.560 1258.490 1352.620 ;
        RECT 1258.170 1221.860 1258.490 1221.920 ;
        RECT 1257.800 1221.720 1258.490 1221.860 ;
        RECT 1257.800 1221.240 1257.940 1221.720 ;
        RECT 1258.170 1221.660 1258.490 1221.720 ;
        RECT 1257.710 1220.980 1258.030 1221.240 ;
        RECT 1257.710 1103.880 1258.030 1103.940 ;
        RECT 1257.515 1103.740 1258.030 1103.880 ;
        RECT 1257.710 1103.680 1258.030 1103.740 ;
        RECT 1257.710 1049.140 1258.030 1049.200 ;
        RECT 1257.515 1049.000 1258.030 1049.140 ;
        RECT 1257.710 1048.940 1258.030 1049.000 ;
        RECT 1257.710 1007.320 1258.030 1007.380 ;
        RECT 1258.630 1007.320 1258.950 1007.380 ;
        RECT 1257.710 1007.180 1258.950 1007.320 ;
        RECT 1257.710 1007.120 1258.030 1007.180 ;
        RECT 1258.630 1007.120 1258.950 1007.180 ;
        RECT 1258.170 869.620 1258.490 869.680 ;
        RECT 1258.630 869.620 1258.950 869.680 ;
        RECT 1258.170 869.480 1258.950 869.620 ;
        RECT 1258.170 869.420 1258.490 869.480 ;
        RECT 1258.630 869.420 1258.950 869.480 ;
        RECT 1257.710 710.840 1258.030 710.900 ;
        RECT 1258.170 710.840 1258.490 710.900 ;
        RECT 1257.710 710.700 1258.490 710.840 ;
        RECT 1257.710 710.640 1258.030 710.700 ;
        RECT 1258.170 710.640 1258.490 710.700 ;
        RECT 1256.790 652.020 1257.110 652.080 ;
        RECT 1257.710 652.020 1258.030 652.080 ;
        RECT 1256.790 651.880 1258.030 652.020 ;
        RECT 1256.790 651.820 1257.110 651.880 ;
        RECT 1257.710 651.820 1258.030 651.880 ;
        RECT 1257.710 510.580 1258.030 510.640 ;
        RECT 1258.185 510.580 1258.475 510.625 ;
        RECT 1257.710 510.440 1258.475 510.580 ;
        RECT 1257.710 510.380 1258.030 510.440 ;
        RECT 1258.185 510.395 1258.475 510.440 ;
        RECT 1258.185 421.500 1258.475 421.545 ;
        RECT 1257.800 421.360 1258.475 421.500 ;
        RECT 1257.800 420.820 1257.940 421.360 ;
        RECT 1258.185 421.315 1258.475 421.360 ;
        RECT 1258.170 420.820 1258.490 420.880 ;
        RECT 1257.800 420.680 1258.490 420.820 ;
        RECT 1258.170 420.620 1258.490 420.680 ;
        RECT 1257.710 283.120 1258.030 283.180 ;
        RECT 1259.090 283.120 1259.410 283.180 ;
        RECT 1257.710 282.980 1259.410 283.120 ;
        RECT 1257.710 282.920 1258.030 282.980 ;
        RECT 1259.090 282.920 1259.410 282.980 ;
        RECT 1258.185 275.980 1258.475 276.025 ;
        RECT 1259.090 275.980 1259.410 276.040 ;
        RECT 1258.185 275.840 1259.410 275.980 ;
        RECT 1258.185 275.795 1258.475 275.840 ;
        RECT 1259.090 275.780 1259.410 275.840 ;
        RECT 1258.170 228.380 1258.490 228.440 ;
        RECT 1257.975 228.240 1258.490 228.380 ;
        RECT 1258.170 228.180 1258.490 228.240 ;
        RECT 1257.710 227.700 1258.030 227.760 ;
        RECT 1258.170 227.700 1258.490 227.760 ;
        RECT 1257.710 227.560 1258.490 227.700 ;
        RECT 1257.710 227.500 1258.030 227.560 ;
        RECT 1258.170 227.500 1258.490 227.560 ;
        RECT 1257.710 145.420 1258.030 145.480 ;
        RECT 1258.170 145.420 1258.490 145.480 ;
        RECT 1257.710 145.280 1258.490 145.420 ;
        RECT 1257.710 145.220 1258.030 145.280 ;
        RECT 1258.170 145.220 1258.490 145.280 ;
        RECT 1257.710 137.940 1258.030 138.000 ;
        RECT 1257.515 137.800 1258.030 137.940 ;
        RECT 1257.710 137.740 1258.030 137.800 ;
        RECT 1257.725 90.000 1258.015 90.045 ;
        RECT 1258.170 90.000 1258.490 90.060 ;
        RECT 1257.725 89.860 1258.490 90.000 ;
        RECT 1257.725 89.815 1258.015 89.860 ;
        RECT 1258.170 89.800 1258.490 89.860 ;
      LAYER via ;
        RECT 1258.200 1683.380 1258.460 1683.640 ;
        RECT 1258.200 1635.440 1258.460 1635.700 ;
        RECT 1257.280 1563.020 1257.540 1563.280 ;
        RECT 1257.740 1497.740 1258.000 1498.000 ;
        RECT 1257.740 1448.440 1258.000 1448.700 ;
        RECT 1259.120 1448.440 1259.380 1448.700 ;
        RECT 1257.280 1352.560 1257.540 1352.820 ;
        RECT 1258.200 1352.560 1258.460 1352.820 ;
        RECT 1258.200 1221.660 1258.460 1221.920 ;
        RECT 1257.740 1220.980 1258.000 1221.240 ;
        RECT 1257.740 1103.680 1258.000 1103.940 ;
        RECT 1257.740 1048.940 1258.000 1049.200 ;
        RECT 1257.740 1007.120 1258.000 1007.380 ;
        RECT 1258.660 1007.120 1258.920 1007.380 ;
        RECT 1258.200 869.420 1258.460 869.680 ;
        RECT 1258.660 869.420 1258.920 869.680 ;
        RECT 1257.740 710.640 1258.000 710.900 ;
        RECT 1258.200 710.640 1258.460 710.900 ;
        RECT 1256.820 651.820 1257.080 652.080 ;
        RECT 1257.740 651.820 1258.000 652.080 ;
        RECT 1257.740 510.380 1258.000 510.640 ;
        RECT 1258.200 420.620 1258.460 420.880 ;
        RECT 1257.740 282.920 1258.000 283.180 ;
        RECT 1259.120 282.920 1259.380 283.180 ;
        RECT 1259.120 275.780 1259.380 276.040 ;
        RECT 1258.200 228.180 1258.460 228.440 ;
        RECT 1257.740 227.500 1258.000 227.760 ;
        RECT 1258.200 227.500 1258.460 227.760 ;
        RECT 1257.740 145.220 1258.000 145.480 ;
        RECT 1258.200 145.220 1258.460 145.480 ;
        RECT 1257.740 137.740 1258.000 138.000 ;
        RECT 1258.200 89.800 1258.460 90.060 ;
      LAYER met2 ;
        RECT 1258.190 1700.000 1258.470 1704.000 ;
        RECT 1258.260 1691.570 1258.400 1700.000 ;
        RECT 1257.800 1691.430 1258.400 1691.570 ;
        RECT 1257.800 1690.890 1257.940 1691.430 ;
        RECT 1257.800 1690.750 1258.400 1690.890 ;
        RECT 1258.260 1683.670 1258.400 1690.750 ;
        RECT 1258.200 1683.350 1258.460 1683.670 ;
        RECT 1258.200 1635.410 1258.460 1635.730 ;
        RECT 1258.260 1618.130 1258.400 1635.410 ;
        RECT 1257.340 1617.990 1258.400 1618.130 ;
        RECT 1257.340 1563.310 1257.480 1617.990 ;
        RECT 1257.280 1562.990 1257.540 1563.310 ;
        RECT 1257.740 1497.710 1258.000 1498.030 ;
        RECT 1257.800 1448.730 1257.940 1497.710 ;
        RECT 1257.740 1448.410 1258.000 1448.730 ;
        RECT 1259.120 1448.410 1259.380 1448.730 ;
        RECT 1259.180 1442.125 1259.320 1448.410 ;
        RECT 1256.810 1441.755 1257.090 1442.125 ;
        RECT 1259.110 1441.755 1259.390 1442.125 ;
        RECT 1256.880 1399.850 1257.020 1441.755 ;
        RECT 1256.880 1399.710 1257.480 1399.850 ;
        RECT 1257.340 1352.850 1257.480 1399.710 ;
        RECT 1257.280 1352.530 1257.540 1352.850 ;
        RECT 1258.200 1352.530 1258.460 1352.850 ;
        RECT 1258.260 1328.450 1258.400 1352.530 ;
        RECT 1258.260 1328.310 1258.860 1328.450 ;
        RECT 1258.720 1273.370 1258.860 1328.310 ;
        RECT 1258.260 1273.230 1258.860 1273.370 ;
        RECT 1258.260 1221.950 1258.400 1273.230 ;
        RECT 1258.200 1221.630 1258.460 1221.950 ;
        RECT 1257.740 1220.950 1258.000 1221.270 ;
        RECT 1257.800 1186.330 1257.940 1220.950 ;
        RECT 1257.800 1186.190 1258.400 1186.330 ;
        RECT 1258.260 1135.330 1258.400 1186.190 ;
        RECT 1257.800 1135.190 1258.400 1135.330 ;
        RECT 1257.800 1103.970 1257.940 1135.190 ;
        RECT 1257.740 1103.650 1258.000 1103.970 ;
        RECT 1257.740 1048.910 1258.000 1049.230 ;
        RECT 1257.800 1007.410 1257.940 1048.910 ;
        RECT 1257.740 1007.090 1258.000 1007.410 ;
        RECT 1258.660 1007.090 1258.920 1007.410 ;
        RECT 1258.720 869.710 1258.860 1007.090 ;
        RECT 1258.200 869.390 1258.460 869.710 ;
        RECT 1258.660 869.390 1258.920 869.710 ;
        RECT 1258.260 835.450 1258.400 869.390 ;
        RECT 1258.260 835.310 1258.860 835.450 ;
        RECT 1258.720 831.370 1258.860 835.310 ;
        RECT 1257.800 831.230 1258.860 831.370 ;
        RECT 1257.800 710.930 1257.940 831.230 ;
        RECT 1257.740 710.610 1258.000 710.930 ;
        RECT 1258.200 710.610 1258.460 710.930 ;
        RECT 1258.260 699.450 1258.400 710.610 ;
        RECT 1257.800 699.310 1258.400 699.450 ;
        RECT 1257.800 652.110 1257.940 699.310 ;
        RECT 1256.820 651.790 1257.080 652.110 ;
        RECT 1257.740 651.790 1258.000 652.110 ;
        RECT 1256.880 628.165 1257.020 651.790 ;
        RECT 1256.810 627.795 1257.090 628.165 ;
        RECT 1257.730 627.795 1258.010 628.165 ;
        RECT 1257.800 603.570 1257.940 627.795 ;
        RECT 1257.800 603.430 1258.400 603.570 ;
        RECT 1258.260 532.285 1258.400 603.430 ;
        RECT 1258.190 531.915 1258.470 532.285 ;
        RECT 1257.730 531.235 1258.010 531.605 ;
        RECT 1257.800 510.670 1257.940 531.235 ;
        RECT 1257.740 510.350 1258.000 510.670 ;
        RECT 1258.200 420.590 1258.460 420.910 ;
        RECT 1258.260 396.170 1258.400 420.590 ;
        RECT 1257.800 396.030 1258.400 396.170 ;
        RECT 1257.800 283.210 1257.940 396.030 ;
        RECT 1257.740 282.890 1258.000 283.210 ;
        RECT 1259.120 282.890 1259.380 283.210 ;
        RECT 1259.180 276.070 1259.320 282.890 ;
        RECT 1259.120 275.750 1259.380 276.070 ;
        RECT 1258.200 228.150 1258.460 228.470 ;
        RECT 1258.260 227.790 1258.400 228.150 ;
        RECT 1257.740 227.470 1258.000 227.790 ;
        RECT 1258.200 227.470 1258.460 227.790 ;
        RECT 1257.800 186.050 1257.940 227.470 ;
        RECT 1257.800 185.910 1258.400 186.050 ;
        RECT 1258.260 145.510 1258.400 185.910 ;
        RECT 1257.740 145.190 1258.000 145.510 ;
        RECT 1258.200 145.190 1258.460 145.510 ;
        RECT 1257.800 138.030 1257.940 145.190 ;
        RECT 1257.740 137.710 1258.000 138.030 ;
        RECT 1258.200 89.770 1258.460 90.090 ;
        RECT 1258.260 44.725 1258.400 89.770 ;
        RECT 401.210 44.355 401.490 44.725 ;
        RECT 1258.190 44.355 1258.470 44.725 ;
        RECT 401.280 2.400 401.420 44.355 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 1256.810 1441.800 1257.090 1442.080 ;
        RECT 1259.110 1441.800 1259.390 1442.080 ;
        RECT 1256.810 627.840 1257.090 628.120 ;
        RECT 1257.730 627.840 1258.010 628.120 ;
        RECT 1258.190 531.960 1258.470 532.240 ;
        RECT 1257.730 531.280 1258.010 531.560 ;
        RECT 401.210 44.400 401.490 44.680 ;
        RECT 1258.190 44.400 1258.470 44.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1257.705 1014.370 1258.035 1014.385 ;
        RECT 1258.625 1014.370 1258.955 1014.385 ;
        RECT 1257.705 1014.070 1258.955 1014.370 ;
        RECT 1257.705 1014.055 1258.035 1014.070 ;
        RECT 1258.625 1014.055 1258.955 1014.070 ;
        RECT 401.185 46.730 401.515 46.745 ;
        RECT 1257.705 46.730 1258.035 46.745 ;
        RECT 401.185 46.430 1258.035 46.730 ;
        RECT 401.185 46.415 401.515 46.430 ;
        RECT 1257.705 46.415 1258.035 46.430 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1256.785 1442.090 1257.115 1442.105 ;
        RECT 1259.085 1442.090 1259.415 1442.105 ;
        RECT 1256.785 1441.790 1259.415 1442.090 ;
        RECT 1256.785 1441.775 1257.115 1441.790 ;
        RECT 1259.085 1441.775 1259.415 1441.790 ;
        RECT 1256.785 628.130 1257.115 628.145 ;
        RECT 1257.705 628.130 1258.035 628.145 ;
        RECT 1256.785 627.830 1258.035 628.130 ;
        RECT 1256.785 627.815 1257.115 627.830 ;
        RECT 1257.705 627.815 1258.035 627.830 ;
        RECT 1258.165 532.250 1258.495 532.265 ;
        RECT 1257.950 531.935 1258.495 532.250 ;
        RECT 1257.950 531.585 1258.250 531.935 ;
        RECT 1257.705 531.270 1258.250 531.585 ;
        RECT 1257.705 531.255 1258.035 531.270 ;
        RECT 401.185 44.690 401.515 44.705 ;
        RECT 1258.165 44.690 1258.495 44.705 ;
        RECT 401.185 44.390 1258.495 44.690 ;
        RECT 401.185 44.375 401.515 44.390 ;
        RECT 1258.165 44.375 1258.495 44.390 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.170 38.320 62.490 38.380 ;
        RECT 1167.090 38.320 1167.410 38.380 ;
        RECT 62.170 38.180 1167.410 38.320 ;
        RECT 62.170 38.120 62.490 38.180 ;
        RECT 1167.090 38.120 1167.410 38.180 ;
      LAYER via ;
        RECT 62.200 38.120 62.460 38.380 ;
        RECT 1167.120 38.120 1167.380 38.380 ;
      LAYER met2 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 62.050 -4.800 62.610 0.300 ;
=======
        RECT 1166.190 1700.410 1166.470 1704.000 ;
        RECT 1166.190 1700.270 1167.320 1700.410 ;
        RECT 1166.190 1700.000 1166.470 1700.270 ;
        RECT 1167.180 38.605 1167.320 1700.270 ;
        RECT 62.190 38.235 62.470 38.605 ;
        RECT 1167.110 38.235 1167.390 38.605 ;
        RECT 62.260 2.400 62.400 38.235 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 62.190 38.280 62.470 38.560 ;
        RECT 1167.110 38.280 1167.390 38.560 ;
      LAYER met3 ;
        RECT 62.165 38.570 62.495 38.585 ;
        RECT 1167.085 38.570 1167.415 38.585 ;
        RECT 62.165 38.270 1167.415 38.570 ;
        RECT 62.165 38.255 62.495 38.270 ;
        RECT 1167.085 38.255 1167.415 38.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1166.650 1700.410 1166.930 1704.000 ;
        RECT 1166.650 1700.270 1167.320 1700.410 ;
        RECT 1166.650 1700.000 1166.930 1700.270 ;
        RECT 1167.180 38.410 1167.320 1700.270 ;
        RECT 62.200 38.090 62.460 38.410 ;
        RECT 1167.120 38.090 1167.380 38.410 ;
        RECT 62.260 2.400 62.400 38.090 ;
        RECT 62.050 -4.800 62.610 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 419.130 45.800 419.450 45.860 ;
        RECT 1263.690 45.800 1264.010 45.860 ;
        RECT 419.130 45.660 1264.010 45.800 ;
        RECT 419.130 45.600 419.450 45.660 ;
        RECT 1263.690 45.600 1264.010 45.660 ;
      LAYER via ;
        RECT 419.160 45.600 419.420 45.860 ;
        RECT 1263.720 45.600 1263.980 45.860 ;
      LAYER met2 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 419.010 -4.800 419.570 0.300 ;
=======
        RECT 1262.790 1700.000 1263.070 1704.000 ;
        RECT 1262.860 47.445 1263.000 1700.000 ;
        RECT 419.150 47.075 419.430 47.445 ;
        RECT 1262.790 47.075 1263.070 47.445 ;
        RECT 419.220 2.400 419.360 47.075 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 419.150 47.120 419.430 47.400 ;
        RECT 1262.790 47.120 1263.070 47.400 ;
      LAYER met3 ;
        RECT 419.125 47.410 419.455 47.425 ;
        RECT 1262.765 47.410 1263.095 47.425 ;
        RECT 419.125 47.110 1263.095 47.410 ;
        RECT 419.125 47.095 419.455 47.110 ;
        RECT 1262.765 47.095 1263.095 47.110 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1263.250 1700.410 1263.530 1704.000 ;
        RECT 1263.250 1700.270 1263.920 1700.410 ;
        RECT 1263.250 1700.000 1263.530 1700.270 ;
        RECT 1263.780 45.890 1263.920 1700.270 ;
        RECT 419.160 45.570 419.420 45.890 ;
        RECT 1263.720 45.570 1263.980 45.890 ;
        RECT 419.220 2.400 419.360 45.570 ;
        RECT 419.010 -4.800 419.570 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 0.300 ;
=======
      LAYER met1 ;
        RECT 1263.230 1665.560 1263.550 1665.620 ;
        RECT 1266.450 1665.560 1266.770 1665.620 ;
        RECT 1263.230 1665.420 1266.770 1665.560 ;
        RECT 1263.230 1665.360 1263.550 1665.420 ;
        RECT 1266.450 1665.360 1266.770 1665.420 ;
      LAYER via ;
        RECT 1263.260 1665.360 1263.520 1665.620 ;
        RECT 1266.480 1665.360 1266.740 1665.620 ;
      LAYER met2 ;
        RECT 1267.390 1700.410 1267.670 1704.000 ;
        RECT 1266.540 1700.270 1267.670 1700.410 ;
        RECT 1266.540 1665.650 1266.680 1700.270 ;
        RECT 1267.390 1700.000 1267.670 1700.270 ;
        RECT 1263.260 1665.330 1263.520 1665.650 ;
        RECT 1266.480 1665.330 1266.740 1665.650 ;
        RECT 1263.320 48.125 1263.460 1665.330 ;
        RECT 436.630 47.755 436.910 48.125 ;
        RECT 1263.250 47.755 1263.530 48.125 ;
        RECT 436.700 2.400 436.840 47.755 ;
=======
      LAYER li1 ;
        RECT 1265.145 869.465 1265.315 932.535 ;
        RECT 1265.145 752.165 1265.315 759.475 ;
        RECT 1265.145 614.125 1265.315 662.235 ;
        RECT 1265.605 462.485 1265.775 510.595 ;
        RECT 1265.145 372.725 1265.315 420.835 ;
        RECT 1265.145 241.485 1265.315 265.795 ;
      LAYER mcon ;
        RECT 1265.145 932.365 1265.315 932.535 ;
        RECT 1265.145 759.305 1265.315 759.475 ;
        RECT 1265.145 662.065 1265.315 662.235 ;
        RECT 1265.605 510.425 1265.775 510.595 ;
        RECT 1265.145 420.665 1265.315 420.835 ;
        RECT 1265.145 265.625 1265.315 265.795 ;
      LAYER met1 ;
        RECT 1265.070 1545.880 1265.390 1545.940 ;
        RECT 1265.530 1545.880 1265.850 1545.940 ;
        RECT 1265.070 1545.740 1265.850 1545.880 ;
        RECT 1265.070 1545.680 1265.390 1545.740 ;
        RECT 1265.530 1545.680 1265.850 1545.740 ;
        RECT 1265.070 1497.600 1265.390 1497.660 ;
        RECT 1265.530 1497.600 1265.850 1497.660 ;
        RECT 1265.070 1497.460 1265.850 1497.600 ;
        RECT 1265.070 1497.400 1265.390 1497.460 ;
        RECT 1265.530 1497.400 1265.850 1497.460 ;
        RECT 1265.530 1449.660 1265.850 1449.720 ;
        RECT 1265.160 1449.520 1265.850 1449.660 ;
        RECT 1265.160 1449.040 1265.300 1449.520 ;
        RECT 1265.530 1449.460 1265.850 1449.520 ;
        RECT 1265.070 1448.780 1265.390 1449.040 ;
        RECT 1265.070 1352.760 1265.390 1352.820 ;
        RECT 1265.530 1352.760 1265.850 1352.820 ;
        RECT 1265.070 1352.620 1265.850 1352.760 ;
        RECT 1265.070 1352.560 1265.390 1352.620 ;
        RECT 1265.530 1352.560 1265.850 1352.620 ;
        RECT 1264.610 1249.060 1264.930 1249.120 ;
        RECT 1265.530 1249.060 1265.850 1249.120 ;
        RECT 1264.610 1248.920 1265.850 1249.060 ;
        RECT 1264.610 1248.860 1264.930 1248.920 ;
        RECT 1265.530 1248.860 1265.850 1248.920 ;
        RECT 1264.610 1200.780 1264.930 1200.840 ;
        RECT 1265.070 1200.780 1265.390 1200.840 ;
        RECT 1264.610 1200.640 1265.390 1200.780 ;
        RECT 1264.610 1200.580 1264.930 1200.640 ;
        RECT 1265.070 1200.580 1265.390 1200.640 ;
        RECT 1265.070 1007.320 1265.390 1007.380 ;
        RECT 1265.990 1007.320 1266.310 1007.380 ;
        RECT 1265.070 1007.180 1266.310 1007.320 ;
        RECT 1265.070 1007.120 1265.390 1007.180 ;
        RECT 1265.990 1007.120 1266.310 1007.180 ;
        RECT 1265.085 932.520 1265.375 932.565 ;
        RECT 1265.990 932.520 1266.310 932.580 ;
        RECT 1265.085 932.380 1266.310 932.520 ;
        RECT 1265.085 932.335 1265.375 932.380 ;
        RECT 1265.990 932.320 1266.310 932.380 ;
        RECT 1265.085 869.620 1265.375 869.665 ;
        RECT 1265.530 869.620 1265.850 869.680 ;
        RECT 1265.085 869.480 1265.850 869.620 ;
        RECT 1265.085 869.435 1265.375 869.480 ;
        RECT 1265.530 869.420 1265.850 869.480 ;
        RECT 1265.085 759.460 1265.375 759.505 ;
        RECT 1265.530 759.460 1265.850 759.520 ;
        RECT 1265.085 759.320 1265.850 759.460 ;
        RECT 1265.085 759.275 1265.375 759.320 ;
        RECT 1265.530 759.260 1265.850 759.320 ;
        RECT 1265.070 752.320 1265.390 752.380 ;
        RECT 1264.875 752.180 1265.390 752.320 ;
        RECT 1265.070 752.120 1265.390 752.180 ;
        RECT 1265.070 662.220 1265.390 662.280 ;
        RECT 1264.875 662.080 1265.390 662.220 ;
        RECT 1265.070 662.020 1265.390 662.080 ;
        RECT 1265.070 614.280 1265.390 614.340 ;
        RECT 1264.875 614.140 1265.390 614.280 ;
        RECT 1265.070 614.080 1265.390 614.140 ;
        RECT 1265.530 510.580 1265.850 510.640 ;
        RECT 1265.335 510.440 1265.850 510.580 ;
        RECT 1265.530 510.380 1265.850 510.440 ;
        RECT 1265.530 462.640 1265.850 462.700 ;
        RECT 1265.530 462.500 1266.045 462.640 ;
        RECT 1265.530 462.440 1265.850 462.500 ;
        RECT 1265.070 420.820 1265.390 420.880 ;
        RECT 1264.875 420.680 1265.390 420.820 ;
        RECT 1265.070 420.620 1265.390 420.680 ;
        RECT 1264.610 372.880 1264.930 372.940 ;
        RECT 1265.085 372.880 1265.375 372.925 ;
        RECT 1264.610 372.740 1265.375 372.880 ;
        RECT 1264.610 372.680 1264.930 372.740 ;
        RECT 1265.085 372.695 1265.375 372.740 ;
        RECT 1264.610 307.260 1264.930 307.320 ;
        RECT 1265.530 307.260 1265.850 307.320 ;
        RECT 1264.610 307.120 1265.850 307.260 ;
        RECT 1264.610 307.060 1264.930 307.120 ;
        RECT 1265.530 307.060 1265.850 307.120 ;
        RECT 1265.085 265.780 1265.375 265.825 ;
        RECT 1265.530 265.780 1265.850 265.840 ;
        RECT 1265.085 265.640 1265.850 265.780 ;
        RECT 1265.085 265.595 1265.375 265.640 ;
        RECT 1265.530 265.580 1265.850 265.640 ;
        RECT 1265.070 241.640 1265.390 241.700 ;
        RECT 1264.875 241.500 1265.390 241.640 ;
        RECT 1265.070 241.440 1265.390 241.500 ;
        RECT 436.610 46.140 436.930 46.200 ;
        RECT 1265.070 46.140 1265.390 46.200 ;
        RECT 436.610 46.000 1265.390 46.140 ;
        RECT 436.610 45.940 436.930 46.000 ;
        RECT 1265.070 45.940 1265.390 46.000 ;
      LAYER via ;
        RECT 1265.100 1545.680 1265.360 1545.940 ;
        RECT 1265.560 1545.680 1265.820 1545.940 ;
        RECT 1265.100 1497.400 1265.360 1497.660 ;
        RECT 1265.560 1497.400 1265.820 1497.660 ;
        RECT 1265.560 1449.460 1265.820 1449.720 ;
        RECT 1265.100 1448.780 1265.360 1449.040 ;
        RECT 1265.100 1352.560 1265.360 1352.820 ;
        RECT 1265.560 1352.560 1265.820 1352.820 ;
        RECT 1264.640 1248.860 1264.900 1249.120 ;
        RECT 1265.560 1248.860 1265.820 1249.120 ;
        RECT 1264.640 1200.580 1264.900 1200.840 ;
        RECT 1265.100 1200.580 1265.360 1200.840 ;
        RECT 1265.100 1007.120 1265.360 1007.380 ;
        RECT 1266.020 1007.120 1266.280 1007.380 ;
        RECT 1266.020 932.320 1266.280 932.580 ;
        RECT 1265.560 869.420 1265.820 869.680 ;
        RECT 1265.560 759.260 1265.820 759.520 ;
        RECT 1265.100 752.120 1265.360 752.380 ;
        RECT 1265.100 662.020 1265.360 662.280 ;
        RECT 1265.100 614.080 1265.360 614.340 ;
        RECT 1265.560 510.380 1265.820 510.640 ;
        RECT 1265.560 462.440 1265.820 462.700 ;
        RECT 1265.100 420.620 1265.360 420.880 ;
        RECT 1264.640 372.680 1264.900 372.940 ;
        RECT 1264.640 307.060 1264.900 307.320 ;
        RECT 1265.560 307.060 1265.820 307.320 ;
        RECT 1265.560 265.580 1265.820 265.840 ;
        RECT 1265.100 241.440 1265.360 241.700 ;
        RECT 436.640 45.940 436.900 46.200 ;
        RECT 1265.100 45.940 1265.360 46.200 ;
      LAYER met2 ;
        RECT 1267.850 1700.410 1268.130 1704.000 ;
        RECT 1267.000 1700.270 1268.130 1700.410 ;
        RECT 1267.000 1677.970 1267.140 1700.270 ;
        RECT 1267.850 1700.000 1268.130 1700.270 ;
        RECT 1265.620 1677.830 1267.140 1677.970 ;
        RECT 1265.620 1545.970 1265.760 1677.830 ;
        RECT 1265.100 1545.650 1265.360 1545.970 ;
        RECT 1265.560 1545.650 1265.820 1545.970 ;
        RECT 1265.160 1497.690 1265.300 1545.650 ;
        RECT 1265.100 1497.370 1265.360 1497.690 ;
        RECT 1265.560 1497.370 1265.820 1497.690 ;
        RECT 1265.620 1449.750 1265.760 1497.370 ;
        RECT 1265.560 1449.430 1265.820 1449.750 ;
        RECT 1265.100 1448.750 1265.360 1449.070 ;
        RECT 1265.160 1352.850 1265.300 1448.750 ;
        RECT 1265.100 1352.530 1265.360 1352.850 ;
        RECT 1265.560 1352.530 1265.820 1352.850 ;
        RECT 1265.620 1328.450 1265.760 1352.530 ;
        RECT 1265.160 1328.310 1265.760 1328.450 ;
        RECT 1265.160 1303.970 1265.300 1328.310 ;
        RECT 1264.700 1303.830 1265.300 1303.970 ;
        RECT 1264.700 1249.150 1264.840 1303.830 ;
        RECT 1264.640 1248.830 1264.900 1249.150 ;
        RECT 1265.560 1248.890 1265.820 1249.150 ;
        RECT 1265.160 1248.830 1265.820 1248.890 ;
        RECT 1265.160 1248.750 1265.760 1248.830 ;
        RECT 1265.160 1221.690 1265.300 1248.750 ;
        RECT 1264.700 1221.550 1265.300 1221.690 ;
        RECT 1264.700 1200.870 1264.840 1221.550 ;
        RECT 1265.160 1200.870 1265.300 1201.025 ;
        RECT 1264.640 1200.550 1264.900 1200.870 ;
        RECT 1265.100 1200.610 1265.360 1200.870 ;
        RECT 1265.100 1200.550 1265.760 1200.610 ;
        RECT 1265.160 1200.470 1265.760 1200.550 ;
        RECT 1265.620 1135.330 1265.760 1200.470 ;
        RECT 1265.160 1135.190 1265.760 1135.330 ;
        RECT 1265.160 1104.165 1265.300 1135.190 ;
        RECT 1265.090 1103.795 1265.370 1104.165 ;
        RECT 1266.010 1103.115 1266.290 1103.485 ;
        RECT 1266.080 1007.605 1266.220 1103.115 ;
        RECT 1265.090 1007.235 1265.370 1007.605 ;
        RECT 1266.010 1007.235 1266.290 1007.605 ;
        RECT 1265.100 1007.090 1265.360 1007.235 ;
        RECT 1266.020 1007.090 1266.280 1007.235 ;
        RECT 1266.080 932.610 1266.220 1007.090 ;
        RECT 1266.020 932.290 1266.280 932.610 ;
        RECT 1265.560 869.390 1265.820 869.710 ;
        RECT 1265.620 835.450 1265.760 869.390 ;
        RECT 1265.620 835.310 1266.220 835.450 ;
        RECT 1266.080 832.050 1266.220 835.310 ;
        RECT 1265.620 831.910 1266.220 832.050 ;
        RECT 1265.620 759.550 1265.760 831.910 ;
        RECT 1265.560 759.230 1265.820 759.550 ;
        RECT 1265.100 752.090 1265.360 752.410 ;
        RECT 1265.160 734.810 1265.300 752.090 ;
        RECT 1265.160 734.670 1265.760 734.810 ;
        RECT 1265.620 662.730 1265.760 734.670 ;
        RECT 1265.160 662.590 1265.760 662.730 ;
        RECT 1265.160 662.310 1265.300 662.590 ;
        RECT 1265.100 661.990 1265.360 662.310 ;
        RECT 1265.100 614.050 1265.360 614.370 ;
        RECT 1265.160 566.170 1265.300 614.050 ;
        RECT 1265.160 566.030 1265.760 566.170 ;
        RECT 1265.620 510.670 1265.760 566.030 ;
        RECT 1265.560 510.350 1265.820 510.670 ;
        RECT 1265.560 462.410 1265.820 462.730 ;
        RECT 1265.620 421.330 1265.760 462.410 ;
        RECT 1265.160 421.190 1265.760 421.330 ;
        RECT 1265.160 420.910 1265.300 421.190 ;
        RECT 1265.100 420.590 1265.360 420.910 ;
        RECT 1264.640 372.650 1264.900 372.970 ;
        RECT 1264.700 307.350 1264.840 372.650 ;
        RECT 1264.640 307.030 1264.900 307.350 ;
        RECT 1265.560 307.030 1265.820 307.350 ;
        RECT 1265.620 265.870 1265.760 307.030 ;
        RECT 1265.560 265.550 1265.820 265.870 ;
        RECT 1265.100 241.410 1265.360 241.730 ;
        RECT 1265.160 46.230 1265.300 241.410 ;
        RECT 436.640 45.910 436.900 46.230 ;
        RECT 1265.100 45.910 1265.360 46.230 ;
        RECT 436.700 2.400 436.840 45.910 ;
>>>>>>> re-updated local openlane
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 1265.090 1103.840 1265.370 1104.120 ;
        RECT 1266.010 1103.160 1266.290 1103.440 ;
        RECT 1265.090 1007.280 1265.370 1007.560 ;
        RECT 1266.010 1007.280 1266.290 1007.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 436.605 48.090 436.935 48.105 ;
        RECT 1263.225 48.090 1263.555 48.105 ;
        RECT 436.605 47.790 1263.555 48.090 ;
        RECT 436.605 47.775 436.935 47.790 ;
        RECT 1263.225 47.775 1263.555 47.790 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1265.065 1104.130 1265.395 1104.145 ;
        RECT 1265.065 1103.815 1265.610 1104.130 ;
        RECT 1265.310 1103.450 1265.610 1103.815 ;
        RECT 1265.985 1103.450 1266.315 1103.465 ;
        RECT 1265.310 1103.150 1266.315 1103.450 ;
        RECT 1265.985 1103.135 1266.315 1103.150 ;
        RECT 1265.065 1007.570 1265.395 1007.585 ;
        RECT 1265.985 1007.570 1266.315 1007.585 ;
        RECT 1265.065 1007.270 1266.315 1007.570 ;
        RECT 1265.065 1007.255 1265.395 1007.270 ;
        RECT 1265.985 1007.255 1266.315 1007.270 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 0.300 ;
=======
      LAYER met1 ;
        RECT 454.550 46.480 454.870 46.540 ;
        RECT 1270.590 46.480 1270.910 46.540 ;
        RECT 454.550 46.340 1270.910 46.480 ;
        RECT 454.550 46.280 454.870 46.340 ;
        RECT 1270.590 46.280 1270.910 46.340 ;
      LAYER via ;
        RECT 454.580 46.280 454.840 46.540 ;
        RECT 1270.620 46.280 1270.880 46.540 ;
      LAYER met2 ;
        RECT 1272.910 1700.410 1273.190 1704.000 ;
        RECT 1271.600 1700.270 1273.190 1700.410 ;
        RECT 1271.600 1659.610 1271.740 1700.270 ;
        RECT 1272.910 1700.000 1273.190 1700.270 ;
        RECT 1270.680 1659.470 1271.740 1659.610 ;
        RECT 1270.680 46.570 1270.820 1659.470 ;
        RECT 454.580 46.250 454.840 46.570 ;
        RECT 1270.620 46.250 1270.880 46.570 ;
        RECT 454.640 2.400 454.780 46.250 ;
        RECT 454.430 -4.800 454.990 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 0.300 ;
=======
      LAYER met1 ;
        RECT 472.490 46.820 472.810 46.880 ;
        RECT 1277.490 46.820 1277.810 46.880 ;
        RECT 472.490 46.680 1277.810 46.820 ;
        RECT 472.490 46.620 472.810 46.680 ;
        RECT 1277.490 46.620 1277.810 46.680 ;
      LAYER via ;
        RECT 472.520 46.620 472.780 46.880 ;
        RECT 1277.520 46.620 1277.780 46.880 ;
      LAYER met2 ;
        RECT 1277.510 1700.000 1277.790 1704.000 ;
        RECT 1277.580 46.910 1277.720 1700.000 ;
        RECT 472.520 46.590 472.780 46.910 ;
        RECT 1277.520 46.590 1277.780 46.910 ;
        RECT 472.580 2.400 472.720 46.590 ;
        RECT 472.370 -4.800 472.930 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 0.300 ;
=======
      LAYER li1 ;
        RECT 1278.485 1490.645 1278.655 1538.755 ;
        RECT 1278.025 1401.225 1278.195 1448.995 ;
        RECT 1278.485 45.305 1278.655 131.155 ;
      LAYER mcon ;
        RECT 1278.485 1538.585 1278.655 1538.755 ;
        RECT 1278.025 1448.825 1278.195 1448.995 ;
        RECT 1278.485 130.985 1278.655 131.155 ;
      LAYER met1 ;
        RECT 1278.410 1539.420 1278.730 1539.480 ;
        RECT 1279.330 1539.420 1279.650 1539.480 ;
        RECT 1278.410 1539.280 1279.650 1539.420 ;
        RECT 1278.410 1539.220 1278.730 1539.280 ;
        RECT 1279.330 1539.220 1279.650 1539.280 ;
        RECT 1278.425 1538.740 1278.715 1538.785 ;
        RECT 1279.330 1538.740 1279.650 1538.800 ;
        RECT 1278.425 1538.600 1279.650 1538.740 ;
        RECT 1278.425 1538.555 1278.715 1538.600 ;
        RECT 1279.330 1538.540 1279.650 1538.600 ;
        RECT 1278.410 1490.800 1278.730 1490.860 ;
        RECT 1278.215 1490.660 1278.730 1490.800 ;
        RECT 1278.410 1490.600 1278.730 1490.660 ;
        RECT 1277.965 1448.980 1278.255 1449.025 ;
        RECT 1278.410 1448.980 1278.730 1449.040 ;
        RECT 1277.965 1448.840 1278.730 1448.980 ;
        RECT 1277.965 1448.795 1278.255 1448.840 ;
        RECT 1278.410 1448.780 1278.730 1448.840 ;
        RECT 1277.950 1401.380 1278.270 1401.440 ;
        RECT 1277.755 1401.240 1278.270 1401.380 ;
        RECT 1277.950 1401.180 1278.270 1401.240 ;
        RECT 1277.950 1269.600 1278.270 1269.860 ;
        RECT 1278.040 1269.120 1278.180 1269.600 ;
        RECT 1278.410 1269.120 1278.730 1269.180 ;
        RECT 1278.040 1268.980 1278.730 1269.120 ;
        RECT 1278.410 1268.920 1278.730 1268.980 ;
        RECT 1278.410 1207.920 1278.730 1207.980 ;
        RECT 1278.040 1207.780 1278.730 1207.920 ;
        RECT 1278.040 1207.640 1278.180 1207.780 ;
        RECT 1278.410 1207.720 1278.730 1207.780 ;
        RECT 1277.950 1207.380 1278.270 1207.640 ;
        RECT 1278.410 959.040 1278.730 959.100 ;
        RECT 1279.330 959.040 1279.650 959.100 ;
        RECT 1278.410 958.900 1279.650 959.040 ;
        RECT 1278.410 958.840 1278.730 958.900 ;
        RECT 1279.330 958.840 1279.650 958.900 ;
        RECT 1277.950 910.760 1278.270 910.820 ;
        RECT 1278.870 910.760 1279.190 910.820 ;
        RECT 1277.950 910.620 1279.190 910.760 ;
        RECT 1277.950 910.560 1278.270 910.620 ;
        RECT 1278.870 910.560 1279.190 910.620 ;
        RECT 1277.950 759.120 1278.270 759.180 ;
        RECT 1278.410 759.120 1278.730 759.180 ;
        RECT 1277.950 758.980 1278.730 759.120 ;
        RECT 1277.950 758.920 1278.270 758.980 ;
        RECT 1278.410 758.920 1278.730 758.980 ;
        RECT 1277.950 572.940 1278.270 573.200 ;
        RECT 1278.040 572.800 1278.180 572.940 ;
        RECT 1278.410 572.800 1278.730 572.860 ;
        RECT 1278.040 572.660 1278.730 572.800 ;
        RECT 1278.410 572.600 1278.730 572.660 ;
        RECT 1277.950 476.240 1278.270 476.300 ;
        RECT 1278.410 476.240 1278.730 476.300 ;
        RECT 1277.950 476.100 1278.730 476.240 ;
        RECT 1277.950 476.040 1278.270 476.100 ;
        RECT 1278.410 476.040 1278.730 476.100 ;
        RECT 1277.950 434.560 1278.270 434.820 ;
        RECT 1278.040 434.420 1278.180 434.560 ;
        RECT 1278.410 434.420 1278.730 434.480 ;
        RECT 1278.040 434.280 1278.730 434.420 ;
        RECT 1278.410 434.220 1278.730 434.280 ;
        RECT 1277.950 186.560 1278.270 186.620 ;
        RECT 1278.410 186.560 1278.730 186.620 ;
        RECT 1277.950 186.420 1278.730 186.560 ;
        RECT 1277.950 186.360 1278.270 186.420 ;
        RECT 1278.410 186.360 1278.730 186.420 ;
        RECT 1277.950 137.740 1278.270 138.000 ;
        RECT 1278.040 137.600 1278.180 137.740 ;
        RECT 1278.410 137.600 1278.730 137.660 ;
        RECT 1278.040 137.460 1278.730 137.600 ;
        RECT 1278.410 137.400 1278.730 137.460 ;
        RECT 1278.410 131.140 1278.730 131.200 ;
        RECT 1278.215 131.000 1278.730 131.140 ;
        RECT 1278.410 130.940 1278.730 131.000 ;
        RECT 490.430 45.460 490.750 45.520 ;
        RECT 1278.425 45.460 1278.715 45.505 ;
        RECT 490.430 45.320 1278.715 45.460 ;
        RECT 490.430 45.260 490.750 45.320 ;
        RECT 1278.425 45.275 1278.715 45.320 ;
      LAYER via ;
        RECT 1278.440 1539.220 1278.700 1539.480 ;
        RECT 1279.360 1539.220 1279.620 1539.480 ;
        RECT 1279.360 1538.540 1279.620 1538.800 ;
        RECT 1278.440 1490.600 1278.700 1490.860 ;
        RECT 1278.440 1448.780 1278.700 1449.040 ;
        RECT 1277.980 1401.180 1278.240 1401.440 ;
        RECT 1277.980 1269.600 1278.240 1269.860 ;
        RECT 1278.440 1268.920 1278.700 1269.180 ;
        RECT 1278.440 1207.720 1278.700 1207.980 ;
        RECT 1277.980 1207.380 1278.240 1207.640 ;
        RECT 1278.440 958.840 1278.700 959.100 ;
        RECT 1279.360 958.840 1279.620 959.100 ;
        RECT 1277.980 910.560 1278.240 910.820 ;
        RECT 1278.900 910.560 1279.160 910.820 ;
        RECT 1277.980 758.920 1278.240 759.180 ;
        RECT 1278.440 758.920 1278.700 759.180 ;
        RECT 1277.980 572.940 1278.240 573.200 ;
        RECT 1278.440 572.600 1278.700 572.860 ;
        RECT 1277.980 476.040 1278.240 476.300 ;
        RECT 1278.440 476.040 1278.700 476.300 ;
        RECT 1277.980 434.560 1278.240 434.820 ;
        RECT 1278.440 434.220 1278.700 434.480 ;
        RECT 1277.980 186.360 1278.240 186.620 ;
        RECT 1278.440 186.360 1278.700 186.620 ;
        RECT 1277.980 137.740 1278.240 138.000 ;
        RECT 1278.440 137.400 1278.700 137.660 ;
        RECT 1278.440 130.940 1278.700 131.200 ;
        RECT 490.460 45.260 490.720 45.520 ;
      LAYER met2 ;
        RECT 1282.110 1700.410 1282.390 1704.000 ;
        RECT 1281.260 1700.270 1282.390 1700.410 ;
        RECT 1281.260 1656.210 1281.400 1700.270 ;
        RECT 1282.110 1700.000 1282.390 1700.270 ;
        RECT 1278.500 1656.070 1281.400 1656.210 ;
        RECT 1278.500 1605.210 1278.640 1656.070 ;
        RECT 1278.040 1605.070 1278.640 1605.210 ;
        RECT 1278.040 1603.850 1278.180 1605.070 ;
        RECT 1278.040 1603.710 1278.640 1603.850 ;
        RECT 1278.500 1539.510 1278.640 1603.710 ;
        RECT 1278.440 1539.190 1278.700 1539.510 ;
        RECT 1279.360 1539.190 1279.620 1539.510 ;
        RECT 1279.420 1538.830 1279.560 1539.190 ;
        RECT 1279.360 1538.510 1279.620 1538.830 ;
        RECT 1278.440 1490.570 1278.700 1490.890 ;
        RECT 1278.500 1449.070 1278.640 1490.570 ;
        RECT 1278.440 1448.750 1278.700 1449.070 ;
        RECT 1277.980 1401.150 1278.240 1401.470 ;
        RECT 1278.040 1269.890 1278.180 1401.150 ;
        RECT 1277.980 1269.570 1278.240 1269.890 ;
        RECT 1278.440 1268.890 1278.700 1269.210 ;
        RECT 1278.500 1208.010 1278.640 1268.890 ;
        RECT 1278.440 1207.690 1278.700 1208.010 ;
        RECT 1277.980 1207.350 1278.240 1207.670 ;
        RECT 1278.040 1200.725 1278.180 1207.350 ;
        RECT 1277.970 1200.355 1278.250 1200.725 ;
        RECT 1278.890 1200.355 1279.170 1200.725 ;
        RECT 1278.960 1176.130 1279.100 1200.355 ;
        RECT 1278.500 1175.990 1279.100 1176.130 ;
        RECT 1278.500 1056.565 1278.640 1175.990 ;
        RECT 1278.430 1056.195 1278.710 1056.565 ;
        RECT 1278.430 1055.515 1278.710 1055.885 ;
        RECT 1278.500 959.130 1278.640 1055.515 ;
        RECT 1278.440 958.810 1278.700 959.130 ;
        RECT 1279.360 958.810 1279.620 959.130 ;
        RECT 1279.420 911.045 1279.560 958.810 ;
        RECT 1277.970 910.675 1278.250 911.045 ;
        RECT 1277.980 910.530 1278.240 910.675 ;
        RECT 1278.900 910.530 1279.160 910.850 ;
        RECT 1279.350 910.675 1279.630 911.045 ;
        RECT 1278.960 821.285 1279.100 910.530 ;
        RECT 1277.970 820.915 1278.250 821.285 ;
        RECT 1278.890 820.915 1279.170 821.285 ;
        RECT 1278.040 759.210 1278.180 820.915 ;
        RECT 1277.980 758.890 1278.240 759.210 ;
        RECT 1278.440 758.890 1278.700 759.210 ;
        RECT 1278.500 758.610 1278.640 758.890 ;
        RECT 1278.500 758.470 1279.100 758.610 ;
        RECT 1278.960 688.570 1279.100 758.470 ;
        RECT 1278.500 688.430 1279.100 688.570 ;
        RECT 1278.500 628.845 1278.640 688.430 ;
        RECT 1278.430 628.475 1278.710 628.845 ;
        RECT 1277.970 627.795 1278.250 628.165 ;
        RECT 1278.040 573.230 1278.180 627.795 ;
        RECT 1277.980 572.910 1278.240 573.230 ;
        RECT 1278.440 572.570 1278.700 572.890 ;
        RECT 1278.500 476.330 1278.640 572.570 ;
        RECT 1277.980 476.010 1278.240 476.330 ;
        RECT 1278.440 476.010 1278.700 476.330 ;
        RECT 1278.040 434.850 1278.180 476.010 ;
        RECT 1277.980 434.530 1278.240 434.850 ;
        RECT 1278.440 434.190 1278.700 434.510 ;
        RECT 1278.500 338.370 1278.640 434.190 ;
        RECT 1278.040 338.230 1278.640 338.370 ;
        RECT 1278.040 186.650 1278.180 338.230 ;
        RECT 1277.980 186.330 1278.240 186.650 ;
        RECT 1278.440 186.330 1278.700 186.650 ;
        RECT 1278.500 162.250 1278.640 186.330 ;
        RECT 1278.040 162.110 1278.640 162.250 ;
        RECT 1278.040 138.030 1278.180 162.110 ;
        RECT 1277.980 137.710 1278.240 138.030 ;
        RECT 1278.440 137.370 1278.700 137.690 ;
        RECT 1278.500 131.230 1278.640 137.370 ;
        RECT 1278.440 130.910 1278.700 131.230 ;
        RECT 490.460 45.230 490.720 45.550 ;
        RECT 490.520 2.400 490.660 45.230 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 1277.970 1200.400 1278.250 1200.680 ;
        RECT 1278.890 1200.400 1279.170 1200.680 ;
        RECT 1278.430 1056.240 1278.710 1056.520 ;
        RECT 1278.430 1055.560 1278.710 1055.840 ;
        RECT 1277.970 910.720 1278.250 911.000 ;
        RECT 1279.350 910.720 1279.630 911.000 ;
        RECT 1277.970 820.960 1278.250 821.240 ;
        RECT 1278.890 820.960 1279.170 821.240 ;
        RECT 1278.430 628.520 1278.710 628.800 ;
        RECT 1277.970 627.840 1278.250 628.120 ;
      LAYER met3 ;
        RECT 1277.945 1200.690 1278.275 1200.705 ;
        RECT 1278.865 1200.690 1279.195 1200.705 ;
        RECT 1277.945 1200.390 1279.195 1200.690 ;
        RECT 1277.945 1200.375 1278.275 1200.390 ;
        RECT 1278.865 1200.375 1279.195 1200.390 ;
        RECT 1278.405 1056.530 1278.735 1056.545 ;
        RECT 1278.190 1056.215 1278.735 1056.530 ;
        RECT 1278.190 1055.865 1278.490 1056.215 ;
        RECT 1278.190 1055.550 1278.735 1055.865 ;
        RECT 1278.405 1055.535 1278.735 1055.550 ;
        RECT 1277.945 911.010 1278.275 911.025 ;
        RECT 1279.325 911.010 1279.655 911.025 ;
        RECT 1277.945 910.710 1279.655 911.010 ;
        RECT 1277.945 910.695 1278.275 910.710 ;
        RECT 1279.325 910.695 1279.655 910.710 ;
        RECT 1277.945 821.250 1278.275 821.265 ;
        RECT 1278.865 821.250 1279.195 821.265 ;
        RECT 1277.945 820.950 1279.195 821.250 ;
        RECT 1277.945 820.935 1278.275 820.950 ;
        RECT 1278.865 820.935 1279.195 820.950 ;
        RECT 1278.405 628.810 1278.735 628.825 ;
        RECT 1278.190 628.495 1278.735 628.810 ;
        RECT 1278.190 628.145 1278.490 628.495 ;
        RECT 1277.945 627.830 1278.490 628.145 ;
        RECT 1277.945 627.815 1278.275 627.830 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1277.030 1678.140 1277.350 1678.200 ;
        RECT 1281.170 1678.140 1281.490 1678.200 ;
        RECT 1277.030 1678.000 1281.490 1678.140 ;
        RECT 1277.030 1677.940 1277.350 1678.000 ;
        RECT 1281.170 1677.940 1281.490 1678.000 ;
        RECT 490.430 47.160 490.750 47.220 ;
        RECT 1277.030 47.160 1277.350 47.220 ;
        RECT 490.430 47.020 1277.350 47.160 ;
        RECT 490.430 46.960 490.750 47.020 ;
        RECT 1277.030 46.960 1277.350 47.020 ;
      LAYER via ;
        RECT 1277.060 1677.940 1277.320 1678.200 ;
        RECT 1281.200 1677.940 1281.460 1678.200 ;
        RECT 490.460 46.960 490.720 47.220 ;
        RECT 1277.060 46.960 1277.320 47.220 ;
      LAYER met2 ;
        RECT 1282.570 1700.410 1282.850 1704.000 ;
        RECT 1281.260 1700.270 1282.850 1700.410 ;
        RECT 1281.260 1678.230 1281.400 1700.270 ;
        RECT 1282.570 1700.000 1282.850 1700.270 ;
        RECT 1277.060 1677.910 1277.320 1678.230 ;
        RECT 1281.200 1677.910 1281.460 1678.230 ;
        RECT 1277.120 47.250 1277.260 1677.910 ;
        RECT 490.460 46.930 490.720 47.250 ;
        RECT 1277.060 46.930 1277.320 47.250 ;
        RECT 490.520 2.400 490.660 46.930 ;
        RECT 490.310 -4.800 490.870 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 0.300 ;
=======
      LAYER met1 ;
        RECT 1285.310 690.440 1285.630 690.500 ;
        RECT 1284.940 690.300 1285.630 690.440 ;
        RECT 1284.940 689.820 1285.080 690.300 ;
        RECT 1285.310 690.240 1285.630 690.300 ;
        RECT 1284.850 689.560 1285.170 689.820 ;
        RECT 510.210 54.300 510.530 54.360 ;
        RECT 1284.390 54.300 1284.710 54.360 ;
        RECT 510.210 54.160 1284.710 54.300 ;
        RECT 510.210 54.100 510.530 54.160 ;
        RECT 1284.390 54.100 1284.710 54.160 ;
        RECT 507.910 15.540 508.230 15.600 ;
        RECT 510.210 15.540 510.530 15.600 ;
        RECT 507.910 15.400 510.530 15.540 ;
        RECT 507.910 15.340 508.230 15.400 ;
        RECT 510.210 15.340 510.530 15.400 ;
      LAYER via ;
        RECT 1285.340 690.240 1285.600 690.500 ;
        RECT 1284.880 689.560 1285.140 689.820 ;
        RECT 510.240 54.100 510.500 54.360 ;
        RECT 1284.420 54.100 1284.680 54.360 ;
        RECT 507.940 15.340 508.200 15.600 ;
        RECT 510.240 15.340 510.500 15.600 ;
      LAYER met2 ;
        RECT 1287.630 1700.410 1287.910 1704.000 ;
        RECT 1286.780 1700.270 1287.910 1700.410 ;
        RECT 1286.780 1684.770 1286.920 1700.270 ;
        RECT 1287.630 1700.000 1287.910 1700.270 ;
        RECT 1284.940 1684.630 1286.920 1684.770 ;
        RECT 1284.940 1414.810 1285.080 1684.630 ;
        RECT 1284.480 1414.670 1285.080 1414.810 ;
        RECT 1284.480 1414.130 1284.620 1414.670 ;
        RECT 1284.480 1413.990 1285.080 1414.130 ;
        RECT 1284.940 1318.250 1285.080 1413.990 ;
        RECT 1284.480 1318.110 1285.080 1318.250 ;
        RECT 1284.480 1317.570 1284.620 1318.110 ;
        RECT 1284.480 1317.430 1285.080 1317.570 ;
        RECT 1284.940 1221.690 1285.080 1317.430 ;
        RECT 1284.480 1221.550 1285.080 1221.690 ;
        RECT 1284.480 1221.010 1284.620 1221.550 ;
        RECT 1284.480 1220.870 1285.080 1221.010 ;
        RECT 1284.940 1125.130 1285.080 1220.870 ;
        RECT 1284.480 1124.990 1285.080 1125.130 ;
        RECT 1284.480 1124.450 1284.620 1124.990 ;
        RECT 1284.480 1124.310 1285.080 1124.450 ;
        RECT 1284.940 1028.570 1285.080 1124.310 ;
        RECT 1284.480 1028.430 1285.080 1028.570 ;
        RECT 1284.480 1027.890 1284.620 1028.430 ;
        RECT 1284.480 1027.750 1285.080 1027.890 ;
        RECT 1284.940 932.010 1285.080 1027.750 ;
        RECT 1284.480 931.870 1285.080 932.010 ;
        RECT 1284.480 931.330 1284.620 931.870 ;
        RECT 1284.480 931.190 1285.080 931.330 ;
        RECT 1284.940 835.450 1285.080 931.190 ;
        RECT 1284.480 835.310 1285.080 835.450 ;
        RECT 1284.480 834.770 1284.620 835.310 ;
        RECT 1284.480 834.630 1285.080 834.770 ;
        RECT 1284.940 738.890 1285.080 834.630 ;
        RECT 1284.480 738.750 1285.080 738.890 ;
        RECT 1284.480 738.210 1284.620 738.750 ;
        RECT 1284.480 738.070 1285.540 738.210 ;
        RECT 1285.400 690.530 1285.540 738.070 ;
        RECT 1285.340 690.210 1285.600 690.530 ;
        RECT 1284.880 689.530 1285.140 689.850 ;
        RECT 1284.940 642.330 1285.080 689.530 ;
        RECT 1284.480 642.190 1285.080 642.330 ;
        RECT 1284.480 641.650 1284.620 642.190 ;
        RECT 1284.480 641.510 1285.080 641.650 ;
        RECT 1284.940 545.770 1285.080 641.510 ;
        RECT 1284.480 545.630 1285.080 545.770 ;
        RECT 1284.480 545.090 1284.620 545.630 ;
        RECT 1284.480 544.950 1285.080 545.090 ;
        RECT 1284.940 449.210 1285.080 544.950 ;
        RECT 1284.480 449.070 1285.080 449.210 ;
        RECT 1284.480 448.530 1284.620 449.070 ;
        RECT 1284.480 448.390 1285.080 448.530 ;
        RECT 1284.940 351.970 1285.080 448.390 ;
        RECT 1284.480 351.830 1285.080 351.970 ;
        RECT 1284.480 351.290 1284.620 351.830 ;
        RECT 1284.480 351.150 1285.080 351.290 ;
        RECT 1284.940 255.410 1285.080 351.150 ;
        RECT 1284.480 255.270 1285.080 255.410 ;
        RECT 1284.480 254.730 1284.620 255.270 ;
        RECT 1284.480 254.590 1285.080 254.730 ;
        RECT 1284.940 158.850 1285.080 254.590 ;
        RECT 1284.480 158.710 1285.080 158.850 ;
        RECT 1284.480 158.170 1284.620 158.710 ;
        RECT 1284.480 158.030 1285.080 158.170 ;
        RECT 1284.940 62.290 1285.080 158.030 ;
        RECT 1284.480 62.150 1285.080 62.290 ;
        RECT 1284.480 54.390 1284.620 62.150 ;
        RECT 510.240 54.070 510.500 54.390 ;
        RECT 1284.420 54.070 1284.680 54.390 ;
        RECT 510.300 15.630 510.440 54.070 ;
        RECT 507.940 15.310 508.200 15.630 ;
        RECT 510.240 15.310 510.500 15.630 ;
        RECT 508.000 2.400 508.140 15.310 ;
        RECT 507.790 -4.800 508.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 0.300 ;
=======
      LAYER met1 ;
        RECT 530.910 54.640 531.230 54.700 ;
        RECT 1292.210 54.640 1292.530 54.700 ;
        RECT 530.910 54.500 1292.530 54.640 ;
        RECT 530.910 54.440 531.230 54.500 ;
        RECT 1292.210 54.440 1292.530 54.500 ;
        RECT 525.850 15.540 526.170 15.600 ;
        RECT 530.910 15.540 531.230 15.600 ;
        RECT 525.850 15.400 531.230 15.540 ;
        RECT 525.850 15.340 526.170 15.400 ;
        RECT 530.910 15.340 531.230 15.400 ;
      LAYER via ;
        RECT 530.940 54.440 531.200 54.700 ;
        RECT 1292.240 54.440 1292.500 54.700 ;
        RECT 525.880 15.340 526.140 15.600 ;
        RECT 530.940 15.340 531.200 15.600 ;
      LAYER met2 ;
        RECT 1292.230 1700.000 1292.510 1704.000 ;
        RECT 1292.300 54.730 1292.440 1700.000 ;
        RECT 530.940 54.410 531.200 54.730 ;
        RECT 1292.240 54.410 1292.500 54.730 ;
        RECT 531.000 15.630 531.140 54.410 ;
        RECT 525.880 15.310 526.140 15.630 ;
        RECT 530.940 15.310 531.200 15.630 ;
        RECT 525.940 2.400 526.080 15.310 ;
        RECT 525.730 -4.800 526.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 0.300 ;
=======
      LAYER met1 ;
        RECT 544.710 54.980 545.030 55.040 ;
        RECT 1297.730 54.980 1298.050 55.040 ;
        RECT 544.710 54.840 1298.050 54.980 ;
        RECT 544.710 54.780 545.030 54.840 ;
        RECT 1297.730 54.780 1298.050 54.840 ;
      LAYER via ;
        RECT 544.740 54.780 545.000 55.040 ;
        RECT 1297.760 54.780 1298.020 55.040 ;
      LAYER met2 ;
        RECT 1297.290 1700.410 1297.570 1704.000 ;
        RECT 1297.290 1700.270 1297.960 1700.410 ;
        RECT 1297.290 1700.000 1297.570 1700.270 ;
        RECT 1297.820 55.070 1297.960 1700.270 ;
        RECT 544.740 54.750 545.000 55.070 ;
        RECT 1297.760 54.750 1298.020 55.070 ;
        RECT 544.800 17.410 544.940 54.750 ;
        RECT 543.880 17.270 544.940 17.410 ;
        RECT 543.880 2.400 544.020 17.270 ;
        RECT 543.670 -4.800 544.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 0.300 ;
=======
      LAYER met1 ;
        RECT 1298.190 1678.140 1298.510 1678.200 ;
        RECT 1300.950 1678.140 1301.270 1678.200 ;
        RECT 1298.190 1678.000 1301.270 1678.140 ;
        RECT 1298.190 1677.940 1298.510 1678.000 ;
        RECT 1300.950 1677.940 1301.270 1678.000 ;
        RECT 565.410 51.240 565.730 51.300 ;
        RECT 1298.190 51.240 1298.510 51.300 ;
        RECT 565.410 51.100 1298.510 51.240 ;
        RECT 565.410 51.040 565.730 51.100 ;
        RECT 1298.190 51.040 1298.510 51.100 ;
        RECT 561.730 14.860 562.050 14.920 ;
        RECT 565.410 14.860 565.730 14.920 ;
        RECT 561.730 14.720 565.730 14.860 ;
        RECT 561.730 14.660 562.050 14.720 ;
        RECT 565.410 14.660 565.730 14.720 ;
      LAYER via ;
        RECT 1298.220 1677.940 1298.480 1678.200 ;
        RECT 1300.980 1677.940 1301.240 1678.200 ;
        RECT 565.440 51.040 565.700 51.300 ;
        RECT 1298.220 51.040 1298.480 51.300 ;
        RECT 561.760 14.660 562.020 14.920 ;
        RECT 565.440 14.660 565.700 14.920 ;
      LAYER met2 ;
        RECT 1301.890 1700.410 1302.170 1704.000 ;
        RECT 1301.040 1700.270 1302.170 1700.410 ;
        RECT 1301.040 1678.230 1301.180 1700.270 ;
        RECT 1301.890 1700.000 1302.170 1700.270 ;
        RECT 1298.220 1677.910 1298.480 1678.230 ;
        RECT 1300.980 1677.910 1301.240 1678.230 ;
        RECT 1298.280 51.330 1298.420 1677.910 ;
        RECT 565.440 51.010 565.700 51.330 ;
        RECT 1298.220 51.010 1298.480 51.330 ;
        RECT 565.500 14.950 565.640 51.010 ;
        RECT 561.760 14.630 562.020 14.950 ;
        RECT 565.440 14.630 565.700 14.950 ;
        RECT 561.820 2.400 561.960 14.630 ;
        RECT 561.610 -4.800 562.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 0.300 ;
=======
      LAYER met1 ;
        RECT 585.650 50.900 585.970 50.960 ;
        RECT 1304.630 50.900 1304.950 50.960 ;
        RECT 585.650 50.760 1304.950 50.900 ;
        RECT 585.650 50.700 585.970 50.760 ;
        RECT 1304.630 50.700 1304.950 50.760 ;
        RECT 579.670 14.860 579.990 14.920 ;
        RECT 584.730 14.860 585.050 14.920 ;
        RECT 579.670 14.720 585.050 14.860 ;
        RECT 579.670 14.660 579.990 14.720 ;
        RECT 584.730 14.660 585.050 14.720 ;
      LAYER via ;
        RECT 585.680 50.700 585.940 50.960 ;
        RECT 1304.660 50.700 1304.920 50.960 ;
        RECT 579.700 14.660 579.960 14.920 ;
        RECT 584.760 14.660 585.020 14.920 ;
      LAYER met2 ;
        RECT 1306.950 1700.410 1307.230 1704.000 ;
        RECT 1305.640 1700.270 1307.230 1700.410 ;
        RECT 1305.640 1678.140 1305.780 1700.270 ;
        RECT 1306.950 1700.000 1307.230 1700.270 ;
        RECT 1304.720 1678.000 1305.780 1678.140 ;
        RECT 1304.720 50.990 1304.860 1678.000 ;
        RECT 585.680 50.670 585.940 50.990 ;
        RECT 1304.660 50.670 1304.920 50.990 ;
        RECT 585.740 18.090 585.880 50.670 ;
        RECT 584.820 17.950 585.880 18.090 ;
        RECT 584.820 14.950 584.960 17.950 ;
        RECT 579.700 14.630 579.960 14.950 ;
        RECT 584.760 14.630 585.020 14.950 ;
        RECT 579.760 2.400 579.900 14.630 ;
        RECT 579.550 -4.800 580.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 0.300 ;
=======
      LAYER met1 ;
        RECT 86.550 38.660 86.870 38.720 ;
        RECT 1173.070 38.660 1173.390 38.720 ;
        RECT 86.550 38.520 1173.390 38.660 ;
        RECT 86.550 38.460 86.870 38.520 ;
        RECT 1173.070 38.460 1173.390 38.520 ;
      LAYER via ;
        RECT 86.580 38.460 86.840 38.720 ;
        RECT 1173.100 38.460 1173.360 38.720 ;
      LAYER met2 ;
        RECT 1173.090 1700.000 1173.370 1704.000 ;
        RECT 1173.160 38.750 1173.300 1700.000 ;
        RECT 86.580 38.430 86.840 38.750 ;
        RECT 1173.100 38.430 1173.360 38.750 ;
        RECT 86.640 7.210 86.780 38.430 ;
        RECT 86.180 7.070 86.780 7.210 ;
        RECT 86.180 2.400 86.320 7.070 ;
        RECT 85.970 -4.800 86.530 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 86.110 38.960 86.390 39.240 ;
        RECT 1166.650 38.960 1166.930 39.240 ;
      LAYER met3 ;
        RECT 86.085 39.250 86.415 39.265 ;
        RECT 1166.625 39.250 1166.955 39.265 ;
        RECT 86.085 38.950 1166.955 39.250 ;
        RECT 86.085 38.935 86.415 38.950 ;
        RECT 1166.625 38.935 1166.955 38.950 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 0.300 ;
=======
      LAYER met1 ;
        RECT 599.910 50.560 600.230 50.620 ;
        RECT 1311.990 50.560 1312.310 50.620 ;
        RECT 599.910 50.420 1312.310 50.560 ;
        RECT 599.910 50.360 600.230 50.420 ;
        RECT 1311.990 50.360 1312.310 50.420 ;
        RECT 597.150 14.860 597.470 14.920 ;
        RECT 599.910 14.860 600.230 14.920 ;
        RECT 597.150 14.720 600.230 14.860 ;
        RECT 597.150 14.660 597.470 14.720 ;
        RECT 599.910 14.660 600.230 14.720 ;
      LAYER via ;
        RECT 599.940 50.360 600.200 50.620 ;
        RECT 1312.020 50.360 1312.280 50.620 ;
        RECT 597.180 14.660 597.440 14.920 ;
        RECT 599.940 14.660 600.200 14.920 ;
      LAYER met2 ;
        RECT 1311.550 1700.410 1311.830 1704.000 ;
        RECT 1311.550 1700.270 1312.220 1700.410 ;
        RECT 1311.550 1700.000 1311.830 1700.270 ;
        RECT 1312.080 50.650 1312.220 1700.270 ;
        RECT 599.940 50.330 600.200 50.650 ;
        RECT 1312.020 50.330 1312.280 50.650 ;
        RECT 600.000 14.950 600.140 50.330 ;
        RECT 597.180 14.630 597.440 14.950 ;
        RECT 599.940 14.630 600.200 14.950 ;
        RECT 597.240 2.400 597.380 14.630 ;
        RECT 597.030 -4.800 597.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 0.300 ;
=======
      LAYER met1 ;
        RECT 1311.070 1678.140 1311.390 1678.200 ;
        RECT 1315.210 1678.140 1315.530 1678.200 ;
        RECT 1311.070 1678.000 1315.530 1678.140 ;
        RECT 1311.070 1677.940 1311.390 1678.000 ;
        RECT 1315.210 1677.940 1315.530 1678.000 ;
        RECT 620.610 50.220 620.930 50.280 ;
        RECT 1311.070 50.220 1311.390 50.280 ;
        RECT 620.610 50.080 1311.390 50.220 ;
        RECT 620.610 50.020 620.930 50.080 ;
        RECT 1311.070 50.020 1311.390 50.080 ;
      LAYER via ;
        RECT 1311.100 1677.940 1311.360 1678.200 ;
        RECT 1315.240 1677.940 1315.500 1678.200 ;
        RECT 620.640 50.020 620.900 50.280 ;
        RECT 1311.100 50.020 1311.360 50.280 ;
      LAYER met2 ;
        RECT 1316.610 1700.410 1316.890 1704.000 ;
        RECT 1315.300 1700.270 1316.890 1700.410 ;
        RECT 1315.300 1678.230 1315.440 1700.270 ;
        RECT 1316.610 1700.000 1316.890 1700.270 ;
        RECT 1311.100 1677.910 1311.360 1678.230 ;
        RECT 1315.240 1677.910 1315.500 1678.230 ;
        RECT 1311.160 50.310 1311.300 1677.910 ;
        RECT 620.640 49.990 620.900 50.310 ;
        RECT 1311.100 49.990 1311.360 50.310 ;
        RECT 620.700 17.410 620.840 49.990 ;
        RECT 615.180 17.270 620.840 17.410 ;
        RECT 615.180 2.400 615.320 17.270 ;
        RECT 614.970 -4.800 615.530 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 0.300 ;
=======
      LAYER li1 ;
        RECT 1175.445 1569.185 1175.615 1593.835 ;
        RECT 1174.985 669.545 1175.155 717.655 ;
      LAYER mcon ;
        RECT 1175.445 1593.665 1175.615 1593.835 ;
        RECT 1174.985 717.485 1175.155 717.655 ;
      LAYER met1 ;
        RECT 1175.370 1642.440 1175.690 1642.500 ;
        RECT 1178.590 1642.440 1178.910 1642.500 ;
        RECT 1175.370 1642.300 1178.910 1642.440 ;
        RECT 1175.370 1642.240 1175.690 1642.300 ;
        RECT 1178.590 1642.240 1178.910 1642.300 ;
        RECT 1175.370 1593.820 1175.690 1593.880 ;
        RECT 1175.175 1593.680 1175.690 1593.820 ;
        RECT 1175.370 1593.620 1175.690 1593.680 ;
        RECT 1175.370 1569.340 1175.690 1569.400 ;
        RECT 1175.175 1569.200 1175.690 1569.340 ;
        RECT 1175.370 1569.140 1175.690 1569.200 ;
        RECT 1174.450 741.780 1174.770 741.840 ;
        RECT 1175.370 741.780 1175.690 741.840 ;
        RECT 1174.450 741.640 1175.690 741.780 ;
        RECT 1174.450 741.580 1174.770 741.640 ;
        RECT 1175.370 741.580 1175.690 741.640 ;
        RECT 1174.910 717.640 1175.230 717.700 ;
        RECT 1174.715 717.500 1175.230 717.640 ;
        RECT 1174.910 717.440 1175.230 717.500 ;
        RECT 1174.910 669.700 1175.230 669.760 ;
        RECT 1174.715 669.560 1175.230 669.700 ;
        RECT 1174.910 669.500 1175.230 669.560 ;
        RECT 109.550 39.000 109.870 39.060 ;
        RECT 1174.910 39.000 1175.230 39.060 ;
        RECT 109.550 38.860 1175.230 39.000 ;
        RECT 109.550 38.800 109.870 38.860 ;
        RECT 1174.910 38.800 1175.230 38.860 ;
      LAYER via ;
        RECT 1175.400 1642.240 1175.660 1642.500 ;
        RECT 1178.620 1642.240 1178.880 1642.500 ;
        RECT 1175.400 1593.620 1175.660 1593.880 ;
        RECT 1175.400 1569.140 1175.660 1569.400 ;
        RECT 1174.480 741.580 1174.740 741.840 ;
        RECT 1175.400 741.580 1175.660 741.840 ;
        RECT 1174.940 717.440 1175.200 717.700 ;
        RECT 1174.940 669.500 1175.200 669.760 ;
        RECT 109.580 38.800 109.840 39.060 ;
        RECT 1174.940 38.800 1175.200 39.060 ;
      LAYER met2 ;
        RECT 1179.530 1700.410 1179.810 1704.000 ;
        RECT 1178.680 1700.270 1179.810 1700.410 ;
        RECT 1178.680 1642.530 1178.820 1700.270 ;
        RECT 1179.530 1700.000 1179.810 1700.270 ;
        RECT 1175.400 1642.210 1175.660 1642.530 ;
        RECT 1178.620 1642.210 1178.880 1642.530 ;
        RECT 1175.460 1593.910 1175.600 1642.210 ;
        RECT 1175.400 1593.590 1175.660 1593.910 ;
        RECT 1175.400 1569.110 1175.660 1569.430 ;
        RECT 1175.460 1414.810 1175.600 1569.110 ;
        RECT 1175.000 1414.670 1175.600 1414.810 ;
        RECT 1175.000 1414.130 1175.140 1414.670 ;
        RECT 1175.000 1413.990 1175.600 1414.130 ;
        RECT 1175.460 1318.250 1175.600 1413.990 ;
        RECT 1175.000 1318.110 1175.600 1318.250 ;
        RECT 1175.000 1317.570 1175.140 1318.110 ;
        RECT 1175.000 1317.430 1175.600 1317.570 ;
        RECT 1175.460 1221.690 1175.600 1317.430 ;
        RECT 1175.000 1221.550 1175.600 1221.690 ;
        RECT 1175.000 1221.010 1175.140 1221.550 ;
        RECT 1175.000 1220.870 1175.600 1221.010 ;
        RECT 1175.460 1125.130 1175.600 1220.870 ;
        RECT 1175.000 1124.990 1175.600 1125.130 ;
        RECT 1175.000 1124.450 1175.140 1124.990 ;
        RECT 1175.000 1124.310 1175.600 1124.450 ;
        RECT 1175.460 1028.570 1175.600 1124.310 ;
        RECT 1175.000 1028.430 1175.600 1028.570 ;
        RECT 1175.000 1027.890 1175.140 1028.430 ;
        RECT 1175.000 1027.750 1175.600 1027.890 ;
        RECT 1175.460 932.010 1175.600 1027.750 ;
        RECT 1175.000 931.870 1175.600 932.010 ;
        RECT 1175.000 931.330 1175.140 931.870 ;
        RECT 1175.000 931.190 1175.600 931.330 ;
        RECT 1175.460 835.450 1175.600 931.190 ;
        RECT 1175.000 835.310 1175.600 835.450 ;
        RECT 1175.000 834.770 1175.140 835.310 ;
        RECT 1175.000 834.630 1175.600 834.770 ;
        RECT 1175.460 741.870 1175.600 834.630 ;
        RECT 1174.480 741.550 1174.740 741.870 ;
        RECT 1175.400 741.550 1175.660 741.870 ;
        RECT 1174.540 717.810 1174.680 741.550 ;
        RECT 1174.540 717.730 1175.140 717.810 ;
        RECT 1174.540 717.670 1175.200 717.730 ;
        RECT 1174.940 717.410 1175.200 717.670 ;
        RECT 1174.940 669.470 1175.200 669.790 ;
        RECT 1175.000 650.490 1175.140 669.470 ;
        RECT 1175.000 650.350 1175.600 650.490 ;
        RECT 1175.460 545.770 1175.600 650.350 ;
        RECT 1175.000 545.630 1175.600 545.770 ;
        RECT 1175.000 545.090 1175.140 545.630 ;
        RECT 1175.000 544.950 1175.600 545.090 ;
        RECT 1175.460 449.210 1175.600 544.950 ;
        RECT 1175.000 449.070 1175.600 449.210 ;
        RECT 1175.000 448.530 1175.140 449.070 ;
        RECT 1175.000 448.390 1175.600 448.530 ;
        RECT 1175.460 351.970 1175.600 448.390 ;
        RECT 1175.000 351.830 1175.600 351.970 ;
        RECT 1175.000 351.290 1175.140 351.830 ;
        RECT 1175.000 351.150 1175.600 351.290 ;
        RECT 1175.460 255.410 1175.600 351.150 ;
        RECT 1175.000 255.270 1175.600 255.410 ;
        RECT 1175.000 254.730 1175.140 255.270 ;
        RECT 1175.000 254.590 1175.600 254.730 ;
        RECT 1175.460 158.850 1175.600 254.590 ;
        RECT 1175.000 158.710 1175.600 158.850 ;
        RECT 1175.000 158.170 1175.140 158.710 ;
        RECT 1175.000 158.030 1175.600 158.170 ;
        RECT 1175.460 62.290 1175.600 158.030 ;
        RECT 1175.000 62.150 1175.600 62.290 ;
        RECT 1175.000 39.090 1175.140 62.150 ;
        RECT 109.580 38.770 109.840 39.090 ;
        RECT 1174.940 38.770 1175.200 39.090 ;
        RECT 109.640 2.400 109.780 38.770 ;
        RECT 109.430 -4.800 109.990 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1174.470 1207.200 1174.750 1207.480 ;
        RECT 1175.390 1207.200 1175.670 1207.480 ;
        RECT 1174.470 1110.640 1174.750 1110.920 ;
        RECT 1175.390 1110.640 1175.670 1110.920 ;
        RECT 1175.390 814.840 1175.670 815.120 ;
        RECT 1174.930 814.160 1175.210 814.440 ;
        RECT 1175.390 435.400 1175.670 435.680 ;
        RECT 1174.930 434.720 1175.210 435.000 ;
        RECT 109.570 39.640 109.850 39.920 ;
        RECT 1174.470 39.640 1174.750 39.920 ;
      LAYER met3 ;
        RECT 1174.445 1207.490 1174.775 1207.505 ;
        RECT 1175.365 1207.490 1175.695 1207.505 ;
        RECT 1174.445 1207.190 1175.695 1207.490 ;
        RECT 1174.445 1207.175 1174.775 1207.190 ;
        RECT 1175.365 1207.175 1175.695 1207.190 ;
        RECT 1174.445 1110.930 1174.775 1110.945 ;
        RECT 1175.365 1110.930 1175.695 1110.945 ;
        RECT 1174.445 1110.630 1175.695 1110.930 ;
        RECT 1174.445 1110.615 1174.775 1110.630 ;
        RECT 1175.365 1110.615 1175.695 1110.630 ;
        RECT 1175.365 815.130 1175.695 815.145 ;
        RECT 1175.150 814.815 1175.695 815.130 ;
        RECT 1175.150 814.465 1175.450 814.815 ;
        RECT 1174.905 814.150 1175.450 814.465 ;
        RECT 1174.905 814.135 1175.235 814.150 ;
        RECT 1175.365 435.690 1175.695 435.705 ;
        RECT 1175.150 435.375 1175.695 435.690 ;
        RECT 1175.150 435.025 1175.450 435.375 ;
        RECT 1174.905 434.710 1175.450 435.025 ;
        RECT 1174.905 434.695 1175.235 434.710 ;
        RECT 109.545 39.930 109.875 39.945 ;
        RECT 1174.445 39.930 1174.775 39.945 ;
        RECT 109.545 39.630 1174.775 39.930 ;
        RECT 109.545 39.615 109.875 39.630 ;
        RECT 1174.445 39.615 1174.775 39.630 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 0.300 ;
=======
      LAYER li1 ;
        RECT 1182.345 89.845 1182.515 137.955 ;
        RECT 1181.885 48.365 1182.055 62.815 ;
      LAYER mcon ;
        RECT 1182.345 137.785 1182.515 137.955 ;
        RECT 1181.885 62.645 1182.055 62.815 ;
      LAYER met1 ;
        RECT 1182.270 1559.820 1182.590 1559.880 ;
        RECT 1181.900 1559.680 1182.590 1559.820 ;
        RECT 1181.900 1559.540 1182.040 1559.680 ;
        RECT 1182.270 1559.620 1182.590 1559.680 ;
        RECT 1181.810 1559.280 1182.130 1559.540 ;
        RECT 1180.890 741.780 1181.210 741.840 ;
        RECT 1181.810 741.780 1182.130 741.840 ;
        RECT 1180.890 741.640 1182.130 741.780 ;
        RECT 1180.890 741.580 1181.210 741.640 ;
        RECT 1181.810 741.580 1182.130 741.640 ;
        RECT 1181.350 717.640 1181.670 717.700 ;
        RECT 1182.270 717.640 1182.590 717.700 ;
        RECT 1181.350 717.500 1182.590 717.640 ;
        RECT 1181.350 717.440 1181.670 717.500 ;
        RECT 1182.270 717.440 1182.590 717.500 ;
        RECT 1181.350 145.080 1181.670 145.140 ;
        RECT 1182.270 145.080 1182.590 145.140 ;
        RECT 1181.350 144.940 1182.590 145.080 ;
        RECT 1181.350 144.880 1181.670 144.940 ;
        RECT 1182.270 144.880 1182.590 144.940 ;
        RECT 1182.270 137.940 1182.590 138.000 ;
        RECT 1182.075 137.800 1182.590 137.940 ;
        RECT 1182.270 137.740 1182.590 137.800 ;
        RECT 1182.270 90.000 1182.590 90.060 ;
        RECT 1182.075 89.860 1182.590 90.000 ;
        RECT 1182.270 89.800 1182.590 89.860 ;
        RECT 1181.825 62.800 1182.115 62.845 ;
        RECT 1182.270 62.800 1182.590 62.860 ;
        RECT 1181.825 62.660 1182.590 62.800 ;
        RECT 1181.825 62.615 1182.115 62.660 ;
        RECT 1182.270 62.600 1182.590 62.660 ;
        RECT 1181.810 48.520 1182.130 48.580 ;
        RECT 1181.615 48.380 1182.130 48.520 ;
        RECT 1181.810 48.320 1182.130 48.380 ;
        RECT 133.470 39.340 133.790 39.400 ;
        RECT 1181.810 39.340 1182.130 39.400 ;
        RECT 133.470 39.200 1182.130 39.340 ;
        RECT 133.470 39.140 133.790 39.200 ;
        RECT 1181.810 39.140 1182.130 39.200 ;
      LAYER via ;
        RECT 1182.300 1559.620 1182.560 1559.880 ;
        RECT 1181.840 1559.280 1182.100 1559.540 ;
        RECT 1180.920 741.580 1181.180 741.840 ;
        RECT 1181.840 741.580 1182.100 741.840 ;
        RECT 1181.380 717.440 1181.640 717.700 ;
        RECT 1182.300 717.440 1182.560 717.700 ;
        RECT 1181.380 144.880 1181.640 145.140 ;
        RECT 1182.300 144.880 1182.560 145.140 ;
        RECT 1182.300 137.740 1182.560 138.000 ;
        RECT 1182.300 89.800 1182.560 90.060 ;
        RECT 1182.300 62.600 1182.560 62.860 ;
        RECT 1181.840 48.320 1182.100 48.580 ;
        RECT 133.500 39.140 133.760 39.400 ;
        RECT 1181.840 39.140 1182.100 39.400 ;
      LAYER met2 ;
        RECT 1185.970 1700.410 1186.250 1704.000 ;
        RECT 1185.120 1700.270 1186.250 1700.410 ;
        RECT 1185.120 1676.610 1185.260 1700.270 ;
        RECT 1185.970 1700.000 1186.250 1700.270 ;
        RECT 1182.360 1676.470 1185.260 1676.610 ;
        RECT 1182.360 1559.910 1182.500 1676.470 ;
        RECT 1182.300 1559.590 1182.560 1559.910 ;
        RECT 1181.840 1559.250 1182.100 1559.570 ;
        RECT 1181.900 1414.810 1182.040 1559.250 ;
        RECT 1181.440 1414.670 1182.040 1414.810 ;
        RECT 1181.440 1414.130 1181.580 1414.670 ;
        RECT 1181.440 1413.990 1182.040 1414.130 ;
        RECT 1181.900 1318.250 1182.040 1413.990 ;
        RECT 1181.440 1318.110 1182.040 1318.250 ;
        RECT 1181.440 1317.570 1181.580 1318.110 ;
        RECT 1181.440 1317.430 1182.040 1317.570 ;
        RECT 1181.900 1221.690 1182.040 1317.430 ;
        RECT 1181.440 1221.550 1182.040 1221.690 ;
        RECT 1181.440 1221.010 1181.580 1221.550 ;
        RECT 1181.440 1220.870 1182.040 1221.010 ;
        RECT 1181.900 1125.130 1182.040 1220.870 ;
        RECT 1181.440 1124.990 1182.040 1125.130 ;
        RECT 1181.440 1124.450 1181.580 1124.990 ;
        RECT 1181.440 1124.310 1182.040 1124.450 ;
        RECT 1181.900 1028.570 1182.040 1124.310 ;
        RECT 1181.440 1028.430 1182.040 1028.570 ;
        RECT 1181.440 1027.890 1181.580 1028.430 ;
        RECT 1181.440 1027.750 1182.040 1027.890 ;
        RECT 1181.900 932.010 1182.040 1027.750 ;
        RECT 1181.440 931.870 1182.040 932.010 ;
        RECT 1181.440 931.330 1181.580 931.870 ;
        RECT 1181.440 931.190 1182.040 931.330 ;
        RECT 1181.900 835.450 1182.040 931.190 ;
        RECT 1181.440 835.310 1182.040 835.450 ;
        RECT 1181.440 834.770 1181.580 835.310 ;
        RECT 1181.440 834.630 1182.040 834.770 ;
        RECT 1181.900 741.870 1182.040 834.630 ;
        RECT 1180.920 741.550 1181.180 741.870 ;
        RECT 1181.840 741.550 1182.100 741.870 ;
        RECT 1180.980 717.810 1181.120 741.550 ;
        RECT 1180.980 717.730 1181.580 717.810 ;
        RECT 1180.980 717.670 1181.640 717.730 ;
        RECT 1181.380 717.410 1181.640 717.670 ;
        RECT 1182.300 717.410 1182.560 717.730 ;
        RECT 1182.360 669.645 1182.500 717.410 ;
        RECT 1181.370 669.275 1181.650 669.645 ;
        RECT 1182.290 669.275 1182.570 669.645 ;
        RECT 1181.440 650.490 1181.580 669.275 ;
        RECT 1181.440 650.350 1182.040 650.490 ;
        RECT 1181.900 545.770 1182.040 650.350 ;
        RECT 1181.440 545.630 1182.040 545.770 ;
        RECT 1181.440 545.090 1181.580 545.630 ;
        RECT 1181.440 544.950 1182.040 545.090 ;
        RECT 1181.900 449.210 1182.040 544.950 ;
        RECT 1181.440 449.070 1182.040 449.210 ;
        RECT 1181.440 448.530 1181.580 449.070 ;
        RECT 1181.440 448.390 1182.040 448.530 ;
        RECT 1181.900 351.970 1182.040 448.390 ;
        RECT 1181.440 351.830 1182.040 351.970 ;
        RECT 1181.440 351.290 1181.580 351.830 ;
        RECT 1181.440 351.150 1182.040 351.290 ;
        RECT 1181.900 255.410 1182.040 351.150 ;
        RECT 1181.440 255.270 1182.040 255.410 ;
        RECT 1181.440 254.730 1181.580 255.270 ;
        RECT 1181.440 254.590 1182.040 254.730 ;
        RECT 1181.900 184.010 1182.040 254.590 ;
        RECT 1181.440 183.870 1182.040 184.010 ;
        RECT 1181.440 145.170 1181.580 183.870 ;
        RECT 1181.380 144.850 1181.640 145.170 ;
        RECT 1182.300 144.850 1182.560 145.170 ;
        RECT 1182.360 138.030 1182.500 144.850 ;
        RECT 1182.300 137.710 1182.560 138.030 ;
        RECT 1182.300 89.770 1182.560 90.090 ;
        RECT 1182.360 62.890 1182.500 89.770 ;
        RECT 1182.300 62.570 1182.560 62.890 ;
        RECT 1181.840 48.290 1182.100 48.610 ;
        RECT 1181.900 39.430 1182.040 48.290 ;
        RECT 133.500 39.110 133.760 39.430 ;
        RECT 1181.840 39.110 1182.100 39.430 ;
        RECT 133.560 2.400 133.700 39.110 ;
        RECT 133.350 -4.800 133.910 2.400 ;
      LAYER via2 ;
        RECT 1181.370 669.320 1181.650 669.600 ;
        RECT 1182.290 669.320 1182.570 669.600 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1181.345 724.690 1181.675 724.705 ;
        RECT 1182.265 724.690 1182.595 724.705 ;
        RECT 1181.345 724.390 1182.595 724.690 ;
        RECT 1181.345 724.375 1181.675 724.390 ;
        RECT 1182.265 724.375 1182.595 724.390 ;
        RECT 1181.345 628.810 1181.675 628.825 ;
        RECT 1181.345 628.495 1181.890 628.810 ;
        RECT 1181.590 628.145 1181.890 628.495 ;
        RECT 1181.345 627.830 1181.890 628.145 ;
        RECT 1181.345 627.815 1181.675 627.830 ;
        RECT 1180.885 470.370 1181.215 470.385 ;
        RECT 1180.885 470.070 1181.890 470.370 ;
        RECT 1180.885 470.055 1181.215 470.070 ;
        RECT 1180.885 469.010 1181.215 469.025 ;
        RECT 1181.590 469.010 1181.890 470.070 ;
        RECT 1180.885 468.710 1181.890 469.010 ;
        RECT 1180.885 468.695 1181.215 468.710 ;
        RECT 133.465 40.610 133.795 40.625 ;
        RECT 1181.345 40.610 1181.675 40.625 ;
        RECT 133.465 40.310 1181.675 40.610 ;
        RECT 133.465 40.295 133.795 40.310 ;
        RECT 1181.345 40.295 1181.675 40.310 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1181.345 669.610 1181.675 669.625 ;
        RECT 1182.265 669.610 1182.595 669.625 ;
        RECT 1181.345 669.310 1182.595 669.610 ;
        RECT 1181.345 669.295 1181.675 669.310 ;
        RECT 1182.265 669.295 1182.595 669.310 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 0.300 ;
=======
      LAYER met1 ;
        RECT 1187.790 717.640 1188.110 717.700 ;
        RECT 1188.710 717.640 1189.030 717.700 ;
        RECT 1187.790 717.500 1189.030 717.640 ;
        RECT 1187.790 717.440 1188.110 717.500 ;
        RECT 1188.710 717.440 1189.030 717.500 ;
        RECT 151.410 45.120 151.730 45.180 ;
        RECT 1187.790 45.120 1188.110 45.180 ;
        RECT 151.410 44.980 1188.110 45.120 ;
        RECT 151.410 44.920 151.730 44.980 ;
        RECT 1187.790 44.920 1188.110 44.980 ;
      LAYER via ;
        RECT 1187.820 717.440 1188.080 717.700 ;
        RECT 1188.740 717.440 1189.000 717.700 ;
        RECT 151.440 44.920 151.700 45.180 ;
        RECT 1187.820 44.920 1188.080 45.180 ;
      LAYER met2 ;
        RECT 1190.570 1700.410 1190.850 1704.000 ;
        RECT 1190.180 1700.270 1190.850 1700.410 ;
        RECT 1190.180 1684.770 1190.320 1700.270 ;
        RECT 1190.570 1700.000 1190.850 1700.270 ;
        RECT 1188.800 1684.630 1190.320 1684.770 ;
        RECT 1188.800 1582.770 1188.940 1684.630 ;
        RECT 1187.880 1582.630 1188.940 1582.770 ;
        RECT 1187.880 1558.970 1188.020 1582.630 ;
        RECT 1187.880 1558.830 1188.480 1558.970 ;
        RECT 1188.340 1414.810 1188.480 1558.830 ;
        RECT 1187.880 1414.670 1188.480 1414.810 ;
        RECT 1187.880 1414.130 1188.020 1414.670 ;
        RECT 1187.880 1413.990 1188.480 1414.130 ;
        RECT 1188.340 1318.250 1188.480 1413.990 ;
        RECT 1187.880 1318.110 1188.480 1318.250 ;
        RECT 1187.880 1317.570 1188.020 1318.110 ;
        RECT 1187.880 1317.430 1188.480 1317.570 ;
        RECT 1188.340 1221.690 1188.480 1317.430 ;
        RECT 1187.880 1221.550 1188.480 1221.690 ;
        RECT 1187.880 1221.010 1188.020 1221.550 ;
        RECT 1187.880 1220.870 1188.480 1221.010 ;
        RECT 1188.340 1125.130 1188.480 1220.870 ;
        RECT 1187.880 1124.990 1188.480 1125.130 ;
        RECT 1187.880 1124.450 1188.020 1124.990 ;
        RECT 1187.880 1124.310 1188.480 1124.450 ;
        RECT 1188.340 1028.570 1188.480 1124.310 ;
        RECT 1187.880 1028.430 1188.480 1028.570 ;
        RECT 1187.880 1027.890 1188.020 1028.430 ;
        RECT 1187.880 1027.750 1188.480 1027.890 ;
        RECT 1188.340 932.010 1188.480 1027.750 ;
        RECT 1187.880 931.870 1188.480 932.010 ;
        RECT 1187.880 931.330 1188.020 931.870 ;
        RECT 1187.880 931.190 1188.480 931.330 ;
        RECT 1188.340 835.450 1188.480 931.190 ;
        RECT 1187.880 835.310 1188.480 835.450 ;
        RECT 1187.880 834.770 1188.020 835.310 ;
        RECT 1187.880 834.630 1188.480 834.770 ;
        RECT 1188.340 738.890 1188.480 834.630 ;
        RECT 1188.340 738.750 1188.940 738.890 ;
        RECT 1188.800 717.925 1188.940 738.750 ;
        RECT 1187.810 717.555 1188.090 717.925 ;
        RECT 1188.730 717.555 1189.010 717.925 ;
        RECT 1187.820 717.410 1188.080 717.555 ;
        RECT 1188.740 717.410 1189.000 717.555 ;
        RECT 1188.800 669.645 1188.940 717.410 ;
        RECT 1187.810 669.275 1188.090 669.645 ;
        RECT 1188.730 669.275 1189.010 669.645 ;
        RECT 1187.880 650.490 1188.020 669.275 ;
        RECT 1187.880 650.350 1188.480 650.490 ;
        RECT 1188.340 545.770 1188.480 650.350 ;
        RECT 1187.880 545.630 1188.480 545.770 ;
        RECT 1187.880 545.090 1188.020 545.630 ;
        RECT 1187.880 544.950 1188.480 545.090 ;
        RECT 1188.340 449.210 1188.480 544.950 ;
        RECT 1187.880 449.070 1188.480 449.210 ;
        RECT 1187.880 448.530 1188.020 449.070 ;
        RECT 1187.880 448.390 1188.480 448.530 ;
        RECT 1188.340 351.970 1188.480 448.390 ;
        RECT 1187.880 351.830 1188.480 351.970 ;
        RECT 1187.880 351.290 1188.020 351.830 ;
        RECT 1187.880 351.150 1188.480 351.290 ;
        RECT 1188.340 255.410 1188.480 351.150 ;
        RECT 1187.880 255.270 1188.480 255.410 ;
        RECT 1187.880 254.730 1188.020 255.270 ;
        RECT 1187.880 254.590 1188.480 254.730 ;
        RECT 1188.340 158.850 1188.480 254.590 ;
        RECT 1187.880 158.710 1188.480 158.850 ;
        RECT 1187.880 158.170 1188.020 158.710 ;
        RECT 1187.880 158.030 1188.480 158.170 ;
        RECT 1188.340 62.290 1188.480 158.030 ;
        RECT 1187.880 62.150 1188.480 62.290 ;
        RECT 1187.880 45.210 1188.020 62.150 ;
        RECT 151.440 44.890 151.700 45.210 ;
        RECT 1187.820 44.890 1188.080 45.210 ;
        RECT 151.500 2.400 151.640 44.890 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 1187.810 717.600 1188.090 717.880 ;
        RECT 1188.730 717.600 1189.010 717.880 ;
        RECT 1187.810 669.320 1188.090 669.600 ;
        RECT 1188.730 669.320 1189.010 669.600 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 151.405 45.370 151.735 45.385 ;
        RECT 1187.785 45.370 1188.115 45.385 ;
        RECT 151.405 45.070 1188.115 45.370 ;
        RECT 151.405 45.055 151.735 45.070 ;
        RECT 1187.785 45.055 1188.115 45.070 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1187.785 717.890 1188.115 717.905 ;
        RECT 1188.705 717.890 1189.035 717.905 ;
        RECT 1187.785 717.590 1189.035 717.890 ;
        RECT 1187.785 717.575 1188.115 717.590 ;
        RECT 1188.705 717.575 1189.035 717.590 ;
        RECT 1187.785 669.610 1188.115 669.625 ;
        RECT 1188.705 669.610 1189.035 669.625 ;
        RECT 1187.785 669.310 1189.035 669.610 ;
        RECT 1187.785 669.295 1188.115 669.310 ;
        RECT 1188.705 669.295 1189.035 669.310 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 169.350 45.460 169.670 45.520 ;
        RECT 1194.230 45.460 1194.550 45.520 ;
        RECT 169.350 45.320 1194.550 45.460 ;
        RECT 169.350 45.260 169.670 45.320 ;
        RECT 1194.230 45.260 1194.550 45.320 ;
      LAYER via ;
        RECT 169.380 45.260 169.640 45.520 ;
        RECT 1194.260 45.260 1194.520 45.520 ;
      LAYER met2 ;
<<<<<<< HEAD
<<<<<<< HEAD
        RECT 169.230 -4.800 169.790 0.300 ;
=======
        RECT 1195.170 1700.410 1195.450 1704.000 ;
        RECT 1194.780 1700.270 1195.450 1700.410 ;
        RECT 1194.780 46.085 1194.920 1700.270 ;
        RECT 1195.170 1700.000 1195.450 1700.270 ;
        RECT 169.370 45.715 169.650 46.085 ;
        RECT 1194.710 45.715 1194.990 46.085 ;
        RECT 169.440 2.400 169.580 45.715 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 169.370 45.760 169.650 46.040 ;
        RECT 1194.710 45.760 1194.990 46.040 ;
      LAYER met3 ;
        RECT 169.345 46.050 169.675 46.065 ;
        RECT 1194.685 46.050 1195.015 46.065 ;
        RECT 169.345 45.750 1195.015 46.050 ;
        RECT 169.345 45.735 169.675 45.750 ;
        RECT 1194.685 45.735 1195.015 45.750 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1195.630 1700.410 1195.910 1704.000 ;
        RECT 1194.320 1700.270 1195.910 1700.410 ;
        RECT 1194.320 45.550 1194.460 1700.270 ;
        RECT 1195.630 1700.000 1195.910 1700.270 ;
        RECT 169.380 45.230 169.640 45.550 ;
        RECT 1194.260 45.230 1194.520 45.550 ;
        RECT 169.440 2.400 169.580 45.230 ;
        RECT 169.230 -4.800 169.790 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 0.300 ;
=======
      LAYER li1 ;
        RECT 1196.145 675.665 1196.315 717.655 ;
        RECT 1196.605 469.285 1196.775 517.395 ;
        RECT 1196.145 385.645 1196.315 427.635 ;
      LAYER mcon ;
        RECT 1196.145 717.485 1196.315 717.655 ;
        RECT 1196.605 517.225 1196.775 517.395 ;
        RECT 1196.145 427.465 1196.315 427.635 ;
      LAYER met1 ;
        RECT 1196.530 1558.940 1196.850 1559.200 ;
        RECT 1196.620 1558.520 1196.760 1558.940 ;
        RECT 1196.530 1558.260 1196.850 1558.520 ;
        RECT 1196.530 1462.380 1196.850 1462.640 ;
        RECT 1196.620 1461.960 1196.760 1462.380 ;
        RECT 1196.530 1461.700 1196.850 1461.960 ;
        RECT 1196.530 1365.820 1196.850 1366.080 ;
        RECT 1196.620 1365.400 1196.760 1365.820 ;
        RECT 1196.530 1365.140 1196.850 1365.400 ;
        RECT 1196.530 1269.260 1196.850 1269.520 ;
        RECT 1196.620 1268.840 1196.760 1269.260 ;
        RECT 1196.530 1268.580 1196.850 1268.840 ;
        RECT 1196.530 1172.700 1196.850 1172.960 ;
        RECT 1196.620 1172.280 1196.760 1172.700 ;
        RECT 1196.530 1172.020 1196.850 1172.280 ;
        RECT 1196.530 1076.140 1196.850 1076.400 ;
        RECT 1196.620 1075.720 1196.760 1076.140 ;
        RECT 1196.530 1075.460 1196.850 1075.720 ;
        RECT 1196.070 772.720 1196.390 772.780 ;
        RECT 1196.530 772.720 1196.850 772.780 ;
        RECT 1196.070 772.580 1196.850 772.720 ;
        RECT 1196.070 772.520 1196.390 772.580 ;
        RECT 1196.530 772.520 1196.850 772.580 ;
        RECT 1196.070 717.640 1196.390 717.700 ;
        RECT 1195.875 717.500 1196.390 717.640 ;
        RECT 1196.070 717.440 1196.390 717.500 ;
        RECT 1196.085 675.820 1196.375 675.865 ;
        RECT 1196.990 675.820 1197.310 675.880 ;
        RECT 1196.085 675.680 1197.310 675.820 ;
        RECT 1196.085 675.635 1196.375 675.680 ;
        RECT 1196.990 675.620 1197.310 675.680 ;
        RECT 1196.530 628.220 1196.850 628.280 ;
        RECT 1196.990 628.220 1197.310 628.280 ;
        RECT 1196.530 628.080 1197.310 628.220 ;
        RECT 1196.530 628.020 1196.850 628.080 ;
        RECT 1196.990 628.020 1197.310 628.080 ;
        RECT 1196.070 572.460 1196.390 572.520 ;
        RECT 1196.990 572.460 1197.310 572.520 ;
        RECT 1196.070 572.320 1197.310 572.460 ;
        RECT 1196.070 572.260 1196.390 572.320 ;
        RECT 1196.990 572.260 1197.310 572.320 ;
        RECT 1196.530 517.380 1196.850 517.440 ;
        RECT 1196.335 517.240 1196.850 517.380 ;
        RECT 1196.530 517.180 1196.850 517.240 ;
        RECT 1196.530 469.440 1196.850 469.500 ;
        RECT 1196.335 469.300 1196.850 469.440 ;
        RECT 1196.530 469.240 1196.850 469.300 ;
        RECT 1196.070 427.620 1196.390 427.680 ;
        RECT 1195.875 427.480 1196.390 427.620 ;
        RECT 1196.070 427.420 1196.390 427.480 ;
        RECT 1196.085 385.800 1196.375 385.845 ;
        RECT 1196.990 385.800 1197.310 385.860 ;
        RECT 1196.085 385.660 1197.310 385.800 ;
        RECT 1196.085 385.615 1196.375 385.660 ;
        RECT 1196.990 385.600 1197.310 385.660 ;
        RECT 1196.530 338.200 1196.850 338.260 ;
        RECT 1196.990 338.200 1197.310 338.260 ;
        RECT 1196.530 338.060 1197.310 338.200 ;
        RECT 1196.530 338.000 1196.850 338.060 ;
        RECT 1196.990 338.000 1197.310 338.060 ;
        RECT 1196.070 158.820 1196.390 159.080 ;
        RECT 1196.160 158.000 1196.300 158.820 ;
        RECT 1196.530 158.000 1196.850 158.060 ;
        RECT 1196.160 157.860 1196.850 158.000 ;
        RECT 1196.530 157.800 1196.850 157.860 ;
        RECT 1196.530 137.740 1196.850 138.000 ;
        RECT 1196.620 137.320 1196.760 137.740 ;
        RECT 1196.530 137.060 1196.850 137.320 ;
      LAYER via ;
        RECT 1196.560 1558.940 1196.820 1559.200 ;
        RECT 1196.560 1558.260 1196.820 1558.520 ;
        RECT 1196.560 1462.380 1196.820 1462.640 ;
        RECT 1196.560 1461.700 1196.820 1461.960 ;
        RECT 1196.560 1365.820 1196.820 1366.080 ;
        RECT 1196.560 1365.140 1196.820 1365.400 ;
        RECT 1196.560 1269.260 1196.820 1269.520 ;
        RECT 1196.560 1268.580 1196.820 1268.840 ;
        RECT 1196.560 1172.700 1196.820 1172.960 ;
        RECT 1196.560 1172.020 1196.820 1172.280 ;
        RECT 1196.560 1076.140 1196.820 1076.400 ;
        RECT 1196.560 1075.460 1196.820 1075.720 ;
        RECT 1196.100 772.520 1196.360 772.780 ;
        RECT 1196.560 772.520 1196.820 772.780 ;
        RECT 1196.100 717.440 1196.360 717.700 ;
        RECT 1197.020 675.620 1197.280 675.880 ;
        RECT 1196.560 628.020 1196.820 628.280 ;
        RECT 1197.020 628.020 1197.280 628.280 ;
        RECT 1196.100 572.260 1196.360 572.520 ;
        RECT 1197.020 572.260 1197.280 572.520 ;
        RECT 1196.560 517.180 1196.820 517.440 ;
        RECT 1196.560 469.240 1196.820 469.500 ;
        RECT 1196.100 427.420 1196.360 427.680 ;
        RECT 1197.020 385.600 1197.280 385.860 ;
        RECT 1196.560 338.000 1196.820 338.260 ;
        RECT 1197.020 338.000 1197.280 338.260 ;
        RECT 1196.100 158.820 1196.360 159.080 ;
        RECT 1196.560 157.800 1196.820 158.060 ;
        RECT 1196.560 137.740 1196.820 138.000 ;
        RECT 1196.560 137.060 1196.820 137.320 ;
=======
      LAYER met1 ;
        RECT 1194.690 1678.140 1195.010 1678.200 ;
        RECT 1199.290 1678.140 1199.610 1678.200 ;
        RECT 1194.690 1678.000 1199.610 1678.140 ;
        RECT 1194.690 1677.940 1195.010 1678.000 ;
        RECT 1199.290 1677.940 1199.610 1678.000 ;
        RECT 192.350 51.580 192.670 51.640 ;
        RECT 1194.690 51.580 1195.010 51.640 ;
        RECT 192.350 51.440 1195.010 51.580 ;
        RECT 192.350 51.380 192.670 51.440 ;
        RECT 1194.690 51.380 1195.010 51.440 ;
        RECT 186.830 15.200 187.150 15.260 ;
        RECT 192.350 15.200 192.670 15.260 ;
        RECT 186.830 15.060 192.670 15.200 ;
        RECT 186.830 15.000 187.150 15.060 ;
        RECT 192.350 15.000 192.670 15.060 ;
      LAYER via ;
        RECT 1194.720 1677.940 1194.980 1678.200 ;
        RECT 1199.320 1677.940 1199.580 1678.200 ;
        RECT 192.380 51.380 192.640 51.640 ;
        RECT 1194.720 51.380 1194.980 51.640 ;
        RECT 186.860 15.000 187.120 15.260 ;
        RECT 192.380 15.000 192.640 15.260 ;
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1200.230 1700.410 1200.510 1704.000 ;
        RECT 1199.380 1700.270 1200.510 1700.410 ;
        RECT 1199.380 1678.230 1199.520 1700.270 ;
        RECT 1200.230 1700.000 1200.510 1700.270 ;
        RECT 1194.720 1677.910 1194.980 1678.230 ;
        RECT 1199.320 1677.910 1199.580 1678.230 ;
        RECT 1194.780 51.670 1194.920 1677.910 ;
        RECT 192.380 51.350 192.640 51.670 ;
        RECT 1194.720 51.350 1194.980 51.670 ;
        RECT 192.440 15.290 192.580 51.350 ;
        RECT 186.860 14.970 187.120 15.290 ;
        RECT 192.380 14.970 192.640 15.290 ;
        RECT 186.920 2.400 187.060 14.970 ;
        RECT 186.710 -4.800 187.270 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1196.550 435.400 1196.830 435.680 ;
        RECT 1196.090 434.720 1196.370 435.000 ;
        RECT 186.850 51.200 187.130 51.480 ;
        RECT 1196.550 51.200 1196.830 51.480 ;
      LAYER met3 ;
        RECT 1196.525 435.690 1196.855 435.705 ;
        RECT 1196.310 435.375 1196.855 435.690 ;
        RECT 1196.310 435.025 1196.610 435.375 ;
        RECT 1196.065 434.710 1196.610 435.025 ;
        RECT 1196.065 434.695 1196.395 434.710 ;
        RECT 186.825 51.490 187.155 51.505 ;
        RECT 1196.525 51.490 1196.855 51.505 ;
        RECT 186.825 51.190 1196.855 51.490 ;
        RECT 186.825 51.175 187.155 51.190 ;
        RECT 1196.525 51.175 1196.855 51.190 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 204.650 -4.800 205.210 0.300 ;
=======
        RECT 1204.830 1700.410 1205.110 1704.000 ;
        RECT 1203.980 1700.270 1205.110 1700.410 ;
        RECT 1203.980 1678.140 1204.120 1700.270 ;
        RECT 1204.830 1700.000 1205.110 1700.270 ;
        RECT 1201.220 1678.000 1204.120 1678.140 ;
        RECT 1201.220 52.205 1201.360 1678.000 ;
        RECT 204.790 51.835 205.070 52.205 ;
        RECT 1201.150 51.835 1201.430 52.205 ;
        RECT 204.860 2.400 205.000 51.835 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 204.790 51.880 205.070 52.160 ;
        RECT 1201.150 51.880 1201.430 52.160 ;
      LAYER met3 ;
        RECT 204.765 52.170 205.095 52.185 ;
        RECT 1201.125 52.170 1201.455 52.185 ;
        RECT 204.765 51.870 1201.455 52.170 ;
        RECT 204.765 51.855 205.095 51.870 ;
        RECT 1201.125 51.855 1201.455 51.870 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1201.130 1678.140 1201.450 1678.200 ;
        RECT 1203.890 1678.140 1204.210 1678.200 ;
        RECT 1201.130 1678.000 1204.210 1678.140 ;
        RECT 1201.130 1677.940 1201.450 1678.000 ;
        RECT 1203.890 1677.940 1204.210 1678.000 ;
        RECT 206.610 51.920 206.930 51.980 ;
        RECT 1201.130 51.920 1201.450 51.980 ;
        RECT 206.610 51.780 1201.450 51.920 ;
        RECT 206.610 51.720 206.930 51.780 ;
        RECT 1201.130 51.720 1201.450 51.780 ;
      LAYER via ;
        RECT 1201.160 1677.940 1201.420 1678.200 ;
        RECT 1203.920 1677.940 1204.180 1678.200 ;
        RECT 206.640 51.720 206.900 51.980 ;
        RECT 1201.160 51.720 1201.420 51.980 ;
      LAYER met2 ;
        RECT 1205.290 1700.410 1205.570 1704.000 ;
        RECT 1203.980 1700.270 1205.570 1700.410 ;
        RECT 1203.980 1678.230 1204.120 1700.270 ;
        RECT 1205.290 1700.000 1205.570 1700.270 ;
        RECT 1201.160 1677.910 1201.420 1678.230 ;
        RECT 1203.920 1677.910 1204.180 1678.230 ;
        RECT 1201.220 52.010 1201.360 1677.910 ;
        RECT 206.640 51.690 206.900 52.010 ;
        RECT 1201.160 51.690 1201.420 52.010 ;
        RECT 206.700 17.410 206.840 51.690 ;
        RECT 204.860 17.270 206.840 17.410 ;
        RECT 204.860 2.400 205.000 17.270 ;
        RECT 204.650 -4.800 205.210 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 0.300 ;
=======
      LAYER met1 ;
        RECT 227.310 52.260 227.630 52.320 ;
        RECT 1208.030 52.260 1208.350 52.320 ;
        RECT 227.310 52.120 1208.350 52.260 ;
        RECT 227.310 52.060 227.630 52.120 ;
        RECT 1208.030 52.060 1208.350 52.120 ;
        RECT 222.710 15.200 223.030 15.260 ;
        RECT 227.310 15.200 227.630 15.260 ;
        RECT 222.710 15.060 227.630 15.200 ;
        RECT 222.710 15.000 223.030 15.060 ;
        RECT 227.310 15.000 227.630 15.060 ;
      LAYER via ;
        RECT 227.340 52.060 227.600 52.320 ;
        RECT 1208.060 52.060 1208.320 52.320 ;
        RECT 222.740 15.000 223.000 15.260 ;
        RECT 227.340 15.000 227.600 15.260 ;
      LAYER met2 ;
        RECT 1209.890 1700.410 1210.170 1704.000 ;
        RECT 1209.040 1700.270 1210.170 1700.410 ;
        RECT 1209.040 1678.140 1209.180 1700.270 ;
        RECT 1209.890 1700.000 1210.170 1700.270 ;
        RECT 1208.120 1678.000 1209.180 1678.140 ;
        RECT 1208.120 52.350 1208.260 1678.000 ;
        RECT 227.340 52.030 227.600 52.350 ;
        RECT 1208.060 52.030 1208.320 52.350 ;
        RECT 227.400 15.290 227.540 52.030 ;
        RECT 222.740 14.970 223.000 15.290 ;
        RECT 227.340 14.970 227.600 15.290 ;
        RECT 222.800 2.400 222.940 14.970 ;
        RECT 222.590 -4.800 223.150 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 227.330 52.560 227.610 52.840 ;
        RECT 1209.430 52.560 1209.710 52.840 ;
      LAYER met3 ;
        RECT 227.305 52.850 227.635 52.865 ;
        RECT 1209.405 52.850 1209.735 52.865 ;
        RECT 227.305 52.550 1209.735 52.850 ;
        RECT 227.305 52.535 227.635 52.550 ;
        RECT 1209.405 52.535 1209.735 52.550 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 37.980 20.630 38.040 ;
        RECT 1153.290 37.980 1153.610 38.040 ;
        RECT 20.310 37.840 1153.610 37.980 ;
        RECT 20.310 37.780 20.630 37.840 ;
        RECT 1153.290 37.780 1153.610 37.840 ;
      LAYER via ;
        RECT 20.340 37.780 20.600 38.040 ;
        RECT 1153.320 37.780 1153.580 38.040 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 20.190 -4.800 20.750 0.300 ;
=======
        RECT 1155.150 1700.410 1155.430 1704.000 ;
        RECT 1154.300 1700.270 1155.430 1700.410 ;
        RECT 1154.300 1661.650 1154.440 1700.270 ;
        RECT 1155.150 1700.000 1155.430 1700.270 ;
        RECT 1153.380 1661.510 1154.440 1661.650 ;
        RECT 1153.380 38.070 1153.520 1661.510 ;
        RECT 20.340 37.750 20.600 38.070 ;
        RECT 1153.320 37.750 1153.580 38.070 ;
        RECT 20.400 2.400 20.540 37.750 ;
        RECT 20.190 -4.800 20.750 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 20.330 37.600 20.610 37.880 ;
        RECT 1154.230 37.600 1154.510 37.880 ;
      LAYER met3 ;
        RECT 20.305 37.890 20.635 37.905 ;
        RECT 1154.205 37.890 1154.535 37.905 ;
        RECT 20.305 37.590 1154.535 37.890 ;
        RECT 20.305 37.575 20.635 37.590 ;
        RECT 1154.205 37.575 1154.535 37.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 44.110 -4.800 44.670 0.300 ;
=======
        RECT 1161.590 1700.410 1161.870 1704.000 ;
        RECT 1160.740 1700.270 1161.870 1700.410 ;
        RECT 1160.740 44.725 1160.880 1700.270 ;
        RECT 1161.590 1700.000 1161.870 1700.270 ;
        RECT 44.250 44.355 44.530 44.725 ;
        RECT 1160.670 44.355 1160.950 44.725 ;
        RECT 44.320 2.400 44.460 44.355 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 44.250 44.400 44.530 44.680 ;
        RECT 1160.670 44.400 1160.950 44.680 ;
      LAYER met3 ;
        RECT 44.225 44.690 44.555 44.705 ;
        RECT 1160.645 44.690 1160.975 44.705 ;
        RECT 44.225 44.390 1160.975 44.690 ;
        RECT 44.225 44.375 44.555 44.390 ;
        RECT 1160.645 44.375 1160.975 44.390 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1159.730 1679.840 1160.050 1679.900 ;
        RECT 1161.570 1679.840 1161.890 1679.900 ;
        RECT 1159.730 1679.700 1161.890 1679.840 ;
        RECT 1159.730 1679.640 1160.050 1679.700 ;
        RECT 1161.570 1679.640 1161.890 1679.700 ;
        RECT 44.230 44.780 44.550 44.840 ;
        RECT 1159.730 44.780 1160.050 44.840 ;
        RECT 44.230 44.640 1160.050 44.780 ;
        RECT 44.230 44.580 44.550 44.640 ;
        RECT 1159.730 44.580 1160.050 44.640 ;
      LAYER via ;
        RECT 1159.760 1679.640 1160.020 1679.900 ;
        RECT 1161.600 1679.640 1161.860 1679.900 ;
        RECT 44.260 44.580 44.520 44.840 ;
        RECT 1159.760 44.580 1160.020 44.840 ;
      LAYER met2 ;
        RECT 1161.590 1700.000 1161.870 1704.000 ;
        RECT 1161.660 1679.930 1161.800 1700.000 ;
        RECT 1159.760 1679.610 1160.020 1679.930 ;
        RECT 1161.600 1679.610 1161.860 1679.930 ;
        RECT 1159.820 44.870 1159.960 1679.610 ;
        RECT 44.260 44.550 44.520 44.870 ;
        RECT 1159.760 44.550 1160.020 44.870 ;
        RECT 44.320 2.400 44.460 44.550 ;
        RECT 44.110 -4.800 44.670 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 248.010 52.600 248.330 52.660 ;
        RECT 1215.850 52.600 1216.170 52.660 ;
        RECT 248.010 52.460 1216.170 52.600 ;
        RECT 248.010 52.400 248.330 52.460 ;
        RECT 1215.850 52.400 1216.170 52.460 ;
      LAYER via ;
        RECT 248.040 52.400 248.300 52.660 ;
        RECT 1215.880 52.400 1216.140 52.660 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 246.510 -4.800 247.070 0.300 ;
=======
        RECT 1216.330 1700.410 1216.610 1704.000 ;
        RECT 1215.940 1700.270 1216.610 1700.410 ;
        RECT 1215.940 52.690 1216.080 1700.270 ;
        RECT 1216.330 1700.000 1216.610 1700.270 ;
        RECT 248.040 52.370 248.300 52.690 ;
        RECT 1215.880 52.370 1216.140 52.690 ;
        RECT 248.100 17.410 248.240 52.370 ;
        RECT 246.720 17.270 248.240 17.410 ;
        RECT 246.720 2.400 246.860 17.270 ;
        RECT 246.510 -4.800 247.070 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 248.030 53.240 248.310 53.520 ;
        RECT 1215.870 53.240 1216.150 53.520 ;
      LAYER met3 ;
        RECT 248.005 53.530 248.335 53.545 ;
        RECT 1215.845 53.530 1216.175 53.545 ;
        RECT 248.005 53.230 1216.175 53.530 ;
        RECT 248.005 53.215 248.335 53.230 ;
        RECT 1215.845 53.215 1216.175 53.230 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1221.370 1695.480 1221.690 1695.540 ;
        RECT 1223.210 1695.480 1223.530 1695.540 ;
        RECT 1221.370 1695.340 1223.530 1695.480 ;
        RECT 1221.370 1695.280 1221.690 1695.340 ;
        RECT 1223.210 1695.280 1223.530 1695.340 ;
        RECT 268.710 52.940 269.030 53.000 ;
        RECT 1223.210 52.940 1223.530 53.000 ;
        RECT 268.710 52.800 1223.530 52.940 ;
        RECT 268.710 52.740 269.030 52.800 ;
        RECT 1223.210 52.740 1223.530 52.800 ;
        RECT 264.110 17.580 264.430 17.640 ;
        RECT 268.710 17.580 269.030 17.640 ;
        RECT 264.110 17.440 269.030 17.580 ;
        RECT 264.110 17.380 264.430 17.440 ;
        RECT 268.710 17.380 269.030 17.440 ;
      LAYER via ;
        RECT 1221.400 1695.280 1221.660 1695.540 ;
        RECT 1223.240 1695.280 1223.500 1695.540 ;
        RECT 268.740 52.740 269.000 53.000 ;
        RECT 1223.240 52.740 1223.500 53.000 ;
        RECT 264.140 17.380 264.400 17.640 ;
        RECT 268.740 17.380 269.000 17.640 ;
      LAYER met2 ;
        RECT 1221.390 1700.000 1221.670 1704.000 ;
        RECT 1221.460 1695.570 1221.600 1700.000 ;
        RECT 1221.400 1695.250 1221.660 1695.570 ;
        RECT 1223.240 1695.250 1223.500 1695.570 ;
        RECT 1223.300 53.030 1223.440 1695.250 ;
        RECT 268.740 52.710 269.000 53.030 ;
        RECT 1223.240 52.710 1223.500 53.030 ;
        RECT 268.800 17.670 268.940 52.710 ;
        RECT 264.140 17.350 264.400 17.670 ;
        RECT 268.740 17.350 269.000 17.670 ;
        RECT 264.200 2.400 264.340 17.350 ;
        RECT 263.990 -4.800 264.550 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 268.730 53.920 269.010 54.200 ;
        RECT 1215.410 53.920 1215.690 54.200 ;
      LAYER met3 ;
        RECT 268.705 54.210 269.035 54.225 ;
        RECT 1215.385 54.210 1215.715 54.225 ;
        RECT 268.705 53.910 1215.715 54.210 ;
        RECT 268.705 53.895 269.035 53.910 ;
        RECT 1215.385 53.895 1215.715 53.910 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1222.290 1678.140 1222.610 1678.200 ;
        RECT 1224.590 1678.140 1224.910 1678.200 ;
        RECT 1222.290 1678.000 1224.910 1678.140 ;
        RECT 1222.290 1677.940 1222.610 1678.000 ;
        RECT 1224.590 1677.940 1224.910 1678.000 ;
      LAYER via ;
        RECT 1222.320 1677.940 1222.580 1678.200 ;
        RECT 1224.620 1677.940 1224.880 1678.200 ;
=======
      LAYER li1 ;
        RECT 1225.125 1090.125 1225.295 1138.575 ;
        RECT 1225.585 1041.845 1225.755 1063.095 ;
        RECT 1225.585 951.405 1225.755 993.395 ;
        RECT 1224.665 848.725 1224.835 856.035 ;
        RECT 1225.125 572.645 1225.295 620.755 ;
      LAYER mcon ;
        RECT 1225.125 1138.405 1225.295 1138.575 ;
        RECT 1225.585 1062.925 1225.755 1063.095 ;
        RECT 1225.585 993.225 1225.755 993.395 ;
        RECT 1224.665 855.865 1224.835 856.035 ;
        RECT 1225.125 620.585 1225.295 620.755 ;
      LAYER met1 ;
        RECT 1224.590 1469.720 1224.910 1469.780 ;
        RECT 1225.510 1469.720 1225.830 1469.780 ;
        RECT 1224.590 1469.580 1225.830 1469.720 ;
        RECT 1224.590 1469.520 1224.910 1469.580 ;
        RECT 1225.510 1469.520 1225.830 1469.580 ;
        RECT 1224.590 1401.040 1224.910 1401.100 ;
        RECT 1225.050 1401.040 1225.370 1401.100 ;
        RECT 1224.590 1400.900 1225.370 1401.040 ;
        RECT 1224.590 1400.840 1224.910 1400.900 ;
        RECT 1225.050 1400.840 1225.370 1400.900 ;
        RECT 1224.590 1304.480 1224.910 1304.540 ;
        RECT 1225.050 1304.480 1225.370 1304.540 ;
        RECT 1224.590 1304.340 1225.370 1304.480 ;
        RECT 1224.590 1304.280 1224.910 1304.340 ;
        RECT 1225.050 1304.280 1225.370 1304.340 ;
        RECT 1225.050 1270.140 1225.370 1270.200 ;
        RECT 1224.680 1270.000 1225.370 1270.140 ;
        RECT 1224.680 1269.520 1224.820 1270.000 ;
        RECT 1225.050 1269.940 1225.370 1270.000 ;
        RECT 1224.590 1269.260 1224.910 1269.520 ;
        RECT 1224.590 1207.580 1224.910 1207.640 ;
        RECT 1225.050 1207.580 1225.370 1207.640 ;
        RECT 1224.590 1207.440 1225.370 1207.580 ;
        RECT 1224.590 1207.380 1224.910 1207.440 ;
        RECT 1225.050 1207.380 1225.370 1207.440 ;
        RECT 1225.050 1173.380 1225.370 1173.640 ;
        RECT 1225.140 1172.960 1225.280 1173.380 ;
        RECT 1225.050 1172.700 1225.370 1172.960 ;
        RECT 1225.050 1138.560 1225.370 1138.620 ;
        RECT 1224.855 1138.420 1225.370 1138.560 ;
        RECT 1225.050 1138.360 1225.370 1138.420 ;
        RECT 1225.065 1090.280 1225.355 1090.325 ;
        RECT 1225.510 1090.280 1225.830 1090.340 ;
        RECT 1225.065 1090.140 1225.830 1090.280 ;
        RECT 1225.065 1090.095 1225.355 1090.140 ;
        RECT 1225.510 1090.080 1225.830 1090.140 ;
        RECT 1225.510 1063.080 1225.830 1063.140 ;
        RECT 1225.315 1062.940 1225.830 1063.080 ;
        RECT 1225.510 1062.880 1225.830 1062.940 ;
        RECT 1224.130 1042.000 1224.450 1042.060 ;
        RECT 1225.525 1042.000 1225.815 1042.045 ;
        RECT 1224.130 1041.860 1225.815 1042.000 ;
        RECT 1224.130 1041.800 1224.450 1041.860 ;
        RECT 1225.525 1041.815 1225.815 1041.860 ;
        RECT 1224.130 1041.320 1224.450 1041.380 ;
        RECT 1225.510 1041.320 1225.830 1041.380 ;
        RECT 1224.130 1041.180 1225.830 1041.320 ;
        RECT 1224.130 1041.120 1224.450 1041.180 ;
        RECT 1225.510 1041.120 1225.830 1041.180 ;
        RECT 1225.510 993.380 1225.830 993.440 ;
        RECT 1225.315 993.240 1225.830 993.380 ;
        RECT 1225.510 993.180 1225.830 993.240 ;
        RECT 1225.510 951.560 1225.830 951.620 ;
        RECT 1225.315 951.420 1225.830 951.560 ;
        RECT 1225.510 951.360 1225.830 951.420 ;
        RECT 1224.605 856.020 1224.895 856.065 ;
        RECT 1225.050 856.020 1225.370 856.080 ;
        RECT 1224.605 855.880 1225.370 856.020 ;
        RECT 1224.605 855.835 1224.895 855.880 ;
        RECT 1225.050 855.820 1225.370 855.880 ;
        RECT 1224.590 848.880 1224.910 848.940 ;
        RECT 1224.395 848.740 1224.910 848.880 ;
        RECT 1224.590 848.680 1224.910 848.740 ;
        RECT 1224.590 807.540 1224.910 807.800 ;
        RECT 1224.680 806.720 1224.820 807.540 ;
        RECT 1225.050 806.720 1225.370 806.780 ;
        RECT 1224.680 806.580 1225.370 806.720 ;
        RECT 1225.050 806.520 1225.370 806.580 ;
        RECT 1224.590 734.780 1224.910 735.040 ;
        RECT 1224.680 734.360 1224.820 734.780 ;
        RECT 1224.590 734.100 1224.910 734.360 ;
        RECT 1225.050 620.740 1225.370 620.800 ;
        RECT 1224.855 620.600 1225.370 620.740 ;
        RECT 1225.050 620.540 1225.370 620.600 ;
        RECT 1225.050 572.800 1225.370 572.860 ;
        RECT 1224.855 572.660 1225.370 572.800 ;
        RECT 1225.050 572.600 1225.370 572.660 ;
        RECT 1225.050 476.580 1225.370 476.640 ;
        RECT 1224.680 476.440 1225.370 476.580 ;
        RECT 1224.680 476.300 1224.820 476.440 ;
        RECT 1225.050 476.380 1225.370 476.440 ;
        RECT 1224.590 476.040 1224.910 476.300 ;
        RECT 1225.050 145.080 1225.370 145.140 ;
        RECT 1225.510 145.080 1225.830 145.140 ;
        RECT 1225.050 144.940 1225.830 145.080 ;
        RECT 1225.050 144.880 1225.370 144.940 ;
        RECT 1225.510 144.880 1225.830 144.940 ;
        RECT 1224.590 96.800 1224.910 96.860 ;
        RECT 1225.050 96.800 1225.370 96.860 ;
        RECT 1224.590 96.660 1225.370 96.800 ;
        RECT 1224.590 96.600 1224.910 96.660 ;
        RECT 1225.050 96.600 1225.370 96.660 ;
        RECT 282.050 53.280 282.370 53.340 ;
        RECT 1224.590 53.280 1224.910 53.340 ;
        RECT 282.050 53.140 1224.910 53.280 ;
        RECT 282.050 53.080 282.370 53.140 ;
        RECT 1224.590 53.080 1224.910 53.140 ;
      LAYER via ;
        RECT 1224.620 1469.520 1224.880 1469.780 ;
        RECT 1225.540 1469.520 1225.800 1469.780 ;
        RECT 1224.620 1400.840 1224.880 1401.100 ;
        RECT 1225.080 1400.840 1225.340 1401.100 ;
        RECT 1224.620 1304.280 1224.880 1304.540 ;
        RECT 1225.080 1304.280 1225.340 1304.540 ;
        RECT 1225.080 1269.940 1225.340 1270.200 ;
        RECT 1224.620 1269.260 1224.880 1269.520 ;
        RECT 1224.620 1207.380 1224.880 1207.640 ;
        RECT 1225.080 1207.380 1225.340 1207.640 ;
        RECT 1225.080 1173.380 1225.340 1173.640 ;
        RECT 1225.080 1172.700 1225.340 1172.960 ;
        RECT 1225.080 1138.360 1225.340 1138.620 ;
        RECT 1225.540 1090.080 1225.800 1090.340 ;
        RECT 1225.540 1062.880 1225.800 1063.140 ;
        RECT 1224.160 1041.800 1224.420 1042.060 ;
        RECT 1224.160 1041.120 1224.420 1041.380 ;
        RECT 1225.540 1041.120 1225.800 1041.380 ;
        RECT 1225.540 993.180 1225.800 993.440 ;
        RECT 1225.540 951.360 1225.800 951.620 ;
        RECT 1225.080 855.820 1225.340 856.080 ;
        RECT 1224.620 848.680 1224.880 848.940 ;
        RECT 1224.620 807.540 1224.880 807.800 ;
        RECT 1225.080 806.520 1225.340 806.780 ;
        RECT 1224.620 734.780 1224.880 735.040 ;
        RECT 1224.620 734.100 1224.880 734.360 ;
        RECT 1225.080 620.540 1225.340 620.800 ;
        RECT 1225.080 572.600 1225.340 572.860 ;
        RECT 1225.080 476.380 1225.340 476.640 ;
        RECT 1224.620 476.040 1224.880 476.300 ;
        RECT 1225.080 144.880 1225.340 145.140 ;
        RECT 1225.540 144.880 1225.800 145.140 ;
        RECT 1224.620 96.600 1224.880 96.860 ;
        RECT 1225.080 96.600 1225.340 96.860 ;
        RECT 282.080 53.080 282.340 53.340 ;
        RECT 1224.620 53.080 1224.880 53.340 ;
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1225.990 1700.410 1226.270 1704.000 ;
        RECT 1225.600 1700.270 1226.270 1700.410 ;
        RECT 1225.600 1690.890 1225.740 1700.270 ;
        RECT 1225.990 1700.000 1226.270 1700.270 ;
        RECT 1225.140 1690.750 1225.740 1690.890 ;
        RECT 1225.140 1563.050 1225.280 1690.750 ;
        RECT 1224.680 1562.910 1225.280 1563.050 ;
        RECT 1224.680 1521.570 1224.820 1562.910 ;
        RECT 1224.680 1521.430 1225.740 1521.570 ;
        RECT 1225.600 1469.810 1225.740 1521.430 ;
        RECT 1224.620 1469.490 1224.880 1469.810 ;
        RECT 1225.540 1469.490 1225.800 1469.810 ;
        RECT 1224.680 1401.130 1224.820 1469.490 ;
        RECT 1224.620 1400.810 1224.880 1401.130 ;
        RECT 1225.080 1400.810 1225.340 1401.130 ;
        RECT 1225.140 1369.930 1225.280 1400.810 ;
        RECT 1224.680 1369.790 1225.280 1369.930 ;
        RECT 1224.680 1304.570 1224.820 1369.790 ;
        RECT 1224.620 1304.250 1224.880 1304.570 ;
        RECT 1225.080 1304.250 1225.340 1304.570 ;
        RECT 1225.140 1270.230 1225.280 1304.250 ;
        RECT 1225.080 1269.910 1225.340 1270.230 ;
        RECT 1224.620 1269.230 1224.880 1269.550 ;
        RECT 1224.680 1207.670 1224.820 1269.230 ;
        RECT 1224.620 1207.350 1224.880 1207.670 ;
        RECT 1225.080 1207.350 1225.340 1207.670 ;
        RECT 1225.140 1173.670 1225.280 1207.350 ;
        RECT 1225.080 1173.350 1225.340 1173.670 ;
        RECT 1225.080 1172.670 1225.340 1172.990 ;
        RECT 1225.140 1138.650 1225.280 1172.670 ;
        RECT 1225.080 1138.330 1225.340 1138.650 ;
        RECT 1225.540 1090.050 1225.800 1090.370 ;
        RECT 1225.600 1063.170 1225.740 1090.050 ;
        RECT 1225.540 1062.850 1225.800 1063.170 ;
        RECT 1224.160 1041.770 1224.420 1042.090 ;
        RECT 1224.220 1041.410 1224.360 1041.770 ;
        RECT 1224.160 1041.090 1224.420 1041.410 ;
        RECT 1225.540 1041.090 1225.800 1041.410 ;
        RECT 1225.600 993.470 1225.740 1041.090 ;
        RECT 1225.540 993.150 1225.800 993.470 ;
        RECT 1225.540 951.330 1225.800 951.650 ;
        RECT 1225.600 910.250 1225.740 951.330 ;
        RECT 1225.140 910.110 1225.740 910.250 ;
        RECT 1225.140 856.110 1225.280 910.110 ;
        RECT 1225.080 855.790 1225.340 856.110 ;
        RECT 1224.620 848.650 1224.880 848.970 ;
        RECT 1224.680 807.830 1224.820 848.650 ;
        RECT 1224.620 807.510 1224.880 807.830 ;
        RECT 1225.080 806.490 1225.340 806.810 ;
        RECT 1225.140 759.290 1225.280 806.490 ;
        RECT 1224.680 759.150 1225.280 759.290 ;
        RECT 1224.680 735.070 1224.820 759.150 ;
        RECT 1224.620 734.750 1224.880 735.070 ;
        RECT 1224.620 734.070 1224.880 734.390 ;
        RECT 1224.680 685.850 1224.820 734.070 ;
        RECT 1224.680 685.710 1225.280 685.850 ;
        RECT 1225.140 620.830 1225.280 685.710 ;
        RECT 1225.080 620.510 1225.340 620.830 ;
        RECT 1225.080 572.570 1225.340 572.890 ;
        RECT 1225.140 476.670 1225.280 572.570 ;
        RECT 1225.080 476.350 1225.340 476.670 ;
        RECT 1224.620 476.010 1224.880 476.330 ;
        RECT 1224.680 448.530 1224.820 476.010 ;
        RECT 1224.680 448.390 1225.280 448.530 ;
        RECT 1225.140 303.690 1225.280 448.390 ;
        RECT 1224.680 303.550 1225.280 303.690 ;
        RECT 1224.680 266.290 1224.820 303.550 ;
        RECT 1224.680 266.150 1225.740 266.290 ;
        RECT 1225.600 254.730 1225.740 266.150 ;
        RECT 1225.140 254.590 1225.740 254.730 ;
        RECT 1225.140 193.020 1225.280 254.590 ;
        RECT 1225.140 192.880 1225.740 193.020 ;
        RECT 1225.600 145.170 1225.740 192.880 ;
        RECT 1225.080 144.850 1225.340 145.170 ;
        RECT 1225.540 144.850 1225.800 145.170 ;
        RECT 1225.140 96.890 1225.280 144.850 ;
        RECT 1224.620 96.570 1224.880 96.890 ;
        RECT 1225.080 96.570 1225.340 96.890 ;
        RECT 1224.680 53.370 1224.820 96.570 ;
        RECT 282.080 53.050 282.340 53.370 ;
        RECT 1224.620 53.050 1224.880 53.370 ;
        RECT 282.140 2.400 282.280 53.050 ;
        RECT 281.930 -4.800 282.490 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 282.070 54.600 282.350 54.880 ;
        RECT 1222.310 54.600 1222.590 54.880 ;
      LAYER met3 ;
        RECT 282.045 54.890 282.375 54.905 ;
        RECT 1222.285 54.890 1222.615 54.905 ;
        RECT 282.045 54.590 1222.615 54.890 ;
        RECT 282.045 54.575 282.375 54.590 ;
        RECT 1222.285 54.575 1222.615 54.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 0.300 ;
=======
      LAYER met1 ;
        RECT 303.210 53.620 303.530 53.680 ;
        RECT 1229.650 53.620 1229.970 53.680 ;
        RECT 303.210 53.480 1229.970 53.620 ;
        RECT 303.210 53.420 303.530 53.480 ;
        RECT 1229.650 53.420 1229.970 53.480 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 299.990 16.760 303.530 16.900 ;
        RECT 299.990 16.700 300.310 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 303.240 53.420 303.500 53.680 ;
        RECT 1229.680 53.420 1229.940 53.680 ;
        RECT 300.020 16.700 300.280 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 1231.050 1700.410 1231.330 1704.000 ;
        RECT 1229.740 1700.270 1231.330 1700.410 ;
        RECT 1229.740 53.710 1229.880 1700.270 ;
        RECT 1231.050 1700.000 1231.330 1700.270 ;
        RECT 303.240 53.390 303.500 53.710 ;
        RECT 1229.680 53.390 1229.940 53.710 ;
        RECT 303.300 16.990 303.440 53.390 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 0.300 ;
=======
      LAYER met1 ;
        RECT 323.910 53.960 324.230 54.020 ;
        RECT 1236.090 53.960 1236.410 54.020 ;
        RECT 323.910 53.820 1236.410 53.960 ;
        RECT 323.910 53.760 324.230 53.820 ;
        RECT 1236.090 53.760 1236.410 53.820 ;
        RECT 317.930 16.900 318.250 16.960 ;
        RECT 323.910 16.900 324.230 16.960 ;
        RECT 317.930 16.760 324.230 16.900 ;
        RECT 317.930 16.700 318.250 16.760 ;
        RECT 323.910 16.700 324.230 16.760 ;
      LAYER via ;
        RECT 323.940 53.760 324.200 54.020 ;
        RECT 1236.120 53.760 1236.380 54.020 ;
        RECT 317.960 16.700 318.220 16.960 ;
        RECT 323.940 16.700 324.200 16.960 ;
      LAYER met2 ;
        RECT 1235.650 1700.410 1235.930 1704.000 ;
        RECT 1235.650 1700.270 1236.320 1700.410 ;
        RECT 1235.650 1700.000 1235.930 1700.270 ;
        RECT 1236.180 54.050 1236.320 1700.270 ;
        RECT 323.940 53.730 324.200 54.050 ;
        RECT 1236.120 53.730 1236.380 54.050 ;
        RECT 324.000 16.990 324.140 53.730 ;
        RECT 317.960 16.670 318.220 16.990 ;
        RECT 323.940 16.670 324.200 16.990 ;
        RECT 318.020 2.400 318.160 16.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 0.300 ;
=======
      LAYER li1 ;
        RECT 1237.085 1400.205 1237.255 1414.655 ;
        RECT 1237.545 517.905 1237.715 545.955 ;
        RECT 1237.545 434.605 1237.715 469.115 ;
        RECT 1238.005 258.825 1238.175 305.575 ;
        RECT 1238.005 183.685 1238.175 227.715 ;
      LAYER mcon ;
        RECT 1237.085 1414.485 1237.255 1414.655 ;
        RECT 1237.545 545.785 1237.715 545.955 ;
        RECT 1237.545 468.945 1237.715 469.115 ;
        RECT 1238.005 305.405 1238.175 305.575 ;
        RECT 1238.005 227.545 1238.175 227.715 ;
      LAYER met1 ;
        RECT 1237.930 1559.620 1238.250 1559.880 ;
        RECT 1238.020 1559.200 1238.160 1559.620 ;
        RECT 1237.930 1558.940 1238.250 1559.200 ;
        RECT 1237.025 1414.640 1237.315 1414.685 ;
        RECT 1237.470 1414.640 1237.790 1414.700 ;
        RECT 1237.025 1414.500 1237.790 1414.640 ;
        RECT 1237.025 1414.455 1237.315 1414.500 ;
        RECT 1237.470 1414.440 1237.790 1414.500 ;
        RECT 1237.010 1400.360 1237.330 1400.420 ;
        RECT 1236.815 1400.220 1237.330 1400.360 ;
        RECT 1237.010 1400.160 1237.330 1400.220 ;
        RECT 1237.010 1345.620 1237.330 1345.680 ;
        RECT 1237.930 1345.620 1238.250 1345.680 ;
        RECT 1237.010 1345.480 1238.250 1345.620 ;
        RECT 1237.010 1345.420 1237.330 1345.480 ;
        RECT 1237.930 1345.420 1238.250 1345.480 ;
        RECT 1237.470 1283.400 1237.790 1283.460 ;
        RECT 1238.390 1283.400 1238.710 1283.460 ;
        RECT 1237.470 1283.260 1238.710 1283.400 ;
        RECT 1237.470 1283.200 1237.790 1283.260 ;
        RECT 1238.390 1283.200 1238.710 1283.260 ;
        RECT 1237.930 1159.300 1238.250 1159.360 ;
        RECT 1238.390 1159.300 1238.710 1159.360 ;
        RECT 1237.930 1159.160 1238.710 1159.300 ;
        RECT 1237.930 1159.100 1238.250 1159.160 ;
        RECT 1238.390 1159.100 1238.710 1159.160 ;
        RECT 1237.470 1076.680 1237.790 1076.740 ;
        RECT 1237.470 1076.540 1238.160 1076.680 ;
        RECT 1237.470 1076.480 1237.790 1076.540 ;
        RECT 1238.020 1076.400 1238.160 1076.540 ;
        RECT 1237.930 1076.140 1238.250 1076.400 ;
        RECT 1237.470 724.440 1237.790 724.500 ;
        RECT 1238.390 724.440 1238.710 724.500 ;
        RECT 1237.470 724.300 1238.710 724.440 ;
        RECT 1237.470 724.240 1237.790 724.300 ;
        RECT 1238.390 724.240 1238.710 724.300 ;
        RECT 1237.470 572.800 1237.790 572.860 ;
        RECT 1237.930 572.800 1238.250 572.860 ;
        RECT 1237.470 572.660 1238.250 572.800 ;
        RECT 1237.470 572.600 1237.790 572.660 ;
        RECT 1237.930 572.600 1238.250 572.660 ;
        RECT 1237.470 545.940 1237.790 546.000 ;
        RECT 1237.275 545.800 1237.790 545.940 ;
        RECT 1237.470 545.740 1237.790 545.800 ;
        RECT 1237.470 518.060 1237.790 518.120 ;
        RECT 1237.275 517.920 1237.790 518.060 ;
        RECT 1237.470 517.860 1237.790 517.920 ;
        RECT 1237.010 517.380 1237.330 517.440 ;
        RECT 1237.470 517.380 1237.790 517.440 ;
        RECT 1237.010 517.240 1237.790 517.380 ;
        RECT 1237.010 517.180 1237.330 517.240 ;
        RECT 1237.470 517.180 1237.790 517.240 ;
        RECT 1237.470 469.100 1237.790 469.160 ;
        RECT 1237.275 468.960 1237.790 469.100 ;
        RECT 1237.470 468.900 1237.790 468.960 ;
        RECT 1237.485 434.760 1237.775 434.805 ;
        RECT 1237.930 434.760 1238.250 434.820 ;
        RECT 1237.485 434.620 1238.250 434.760 ;
        RECT 1237.485 434.575 1237.775 434.620 ;
        RECT 1237.930 434.560 1238.250 434.620 ;
        RECT 1237.930 305.560 1238.250 305.620 ;
        RECT 1237.735 305.420 1238.250 305.560 ;
        RECT 1237.930 305.360 1238.250 305.420 ;
        RECT 1237.470 258.980 1237.790 259.040 ;
        RECT 1237.945 258.980 1238.235 259.025 ;
        RECT 1237.470 258.840 1238.235 258.980 ;
        RECT 1237.470 258.780 1237.790 258.840 ;
        RECT 1237.945 258.795 1238.235 258.840 ;
        RECT 1237.930 227.700 1238.250 227.760 ;
        RECT 1237.735 227.560 1238.250 227.700 ;
        RECT 1237.930 227.500 1238.250 227.560 ;
        RECT 1237.930 183.840 1238.250 183.900 ;
        RECT 1237.735 183.700 1238.250 183.840 ;
        RECT 1237.930 183.640 1238.250 183.700 ;
        RECT 1237.930 159.020 1238.250 159.080 ;
        RECT 1237.560 158.880 1238.250 159.020 ;
        RECT 1237.560 158.740 1237.700 158.880 ;
        RECT 1237.930 158.820 1238.250 158.880 ;
        RECT 1237.470 158.480 1237.790 158.740 ;
        RECT 337.710 52.260 338.030 52.320 ;
        RECT 1237.470 52.260 1237.790 52.320 ;
        RECT 337.710 52.120 1237.790 52.260 ;
        RECT 337.710 52.060 338.030 52.120 ;
        RECT 1237.470 52.060 1237.790 52.120 ;
      LAYER via ;
        RECT 1237.960 1559.620 1238.220 1559.880 ;
        RECT 1237.960 1558.940 1238.220 1559.200 ;
        RECT 1237.500 1414.440 1237.760 1414.700 ;
        RECT 1237.040 1400.160 1237.300 1400.420 ;
        RECT 1237.040 1345.420 1237.300 1345.680 ;
        RECT 1237.960 1345.420 1238.220 1345.680 ;
        RECT 1237.500 1283.200 1237.760 1283.460 ;
        RECT 1238.420 1283.200 1238.680 1283.460 ;
        RECT 1237.960 1159.100 1238.220 1159.360 ;
        RECT 1238.420 1159.100 1238.680 1159.360 ;
        RECT 1237.500 1076.480 1237.760 1076.740 ;
        RECT 1237.960 1076.140 1238.220 1076.400 ;
        RECT 1237.500 724.240 1237.760 724.500 ;
        RECT 1238.420 724.240 1238.680 724.500 ;
        RECT 1237.500 572.600 1237.760 572.860 ;
        RECT 1237.960 572.600 1238.220 572.860 ;
        RECT 1237.500 545.740 1237.760 546.000 ;
        RECT 1237.500 517.860 1237.760 518.120 ;
        RECT 1237.040 517.180 1237.300 517.440 ;
        RECT 1237.500 517.180 1237.760 517.440 ;
        RECT 1237.500 468.900 1237.760 469.160 ;
        RECT 1237.960 434.560 1238.220 434.820 ;
        RECT 1237.960 305.360 1238.220 305.620 ;
        RECT 1237.500 258.780 1237.760 259.040 ;
        RECT 1237.960 227.500 1238.220 227.760 ;
        RECT 1237.960 183.640 1238.220 183.900 ;
        RECT 1237.960 158.820 1238.220 159.080 ;
        RECT 1237.500 158.480 1237.760 158.740 ;
        RECT 337.740 52.060 338.000 52.320 ;
        RECT 1237.500 52.060 1237.760 52.320 ;
      LAYER met2 ;
        RECT 1240.250 1700.410 1240.530 1704.000 ;
        RECT 1239.860 1700.270 1240.530 1700.410 ;
        RECT 1239.860 1677.970 1240.000 1700.270 ;
        RECT 1240.250 1700.000 1240.530 1700.270 ;
        RECT 1238.020 1677.830 1240.000 1677.970 ;
        RECT 1238.020 1559.910 1238.160 1677.830 ;
        RECT 1237.960 1559.590 1238.220 1559.910 ;
        RECT 1237.960 1558.910 1238.220 1559.230 ;
        RECT 1238.020 1463.090 1238.160 1558.910 ;
        RECT 1237.560 1462.950 1238.160 1463.090 ;
        RECT 1237.560 1462.410 1237.700 1462.950 ;
        RECT 1237.560 1462.270 1238.160 1462.410 ;
        RECT 1238.020 1442.010 1238.160 1462.270 ;
        RECT 1237.560 1441.870 1238.160 1442.010 ;
        RECT 1237.560 1414.730 1237.700 1441.870 ;
        RECT 1237.500 1414.410 1237.760 1414.730 ;
        RECT 1237.040 1400.130 1237.300 1400.450 ;
        RECT 1237.100 1345.710 1237.240 1400.130 ;
        RECT 1237.040 1345.390 1237.300 1345.710 ;
        RECT 1237.960 1345.390 1238.220 1345.710 ;
        RECT 1238.020 1314.170 1238.160 1345.390 ;
        RECT 1237.560 1314.030 1238.160 1314.170 ;
        RECT 1237.560 1283.490 1237.700 1314.030 ;
        RECT 1237.500 1283.170 1237.760 1283.490 ;
        RECT 1238.420 1283.170 1238.680 1283.490 ;
        RECT 1238.480 1159.390 1238.620 1283.170 ;
        RECT 1237.960 1159.070 1238.220 1159.390 ;
        RECT 1238.420 1159.070 1238.680 1159.390 ;
        RECT 1238.020 1104.050 1238.160 1159.070 ;
        RECT 1237.560 1103.910 1238.160 1104.050 ;
        RECT 1237.560 1076.770 1237.700 1103.910 ;
        RECT 1237.500 1076.450 1237.760 1076.770 ;
        RECT 1237.960 1076.110 1238.220 1076.430 ;
        RECT 1238.020 835.450 1238.160 1076.110 ;
        RECT 1237.560 835.310 1238.160 835.450 ;
        RECT 1237.560 834.770 1237.700 835.310 ;
        RECT 1237.560 834.630 1238.160 834.770 ;
        RECT 1238.020 773.685 1238.160 834.630 ;
        RECT 1237.950 773.315 1238.230 773.685 ;
        RECT 1237.950 772.635 1238.230 773.005 ;
        RECT 1238.020 738.890 1238.160 772.635 ;
        RECT 1238.020 738.750 1238.620 738.890 ;
        RECT 1238.480 724.725 1238.620 738.750 ;
        RECT 1237.490 724.355 1237.770 724.725 ;
        RECT 1238.410 724.355 1238.690 724.725 ;
        RECT 1237.500 724.210 1237.760 724.355 ;
        RECT 1238.420 724.210 1238.680 724.355 ;
        RECT 1238.480 699.450 1238.620 724.210 ;
        RECT 1238.020 699.310 1238.620 699.450 ;
        RECT 1238.020 628.845 1238.160 699.310 ;
        RECT 1237.950 628.475 1238.230 628.845 ;
        RECT 1237.950 627.795 1238.230 628.165 ;
        RECT 1238.020 572.890 1238.160 627.795 ;
        RECT 1237.500 572.570 1237.760 572.890 ;
        RECT 1237.960 572.570 1238.220 572.890 ;
        RECT 1237.560 546.030 1237.700 572.570 ;
        RECT 1237.500 545.710 1237.760 546.030 ;
        RECT 1237.500 517.830 1237.760 518.150 ;
        RECT 1237.560 517.470 1237.700 517.830 ;
        RECT 1237.040 517.150 1237.300 517.470 ;
        RECT 1237.500 517.150 1237.760 517.470 ;
        RECT 1237.100 475.730 1237.240 517.150 ;
        RECT 1237.100 475.590 1237.700 475.730 ;
        RECT 1237.560 469.190 1237.700 475.590 ;
        RECT 1237.500 468.870 1237.760 469.190 ;
        RECT 1237.960 434.530 1238.220 434.850 ;
        RECT 1238.020 305.650 1238.160 434.530 ;
        RECT 1237.960 305.330 1238.220 305.650 ;
        RECT 1237.500 258.750 1237.760 259.070 ;
        RECT 1237.560 235.010 1237.700 258.750 ;
        RECT 1237.560 234.870 1238.160 235.010 ;
        RECT 1238.020 227.790 1238.160 234.870 ;
        RECT 1237.960 227.470 1238.220 227.790 ;
        RECT 1237.960 183.610 1238.220 183.930 ;
        RECT 1238.020 159.110 1238.160 183.610 ;
        RECT 1237.960 158.790 1238.220 159.110 ;
        RECT 1237.500 158.450 1237.760 158.770 ;
        RECT 1237.560 52.350 1237.700 158.450 ;
        RECT 337.740 52.030 338.000 52.350 ;
        RECT 1237.500 52.030 1237.760 52.350 ;
        RECT 337.800 17.410 337.940 52.030 ;
        RECT 335.960 17.270 337.940 17.410 ;
        RECT 335.960 2.400 336.100 17.270 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 1237.950 773.360 1238.230 773.640 ;
        RECT 1237.950 772.680 1238.230 772.960 ;
        RECT 1237.490 724.400 1237.770 724.680 ;
        RECT 1238.410 724.400 1238.690 724.680 ;
        RECT 1237.950 628.520 1238.230 628.800 ;
        RECT 1237.950 627.840 1238.230 628.120 ;
      LAYER met3 ;
        RECT 1237.925 773.650 1238.255 773.665 ;
        RECT 1237.710 773.335 1238.255 773.650 ;
        RECT 1237.710 772.985 1238.010 773.335 ;
        RECT 1237.710 772.670 1238.255 772.985 ;
        RECT 1237.925 772.655 1238.255 772.670 ;
        RECT 1237.465 724.690 1237.795 724.705 ;
        RECT 1238.385 724.690 1238.715 724.705 ;
        RECT 1237.465 724.390 1238.715 724.690 ;
        RECT 1237.465 724.375 1237.795 724.390 ;
        RECT 1238.385 724.375 1238.715 724.390 ;
        RECT 1237.925 628.810 1238.255 628.825 ;
        RECT 1237.710 628.495 1238.255 628.810 ;
        RECT 1237.710 628.145 1238.010 628.495 ;
        RECT 1237.710 627.830 1238.255 628.145 ;
        RECT 1237.925 627.815 1238.255 627.830 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1236.550 1669.640 1236.870 1669.700 ;
        RECT 1239.310 1669.640 1239.630 1669.700 ;
        RECT 1236.550 1669.500 1239.630 1669.640 ;
        RECT 1236.550 1669.440 1236.870 1669.500 ;
        RECT 1239.310 1669.440 1239.630 1669.500 ;
        RECT 337.710 1631.900 338.030 1631.960 ;
        RECT 1236.550 1631.900 1236.870 1631.960 ;
        RECT 337.710 1631.760 1236.870 1631.900 ;
        RECT 337.710 1631.700 338.030 1631.760 ;
        RECT 1236.550 1631.700 1236.870 1631.760 ;
      LAYER via ;
        RECT 1236.580 1669.440 1236.840 1669.700 ;
        RECT 1239.340 1669.440 1239.600 1669.700 ;
        RECT 337.740 1631.700 338.000 1631.960 ;
        RECT 1236.580 1631.700 1236.840 1631.960 ;
      LAYER met2 ;
        RECT 1240.710 1700.410 1240.990 1704.000 ;
        RECT 1239.400 1700.270 1240.990 1700.410 ;
        RECT 1239.400 1669.730 1239.540 1700.270 ;
        RECT 1240.710 1700.000 1240.990 1700.270 ;
        RECT 1236.580 1669.410 1236.840 1669.730 ;
        RECT 1239.340 1669.410 1239.600 1669.730 ;
        RECT 1236.640 1631.990 1236.780 1669.410 ;
        RECT 337.740 1631.670 338.000 1631.990 ;
        RECT 1236.580 1631.670 1236.840 1631.990 ;
        RECT 337.800 3.130 337.940 1631.670 ;
        RECT 335.960 2.990 337.940 3.130 ;
        RECT 335.960 2.400 336.100 2.990 ;
        RECT 335.750 -4.800 336.310 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 0.300 ;
=======
      LAYER met1 ;
        RECT 1244.830 1628.840 1245.150 1628.900 ;
        RECT 1245.290 1628.840 1245.610 1628.900 ;
        RECT 1244.830 1628.700 1245.610 1628.840 ;
        RECT 1244.830 1628.640 1245.150 1628.700 ;
        RECT 1245.290 1628.640 1245.610 1628.700 ;
        RECT 358.410 1576.480 358.730 1576.540 ;
        RECT 1244.830 1576.480 1245.150 1576.540 ;
        RECT 358.410 1576.340 1245.150 1576.480 ;
        RECT 358.410 1576.280 358.730 1576.340 ;
        RECT 1244.830 1576.280 1245.150 1576.340 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 358.410 16.900 358.730 16.960 ;
        RECT 353.350 16.760 358.730 16.900 ;
        RECT 353.350 16.700 353.670 16.760 ;
        RECT 358.410 16.700 358.730 16.760 ;
      LAYER via ;
        RECT 1244.860 1628.640 1245.120 1628.900 ;
        RECT 1245.320 1628.640 1245.580 1628.900 ;
        RECT 358.440 1576.280 358.700 1576.540 ;
        RECT 1244.860 1576.280 1245.120 1576.540 ;
        RECT 353.380 16.700 353.640 16.960 ;
        RECT 358.440 16.700 358.700 16.960 ;
      LAYER met2 ;
        RECT 1245.310 1700.000 1245.590 1704.000 ;
        RECT 1245.380 1628.930 1245.520 1700.000 ;
        RECT 1244.860 1628.610 1245.120 1628.930 ;
        RECT 1245.320 1628.610 1245.580 1628.930 ;
        RECT 1244.920 1576.570 1245.060 1628.610 ;
        RECT 358.440 1576.250 358.700 1576.570 ;
        RECT 1244.860 1576.250 1245.120 1576.570 ;
        RECT 358.500 16.990 358.640 1576.250 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 358.440 16.670 358.700 16.990 ;
        RECT 353.440 2.400 353.580 16.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 0.300 ;
=======
      LAYER li1 ;
        RECT 1250.425 1666.085 1250.595 1679.175 ;
      LAYER mcon ;
        RECT 1250.425 1679.005 1250.595 1679.175 ;
      LAYER met1 ;
        RECT 1250.350 1679.160 1250.670 1679.220 ;
        RECT 1250.155 1679.020 1250.670 1679.160 ;
        RECT 1250.350 1678.960 1250.670 1679.020 ;
        RECT 1250.350 1666.240 1250.670 1666.300 ;
        RECT 1250.155 1666.100 1250.670 1666.240 ;
        RECT 1250.350 1666.040 1250.670 1666.100 ;
        RECT 372.210 1535.340 372.530 1535.400 ;
        RECT 1250.350 1535.340 1250.670 1535.400 ;
        RECT 372.210 1535.200 1250.670 1535.340 ;
        RECT 372.210 1535.140 372.530 1535.200 ;
        RECT 1250.350 1535.140 1250.670 1535.200 ;
        RECT 371.290 2.960 371.610 3.020 ;
        RECT 372.210 2.960 372.530 3.020 ;
        RECT 371.290 2.820 372.530 2.960 ;
        RECT 371.290 2.760 371.610 2.820 ;
        RECT 372.210 2.760 372.530 2.820 ;
      LAYER via ;
        RECT 1250.380 1678.960 1250.640 1679.220 ;
        RECT 1250.380 1666.040 1250.640 1666.300 ;
        RECT 372.240 1535.140 372.500 1535.400 ;
        RECT 1250.380 1535.140 1250.640 1535.400 ;
        RECT 371.320 2.760 371.580 3.020 ;
        RECT 372.240 2.760 372.500 3.020 ;
      LAYER met2 ;
        RECT 1250.370 1700.000 1250.650 1704.000 ;
        RECT 1250.440 1679.250 1250.580 1700.000 ;
        RECT 1250.380 1678.930 1250.640 1679.250 ;
        RECT 1250.380 1666.010 1250.640 1666.330 ;
        RECT 1250.440 1535.430 1250.580 1666.010 ;
        RECT 372.240 1535.110 372.500 1535.430 ;
        RECT 1250.380 1535.110 1250.640 1535.430 ;
        RECT 372.300 3.050 372.440 1535.110 ;
        RECT 371.320 2.730 371.580 3.050 ;
        RECT 372.240 2.730 372.500 3.050 ;
        RECT 371.380 2.400 371.520 2.730 ;
        RECT 371.170 -4.800 371.730 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1248.070 1428.200 1248.350 1428.480 ;
        RECT 1250.830 1428.200 1251.110 1428.480 ;
        RECT 1250.370 1014.080 1250.650 1014.360 ;
        RECT 1250.830 1013.400 1251.110 1013.680 ;
        RECT 1250.370 773.360 1250.650 773.640 ;
        RECT 1249.910 772.680 1250.190 772.960 ;
        RECT 1249.910 435.400 1250.190 435.680 ;
        RECT 1249.910 434.720 1250.190 435.000 ;
      LAYER met3 ;
        RECT 1248.045 1428.490 1248.375 1428.505 ;
        RECT 1250.805 1428.490 1251.135 1428.505 ;
        RECT 1248.045 1428.190 1251.135 1428.490 ;
        RECT 1248.045 1428.175 1248.375 1428.190 ;
        RECT 1250.805 1428.175 1251.135 1428.190 ;
        RECT 1250.345 1014.370 1250.675 1014.385 ;
        RECT 1250.345 1014.055 1250.890 1014.370 ;
        RECT 1250.590 1013.705 1250.890 1014.055 ;
        RECT 1250.590 1013.390 1251.135 1013.705 ;
        RECT 1250.805 1013.375 1251.135 1013.390 ;
        RECT 1250.345 773.650 1250.675 773.665 ;
        RECT 1249.670 773.350 1250.675 773.650 ;
        RECT 1249.670 772.985 1249.970 773.350 ;
        RECT 1250.345 773.335 1250.675 773.350 ;
        RECT 1249.670 772.670 1250.215 772.985 ;
        RECT 1249.885 772.655 1250.215 772.670 ;
        RECT 1249.885 435.690 1250.215 435.705 ;
        RECT 1249.670 435.375 1250.215 435.690 ;
        RECT 1249.670 435.025 1249.970 435.375 ;
        RECT 1249.670 434.710 1250.215 435.025 ;
        RECT 1249.885 434.695 1250.215 434.710 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 0.300 ;
=======
      LAYER li1 ;
        RECT 1251.345 1538.925 1251.515 1587.035 ;
        RECT 1251.345 1386.945 1251.515 1414.995 ;
        RECT 1251.345 1297.185 1251.515 1345.295 ;
        RECT 1251.345 1104.065 1251.515 1140.955 ;
        RECT 1251.805 565.845 1251.975 590.155 ;
        RECT 1251.345 331.245 1251.515 379.355 ;
        RECT 1251.345 59.585 1251.515 96.475 ;
      LAYER mcon ;
        RECT 1251.345 1586.865 1251.515 1587.035 ;
        RECT 1251.345 1414.825 1251.515 1414.995 ;
        RECT 1251.345 1345.125 1251.515 1345.295 ;
        RECT 1251.345 1140.785 1251.515 1140.955 ;
        RECT 1251.805 589.985 1251.975 590.155 ;
        RECT 1251.345 379.185 1251.515 379.355 ;
        RECT 1251.345 96.305 1251.515 96.475 ;
      LAYER met1 ;
        RECT 1251.270 1587.020 1251.590 1587.080 ;
        RECT 1251.075 1586.880 1251.590 1587.020 ;
        RECT 1251.270 1586.820 1251.590 1586.880 ;
        RECT 1251.285 1539.080 1251.575 1539.125 ;
        RECT 1251.730 1539.080 1252.050 1539.140 ;
        RECT 1251.285 1538.940 1252.050 1539.080 ;
        RECT 1251.285 1538.895 1251.575 1538.940 ;
        RECT 1251.730 1538.880 1252.050 1538.940 ;
        RECT 1251.270 1414.980 1251.590 1415.040 ;
        RECT 1251.075 1414.840 1251.590 1414.980 ;
        RECT 1251.270 1414.780 1251.590 1414.840 ;
        RECT 1251.270 1387.100 1251.590 1387.160 ;
        RECT 1251.075 1386.960 1251.590 1387.100 ;
        RECT 1251.270 1386.900 1251.590 1386.960 ;
        RECT 1251.270 1345.280 1251.590 1345.340 ;
        RECT 1251.075 1345.140 1251.590 1345.280 ;
        RECT 1251.270 1345.080 1251.590 1345.140 ;
        RECT 1251.285 1297.340 1251.575 1297.385 ;
        RECT 1252.190 1297.340 1252.510 1297.400 ;
        RECT 1251.285 1297.200 1252.510 1297.340 ;
        RECT 1251.285 1297.155 1251.575 1297.200 ;
        RECT 1252.190 1297.140 1252.510 1297.200 ;
        RECT 1251.270 1249.060 1251.590 1249.120 ;
        RECT 1252.190 1249.060 1252.510 1249.120 ;
        RECT 1251.270 1248.920 1252.510 1249.060 ;
        RECT 1251.270 1248.860 1251.590 1248.920 ;
        RECT 1252.190 1248.860 1252.510 1248.920 ;
        RECT 1251.270 1207.380 1251.590 1207.640 ;
        RECT 1251.360 1207.240 1251.500 1207.380 ;
        RECT 1251.730 1207.240 1252.050 1207.300 ;
        RECT 1251.360 1207.100 1252.050 1207.240 ;
        RECT 1251.730 1207.040 1252.050 1207.100 ;
        RECT 1251.270 1152.500 1251.590 1152.560 ;
        RECT 1252.190 1152.500 1252.510 1152.560 ;
        RECT 1251.270 1152.360 1252.510 1152.500 ;
        RECT 1251.270 1152.300 1251.590 1152.360 ;
        RECT 1252.190 1152.300 1252.510 1152.360 ;
        RECT 1251.270 1140.940 1251.590 1141.000 ;
        RECT 1251.075 1140.800 1251.590 1140.940 ;
        RECT 1251.270 1140.740 1251.590 1140.800 ;
        RECT 1251.285 1104.220 1251.575 1104.265 ;
        RECT 1252.190 1104.220 1252.510 1104.280 ;
        RECT 1251.285 1104.080 1252.510 1104.220 ;
        RECT 1251.285 1104.035 1251.575 1104.080 ;
        RECT 1252.190 1104.020 1252.510 1104.080 ;
        RECT 1252.190 1097.080 1252.510 1097.140 ;
        RECT 1253.110 1097.080 1253.430 1097.140 ;
        RECT 1252.190 1096.940 1253.430 1097.080 ;
        RECT 1252.190 1096.880 1252.510 1096.940 ;
        RECT 1253.110 1096.880 1253.430 1096.940 ;
        RECT 1251.730 1014.800 1252.050 1014.860 ;
        RECT 1251.360 1014.660 1252.050 1014.800 ;
        RECT 1251.360 1014.520 1251.500 1014.660 ;
        RECT 1251.730 1014.600 1252.050 1014.660 ;
        RECT 1251.270 1014.260 1251.590 1014.520 ;
        RECT 1251.270 979.920 1251.590 980.180 ;
        RECT 1251.360 979.500 1251.500 979.920 ;
        RECT 1251.270 979.240 1251.590 979.500 ;
        RECT 1251.270 931.640 1251.590 931.900 ;
        RECT 1251.360 931.160 1251.500 931.640 ;
        RECT 1251.730 931.160 1252.050 931.220 ;
        RECT 1251.360 931.020 1252.050 931.160 ;
        RECT 1251.730 930.960 1252.050 931.020 ;
        RECT 1251.270 869.620 1251.590 869.680 ;
        RECT 1252.190 869.620 1252.510 869.680 ;
        RECT 1251.270 869.480 1252.510 869.620 ;
        RECT 1251.270 869.420 1251.590 869.480 ;
        RECT 1252.190 869.420 1252.510 869.480 ;
        RECT 1251.730 786.660 1252.050 786.720 ;
        RECT 1251.360 786.520 1252.050 786.660 ;
        RECT 1251.360 786.380 1251.500 786.520 ;
        RECT 1251.730 786.460 1252.050 786.520 ;
        RECT 1251.270 786.120 1251.590 786.380 ;
        RECT 1251.270 738.180 1251.590 738.440 ;
        RECT 1251.360 738.040 1251.500 738.180 ;
        RECT 1251.730 738.040 1252.050 738.100 ;
        RECT 1251.360 737.900 1252.050 738.040 ;
        RECT 1251.730 737.840 1252.050 737.900 ;
        RECT 1251.270 676.160 1251.590 676.220 ;
        RECT 1252.190 676.160 1252.510 676.220 ;
        RECT 1251.270 676.020 1252.510 676.160 ;
        RECT 1251.270 675.960 1251.590 676.020 ;
        RECT 1252.190 675.960 1252.510 676.020 ;
        RECT 1251.730 590.140 1252.050 590.200 ;
        RECT 1251.535 590.000 1252.050 590.140 ;
        RECT 1251.730 589.940 1252.050 590.000 ;
        RECT 1251.745 566.000 1252.035 566.045 ;
        RECT 1252.190 566.000 1252.510 566.060 ;
        RECT 1251.745 565.860 1252.510 566.000 ;
        RECT 1251.745 565.815 1252.035 565.860 ;
        RECT 1252.190 565.800 1252.510 565.860 ;
        RECT 1251.270 524.520 1251.590 524.580 ;
        RECT 1252.190 524.520 1252.510 524.580 ;
        RECT 1251.270 524.380 1252.510 524.520 ;
        RECT 1251.270 524.320 1251.590 524.380 ;
        RECT 1252.190 524.320 1252.510 524.380 ;
        RECT 1250.810 469.440 1251.130 469.500 ;
        RECT 1251.730 469.440 1252.050 469.500 ;
        RECT 1250.810 469.300 1252.050 469.440 ;
        RECT 1250.810 469.240 1251.130 469.300 ;
        RECT 1251.730 469.240 1252.050 469.300 ;
        RECT 1251.270 379.340 1251.590 379.400 ;
        RECT 1251.075 379.200 1251.590 379.340 ;
        RECT 1251.270 379.140 1251.590 379.200 ;
        RECT 1251.270 331.400 1251.590 331.460 ;
        RECT 1251.075 331.260 1251.590 331.400 ;
        RECT 1251.270 331.200 1251.590 331.260 ;
        RECT 1251.730 159.020 1252.050 159.080 ;
        RECT 1251.360 158.880 1252.050 159.020 ;
        RECT 1251.360 158.740 1251.500 158.880 ;
        RECT 1251.730 158.820 1252.050 158.880 ;
        RECT 1251.270 158.480 1251.590 158.740 ;
        RECT 1251.270 96.460 1251.590 96.520 ;
        RECT 1251.075 96.320 1251.590 96.460 ;
        RECT 1251.270 96.260 1251.590 96.320 ;
        RECT 392.910 59.740 393.230 59.800 ;
        RECT 1251.285 59.740 1251.575 59.785 ;
        RECT 392.910 59.600 1251.575 59.740 ;
        RECT 392.910 59.540 393.230 59.600 ;
        RECT 1251.285 59.555 1251.575 59.600 ;
=======
      LAYER met1 ;
        RECT 1249.890 1678.140 1250.210 1678.200 ;
        RECT 1254.030 1678.140 1254.350 1678.200 ;
        RECT 1249.890 1678.000 1254.350 1678.140 ;
        RECT 1249.890 1677.940 1250.210 1678.000 ;
        RECT 1254.030 1677.940 1254.350 1678.000 ;
        RECT 392.910 1528.200 393.230 1528.260 ;
        RECT 1249.890 1528.200 1250.210 1528.260 ;
        RECT 392.910 1528.060 1250.210 1528.200 ;
        RECT 392.910 1528.000 393.230 1528.060 ;
        RECT 1249.890 1528.000 1250.210 1528.060 ;
>>>>>>> re-updated local openlane
        RECT 389.230 16.900 389.550 16.960 ;
        RECT 392.910 16.900 393.230 16.960 ;
        RECT 389.230 16.760 393.230 16.900 ;
        RECT 389.230 16.700 389.550 16.760 ;
        RECT 392.910 16.700 393.230 16.760 ;
      LAYER via ;
        RECT 1249.920 1677.940 1250.180 1678.200 ;
        RECT 1254.060 1677.940 1254.320 1678.200 ;
        RECT 392.940 1528.000 393.200 1528.260 ;
        RECT 1249.920 1528.000 1250.180 1528.260 ;
        RECT 389.260 16.700 389.520 16.960 ;
        RECT 392.940 16.700 393.200 16.960 ;
      LAYER met2 ;
        RECT 1254.970 1700.410 1255.250 1704.000 ;
        RECT 1254.120 1700.270 1255.250 1700.410 ;
        RECT 1254.120 1678.230 1254.260 1700.270 ;
        RECT 1254.970 1700.000 1255.250 1700.270 ;
        RECT 1249.920 1677.910 1250.180 1678.230 ;
        RECT 1254.060 1677.910 1254.320 1678.230 ;
        RECT 1249.980 1528.290 1250.120 1677.910 ;
        RECT 392.940 1527.970 393.200 1528.290 ;
        RECT 1249.920 1527.970 1250.180 1528.290 ;
        RECT 393.000 16.990 393.140 1527.970 ;
        RECT 389.260 16.670 389.520 16.990 ;
        RECT 392.940 16.670 393.200 16.990 ;
        RECT 389.320 2.400 389.460 16.670 ;
        RECT 389.110 -4.800 389.670 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1251.750 1048.760 1252.030 1049.040 ;
        RECT 1253.130 1048.760 1253.410 1049.040 ;
        RECT 1251.290 869.240 1251.570 869.520 ;
        RECT 1252.210 869.240 1252.490 869.520 ;
        RECT 1251.750 676.800 1252.030 677.080 ;
        RECT 1251.290 676.120 1251.570 676.400 ;
      LAYER met3 ;
        RECT 1251.725 1049.050 1252.055 1049.065 ;
        RECT 1253.105 1049.050 1253.435 1049.065 ;
        RECT 1251.725 1048.750 1253.435 1049.050 ;
        RECT 1251.725 1048.735 1252.055 1048.750 ;
        RECT 1253.105 1048.735 1253.435 1048.750 ;
        RECT 1251.265 869.530 1251.595 869.545 ;
        RECT 1252.185 869.530 1252.515 869.545 ;
        RECT 1251.265 869.230 1252.515 869.530 ;
        RECT 1251.265 869.215 1251.595 869.230 ;
        RECT 1252.185 869.215 1252.515 869.230 ;
        RECT 1251.725 677.090 1252.055 677.105 ;
        RECT 1251.510 676.775 1252.055 677.090 ;
        RECT 1251.510 676.425 1251.810 676.775 ;
        RECT 1251.265 676.110 1251.810 676.425 ;
        RECT 1251.265 676.095 1251.595 676.110 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1258.630 1695.480 1258.950 1695.540 ;
        RECT 1260.010 1695.480 1260.330 1695.540 ;
        RECT 1258.630 1695.340 1260.330 1695.480 ;
        RECT 1258.630 1695.280 1258.950 1695.340 ;
        RECT 1260.010 1695.280 1260.330 1695.340 ;
        RECT 1256.790 1678.140 1257.110 1678.200 ;
        RECT 1258.630 1678.140 1258.950 1678.200 ;
        RECT 1256.790 1678.000 1258.950 1678.140 ;
        RECT 1256.790 1677.940 1257.110 1678.000 ;
        RECT 1258.630 1677.940 1258.950 1678.000 ;
        RECT 413.610 1638.700 413.930 1638.760 ;
        RECT 1256.790 1638.700 1257.110 1638.760 ;
        RECT 413.610 1638.560 1257.110 1638.700 ;
        RECT 413.610 1638.500 413.930 1638.560 ;
        RECT 1256.790 1638.500 1257.110 1638.560 ;
        RECT 407.170 16.900 407.490 16.960 ;
        RECT 413.610 16.900 413.930 16.960 ;
        RECT 407.170 16.760 413.930 16.900 ;
        RECT 407.170 16.700 407.490 16.760 ;
        RECT 413.610 16.700 413.930 16.760 ;
      LAYER via ;
        RECT 1258.660 1695.280 1258.920 1695.540 ;
        RECT 1260.040 1695.280 1260.300 1695.540 ;
        RECT 1256.820 1677.940 1257.080 1678.200 ;
        RECT 1258.660 1677.940 1258.920 1678.200 ;
        RECT 413.640 1638.500 413.900 1638.760 ;
        RECT 1256.820 1638.500 1257.080 1638.760 ;
        RECT 407.200 16.700 407.460 16.960 ;
        RECT 413.640 16.700 413.900 16.960 ;
      LAYER met2 ;
        RECT 1260.030 1700.000 1260.310 1704.000 ;
        RECT 1260.100 1695.570 1260.240 1700.000 ;
        RECT 1258.660 1695.250 1258.920 1695.570 ;
        RECT 1260.040 1695.250 1260.300 1695.570 ;
        RECT 1258.720 1678.230 1258.860 1695.250 ;
        RECT 1256.820 1677.910 1257.080 1678.230 ;
        RECT 1258.660 1677.910 1258.920 1678.230 ;
        RECT 1256.880 1638.790 1257.020 1677.910 ;
        RECT 413.640 1638.470 413.900 1638.790 ;
        RECT 1256.820 1638.470 1257.080 1638.790 ;
        RECT 413.700 16.990 413.840 1638.470 ;
        RECT 407.200 16.670 407.460 16.990 ;
        RECT 413.640 16.670 413.900 16.990 ;
        RECT 407.260 2.400 407.400 16.670 ;
        RECT 407.050 -4.800 407.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 0.300 ;
=======
      LAYER met1 ;
        RECT 86.090 1555.740 86.410 1555.800 ;
        RECT 1167.550 1555.740 1167.870 1555.800 ;
        RECT 86.090 1555.600 1167.870 1555.740 ;
        RECT 86.090 1555.540 86.410 1555.600 ;
        RECT 1167.550 1555.540 1167.870 1555.600 ;
        RECT 68.150 19.620 68.470 19.680 ;
        RECT 86.090 19.620 86.410 19.680 ;
        RECT 68.150 19.480 86.410 19.620 ;
        RECT 68.150 19.420 68.470 19.480 ;
        RECT 86.090 19.420 86.410 19.480 ;
      LAYER via ;
        RECT 86.120 1555.540 86.380 1555.800 ;
        RECT 1167.580 1555.540 1167.840 1555.800 ;
        RECT 68.180 19.420 68.440 19.680 ;
        RECT 86.120 19.420 86.380 19.680 ;
      LAYER met2 ;
        RECT 1168.030 1700.410 1168.310 1704.000 ;
        RECT 1167.640 1700.270 1168.310 1700.410 ;
        RECT 1167.640 1555.830 1167.780 1700.270 ;
        RECT 1168.030 1700.000 1168.310 1700.270 ;
        RECT 86.120 1555.510 86.380 1555.830 ;
        RECT 1167.580 1555.510 1167.840 1555.830 ;
        RECT 86.180 19.710 86.320 1555.510 ;
        RECT 68.180 19.390 68.440 19.710 ;
        RECT 86.120 19.390 86.380 19.710 ;
        RECT 68.240 2.400 68.380 19.390 ;
        RECT 68.030 -4.800 68.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 0.300 ;
=======
      LAYER met1 ;
        RECT 1257.250 1683.920 1257.570 1683.980 ;
        RECT 1264.610 1683.920 1264.930 1683.980 ;
        RECT 1257.250 1683.780 1264.930 1683.920 ;
        RECT 1257.250 1683.720 1257.570 1683.780 ;
        RECT 1264.610 1683.720 1264.930 1683.780 ;
        RECT 427.410 1659.440 427.730 1659.500 ;
        RECT 1257.250 1659.440 1257.570 1659.500 ;
        RECT 427.410 1659.300 1257.570 1659.440 ;
        RECT 427.410 1659.240 427.730 1659.300 ;
        RECT 1257.250 1659.240 1257.570 1659.300 ;
        RECT 424.650 16.560 424.970 16.620 ;
        RECT 427.410 16.560 427.730 16.620 ;
        RECT 424.650 16.420 427.730 16.560 ;
        RECT 424.650 16.360 424.970 16.420 ;
        RECT 427.410 16.360 427.730 16.420 ;
      LAYER via ;
        RECT 1257.280 1683.720 1257.540 1683.980 ;
        RECT 1264.640 1683.720 1264.900 1683.980 ;
        RECT 427.440 1659.240 427.700 1659.500 ;
        RECT 1257.280 1659.240 1257.540 1659.500 ;
        RECT 424.680 16.360 424.940 16.620 ;
        RECT 427.440 16.360 427.700 16.620 ;
      LAYER met2 ;
        RECT 1264.630 1700.000 1264.910 1704.000 ;
        RECT 1264.700 1684.010 1264.840 1700.000 ;
        RECT 1257.280 1683.690 1257.540 1684.010 ;
        RECT 1264.640 1683.690 1264.900 1684.010 ;
        RECT 1257.340 1659.530 1257.480 1683.690 ;
        RECT 427.440 1659.210 427.700 1659.530 ;
        RECT 1257.280 1659.210 1257.540 1659.530 ;
        RECT 427.500 16.650 427.640 1659.210 ;
        RECT 424.680 16.330 424.940 16.650 ;
        RECT 427.440 16.330 427.700 16.650 ;
        RECT 424.740 2.400 424.880 16.330 ;
        RECT 424.530 -4.800 425.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 0.300 ;
=======
      LAYER met1 ;
        RECT 448.110 1652.640 448.430 1652.700 ;
        RECT 1269.670 1652.640 1269.990 1652.700 ;
        RECT 448.110 1652.500 1269.990 1652.640 ;
        RECT 448.110 1652.440 448.430 1652.500 ;
        RECT 1269.670 1652.440 1269.990 1652.500 ;
        RECT 442.590 15.880 442.910 15.940 ;
        RECT 448.110 15.880 448.430 15.940 ;
        RECT 442.590 15.740 448.430 15.880 ;
        RECT 442.590 15.680 442.910 15.740 ;
        RECT 448.110 15.680 448.430 15.740 ;
      LAYER via ;
        RECT 448.140 1652.440 448.400 1652.700 ;
        RECT 1269.700 1652.440 1269.960 1652.700 ;
        RECT 442.620 15.680 442.880 15.940 ;
        RECT 448.140 15.680 448.400 15.940 ;
      LAYER met2 ;
        RECT 1269.690 1700.000 1269.970 1704.000 ;
        RECT 1269.760 1652.730 1269.900 1700.000 ;
        RECT 448.140 1652.410 448.400 1652.730 ;
        RECT 1269.700 1652.410 1269.960 1652.730 ;
        RECT 448.200 15.970 448.340 1652.410 ;
        RECT 442.620 15.650 442.880 15.970 ;
        RECT 448.140 15.650 448.400 15.970 ;
        RECT 442.680 2.400 442.820 15.650 ;
        RECT 442.470 -4.800 443.030 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 0.300 ;
=======
      LAYER li1 ;
        RECT 1272.045 1449.165 1272.215 1497.275 ;
        RECT 1271.585 710.685 1271.755 738.395 ;
        RECT 1271.585 469.285 1271.755 502.095 ;
        RECT 1271.585 179.605 1271.755 227.715 ;
        RECT 1272.045 60.945 1272.215 131.155 ;
      LAYER mcon ;
        RECT 1272.045 1497.105 1272.215 1497.275 ;
        RECT 1271.585 738.225 1271.755 738.395 ;
        RECT 1271.585 501.925 1271.755 502.095 ;
        RECT 1271.585 227.545 1271.755 227.715 ;
        RECT 1272.045 130.985 1272.215 131.155 ;
      LAYER met1 ;
        RECT 1271.510 1545.880 1271.830 1545.940 ;
        RECT 1271.970 1545.880 1272.290 1545.940 ;
        RECT 1271.510 1545.740 1272.290 1545.880 ;
        RECT 1271.510 1545.680 1271.830 1545.740 ;
        RECT 1271.970 1545.680 1272.290 1545.740 ;
        RECT 1271.510 1511.340 1271.830 1511.600 ;
        RECT 1271.600 1510.520 1271.740 1511.340 ;
        RECT 1271.970 1510.520 1272.290 1510.580 ;
        RECT 1271.600 1510.380 1272.290 1510.520 ;
        RECT 1271.970 1510.320 1272.290 1510.380 ;
        RECT 1271.970 1497.260 1272.290 1497.320 ;
        RECT 1271.775 1497.120 1272.290 1497.260 ;
        RECT 1271.970 1497.060 1272.290 1497.120 ;
        RECT 1271.970 1449.320 1272.290 1449.380 ;
        RECT 1271.775 1449.180 1272.290 1449.320 ;
        RECT 1271.970 1449.120 1272.290 1449.180 ;
        RECT 1271.510 1269.600 1271.830 1269.860 ;
        RECT 1271.600 1269.120 1271.740 1269.600 ;
        RECT 1271.970 1269.120 1272.290 1269.180 ;
        RECT 1271.600 1268.980 1272.290 1269.120 ;
        RECT 1271.970 1268.920 1272.290 1268.980 ;
        RECT 1271.970 1207.920 1272.290 1207.980 ;
        RECT 1271.600 1207.780 1272.290 1207.920 ;
        RECT 1271.600 1207.640 1271.740 1207.780 ;
        RECT 1271.970 1207.720 1272.290 1207.780 ;
        RECT 1271.510 1207.380 1271.830 1207.640 ;
        RECT 1271.510 1152.500 1271.830 1152.560 ;
        RECT 1271.970 1152.500 1272.290 1152.560 ;
        RECT 1271.510 1152.360 1272.290 1152.500 ;
        RECT 1271.510 1152.300 1271.830 1152.360 ;
        RECT 1271.970 1152.300 1272.290 1152.360 ;
        RECT 1271.510 966.180 1271.830 966.240 ;
        RECT 1271.970 966.180 1272.290 966.240 ;
        RECT 1271.510 966.040 1272.290 966.180 ;
        RECT 1271.510 965.980 1271.830 966.040 ;
        RECT 1271.970 965.980 1272.290 966.040 ;
        RECT 1270.590 959.040 1270.910 959.100 ;
        RECT 1271.970 959.040 1272.290 959.100 ;
        RECT 1270.590 958.900 1272.290 959.040 ;
        RECT 1270.590 958.840 1270.910 958.900 ;
        RECT 1271.970 958.840 1272.290 958.900 ;
        RECT 1271.510 910.760 1271.830 910.820 ;
        RECT 1272.430 910.760 1272.750 910.820 ;
        RECT 1271.510 910.620 1272.750 910.760 ;
        RECT 1271.510 910.560 1271.830 910.620 ;
        RECT 1272.430 910.560 1272.750 910.620 ;
        RECT 1271.510 759.260 1271.830 759.520 ;
        RECT 1271.600 758.840 1271.740 759.260 ;
        RECT 1271.510 758.580 1271.830 758.840 ;
        RECT 1271.510 738.380 1271.830 738.440 ;
        RECT 1271.315 738.240 1271.830 738.380 ;
        RECT 1271.510 738.180 1271.830 738.240 ;
        RECT 1271.525 710.840 1271.815 710.885 ;
        RECT 1272.430 710.840 1272.750 710.900 ;
        RECT 1271.525 710.700 1272.750 710.840 ;
        RECT 1271.525 710.655 1271.815 710.700 ;
        RECT 1272.430 710.640 1272.750 710.700 ;
        RECT 1271.510 572.940 1271.830 573.200 ;
        RECT 1271.600 572.800 1271.740 572.940 ;
        RECT 1271.970 572.800 1272.290 572.860 ;
        RECT 1271.600 572.660 1272.290 572.800 ;
        RECT 1271.970 572.600 1272.290 572.660 ;
        RECT 1271.510 502.080 1271.830 502.140 ;
        RECT 1271.315 501.940 1271.830 502.080 ;
        RECT 1271.510 501.880 1271.830 501.940 ;
        RECT 1271.525 469.440 1271.815 469.485 ;
        RECT 1271.970 469.440 1272.290 469.500 ;
        RECT 1271.525 469.300 1272.290 469.440 ;
        RECT 1271.525 469.255 1271.815 469.300 ;
        RECT 1271.970 469.240 1272.290 469.300 ;
        RECT 1271.510 283.120 1271.830 283.180 ;
        RECT 1272.430 283.120 1272.750 283.180 ;
        RECT 1271.510 282.980 1272.750 283.120 ;
        RECT 1271.510 282.920 1271.830 282.980 ;
        RECT 1272.430 282.920 1272.750 282.980 ;
        RECT 1271.510 227.700 1271.830 227.760 ;
        RECT 1271.315 227.560 1271.830 227.700 ;
        RECT 1271.510 227.500 1271.830 227.560 ;
        RECT 1271.525 179.760 1271.815 179.805 ;
        RECT 1272.430 179.760 1272.750 179.820 ;
        RECT 1271.525 179.620 1272.750 179.760 ;
        RECT 1271.525 179.575 1271.815 179.620 ;
        RECT 1272.430 179.560 1272.750 179.620 ;
        RECT 1271.970 131.140 1272.290 131.200 ;
        RECT 1271.775 131.000 1272.290 131.140 ;
        RECT 1271.970 130.940 1272.290 131.000 ;
        RECT 461.910 61.100 462.230 61.160 ;
        RECT 1271.985 61.100 1272.275 61.145 ;
        RECT 461.910 60.960 1272.275 61.100 ;
        RECT 461.910 60.900 462.230 60.960 ;
        RECT 1271.985 60.915 1272.275 60.960 ;
=======
      LAYER met1 ;
        RECT 461.910 1514.600 462.230 1514.660 ;
        RECT 1272.430 1514.600 1272.750 1514.660 ;
        RECT 461.910 1514.460 1272.750 1514.600 ;
        RECT 461.910 1514.400 462.230 1514.460 ;
        RECT 1272.430 1514.400 1272.750 1514.460 ;
>>>>>>> re-updated local openlane
        RECT 460.530 2.960 460.850 3.020 ;
        RECT 461.910 2.960 462.230 3.020 ;
        RECT 460.530 2.820 462.230 2.960 ;
        RECT 460.530 2.760 460.850 2.820 ;
        RECT 461.910 2.760 462.230 2.820 ;
      LAYER via ;
        RECT 461.940 1514.400 462.200 1514.660 ;
        RECT 1272.460 1514.400 1272.720 1514.660 ;
        RECT 460.560 2.760 460.820 3.020 ;
        RECT 461.940 2.760 462.200 3.020 ;
      LAYER met2 ;
        RECT 1274.290 1700.410 1274.570 1704.000 ;
        RECT 1273.900 1700.270 1274.570 1700.410 ;
        RECT 1273.900 1668.450 1274.040 1700.270 ;
        RECT 1274.290 1700.000 1274.570 1700.270 ;
        RECT 1272.980 1668.310 1274.040 1668.450 ;
        RECT 1272.980 1558.970 1273.120 1668.310 ;
        RECT 1272.520 1558.830 1273.120 1558.970 ;
        RECT 1272.520 1514.690 1272.660 1558.830 ;
        RECT 461.940 1514.370 462.200 1514.690 ;
        RECT 1272.460 1514.370 1272.720 1514.690 ;
        RECT 462.000 3.050 462.140 1514.370 ;
        RECT 460.560 2.730 460.820 3.050 ;
        RECT 461.940 2.730 462.200 3.050 ;
        RECT 460.620 2.400 460.760 2.730 ;
        RECT 460.410 -4.800 460.970 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1271.990 1401.680 1272.270 1401.960 ;
        RECT 1271.530 1401.000 1271.810 1401.280 ;
        RECT 1270.610 910.720 1270.890 911.000 ;
        RECT 1271.530 910.720 1271.810 911.000 ;
        RECT 1271.530 820.960 1271.810 821.240 ;
        RECT 1272.450 820.960 1272.730 821.240 ;
        RECT 1271.990 628.520 1272.270 628.800 ;
        RECT 1271.530 627.840 1271.810 628.120 ;
      LAYER met3 ;
        RECT 1271.965 1401.970 1272.295 1401.985 ;
        RECT 1270.830 1401.670 1272.295 1401.970 ;
        RECT 1270.830 1401.290 1271.130 1401.670 ;
        RECT 1271.965 1401.655 1272.295 1401.670 ;
        RECT 1271.505 1401.290 1271.835 1401.305 ;
        RECT 1270.830 1400.990 1271.835 1401.290 ;
        RECT 1271.505 1400.975 1271.835 1400.990 ;
        RECT 1270.585 911.010 1270.915 911.025 ;
        RECT 1271.505 911.010 1271.835 911.025 ;
        RECT 1270.585 910.710 1271.835 911.010 ;
        RECT 1270.585 910.695 1270.915 910.710 ;
        RECT 1271.505 910.695 1271.835 910.710 ;
        RECT 1271.505 821.250 1271.835 821.265 ;
        RECT 1272.425 821.250 1272.755 821.265 ;
        RECT 1271.505 820.950 1272.755 821.250 ;
        RECT 1271.505 820.935 1271.835 820.950 ;
        RECT 1272.425 820.935 1272.755 820.950 ;
        RECT 1271.965 628.810 1272.295 628.825 ;
        RECT 1271.750 628.495 1272.295 628.810 ;
        RECT 1271.750 628.145 1272.050 628.495 ;
        RECT 1271.505 627.830 1272.050 628.145 ;
        RECT 1271.505 627.815 1271.835 627.830 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 0.300 ;
=======
      LAYER met1 ;
        RECT 482.610 1521.400 482.930 1521.460 ;
        RECT 1277.950 1521.400 1278.270 1521.460 ;
        RECT 482.610 1521.260 1278.270 1521.400 ;
        RECT 482.610 1521.200 482.930 1521.260 ;
        RECT 1277.950 1521.200 1278.270 1521.260 ;
        RECT 478.470 15.540 478.790 15.600 ;
        RECT 482.610 15.540 482.930 15.600 ;
        RECT 478.470 15.400 482.930 15.540 ;
        RECT 478.470 15.340 478.790 15.400 ;
        RECT 482.610 15.340 482.930 15.400 ;
      LAYER via ;
        RECT 482.640 1521.200 482.900 1521.460 ;
        RECT 1277.980 1521.200 1278.240 1521.460 ;
        RECT 478.500 15.340 478.760 15.600 ;
        RECT 482.640 15.340 482.900 15.600 ;
      LAYER met2 ;
        RECT 1279.350 1700.410 1279.630 1704.000 ;
        RECT 1278.040 1700.270 1279.630 1700.410 ;
        RECT 1278.040 1521.490 1278.180 1700.270 ;
        RECT 1279.350 1700.000 1279.630 1700.270 ;
        RECT 482.640 1521.170 482.900 1521.490 ;
        RECT 1277.980 1521.170 1278.240 1521.490 ;
        RECT 482.700 15.630 482.840 1521.170 ;
        RECT 478.500 15.310 478.760 15.630 ;
        RECT 482.640 15.310 482.900 15.630 ;
        RECT 478.560 2.400 478.700 15.310 ;
        RECT 478.350 -4.800 478.910 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 0.300 ;
=======
      LAYER met1 ;
        RECT 496.410 61.780 496.730 61.840 ;
        RECT 1284.850 61.780 1285.170 61.840 ;
        RECT 496.410 61.640 1285.170 61.780 ;
        RECT 496.410 61.580 496.730 61.640 ;
        RECT 1284.850 61.580 1285.170 61.640 ;
      LAYER via ;
        RECT 496.440 61.580 496.700 61.840 ;
        RECT 1284.880 61.580 1285.140 61.840 ;
      LAYER met2 ;
        RECT 1283.490 1700.410 1283.770 1704.000 ;
        RECT 1283.490 1700.270 1285.080 1700.410 ;
        RECT 1283.490 1700.000 1283.770 1700.270 ;
        RECT 1284.940 61.870 1285.080 1700.270 ;
        RECT 496.440 61.550 496.700 61.870 ;
        RECT 1284.880 61.550 1285.140 61.870 ;
        RECT 496.500 2.400 496.640 61.550 ;
=======
      LAYER li1 ;
        RECT 1252.265 1635.485 1252.435 1683.595 ;
        RECT 1252.265 1538.925 1252.435 1587.035 ;
      LAYER mcon ;
        RECT 1252.265 1683.425 1252.435 1683.595 ;
        RECT 1252.265 1586.865 1252.435 1587.035 ;
      LAYER met1 ;
        RECT 1252.650 1688.000 1252.970 1688.060 ;
        RECT 1284.390 1688.000 1284.710 1688.060 ;
        RECT 1252.650 1687.860 1284.710 1688.000 ;
        RECT 1252.650 1687.800 1252.970 1687.860 ;
        RECT 1284.390 1687.800 1284.710 1687.860 ;
        RECT 1252.205 1683.580 1252.495 1683.625 ;
        RECT 1252.650 1683.580 1252.970 1683.640 ;
        RECT 1252.205 1683.440 1252.970 1683.580 ;
        RECT 1252.205 1683.395 1252.495 1683.440 ;
        RECT 1252.650 1683.380 1252.970 1683.440 ;
        RECT 1252.190 1635.640 1252.510 1635.700 ;
        RECT 1251.995 1635.500 1252.510 1635.640 ;
        RECT 1252.190 1635.440 1252.510 1635.500 ;
        RECT 1252.190 1587.020 1252.510 1587.080 ;
        RECT 1251.995 1586.880 1252.510 1587.020 ;
        RECT 1252.190 1586.820 1252.510 1586.880 ;
        RECT 1252.190 1539.080 1252.510 1539.140 ;
        RECT 1251.995 1538.940 1252.510 1539.080 ;
        RECT 1252.190 1538.880 1252.510 1538.940 ;
        RECT 1251.730 1111.020 1252.050 1111.080 ;
        RECT 1252.190 1111.020 1252.510 1111.080 ;
        RECT 1251.730 1110.880 1252.510 1111.020 ;
        RECT 1251.730 1110.820 1252.050 1110.880 ;
        RECT 1252.190 1110.820 1252.510 1110.880 ;
        RECT 1251.730 1062.740 1252.050 1062.800 ;
        RECT 1252.190 1062.740 1252.510 1062.800 ;
        RECT 1251.730 1062.600 1252.510 1062.740 ;
        RECT 1251.730 1062.540 1252.050 1062.600 ;
        RECT 1252.190 1062.540 1252.510 1062.600 ;
        RECT 496.410 72.320 496.730 72.380 ;
        RECT 1252.190 72.320 1252.510 72.380 ;
        RECT 496.410 72.180 1252.510 72.320 ;
        RECT 496.410 72.120 496.730 72.180 ;
        RECT 1252.190 72.120 1252.510 72.180 ;
      LAYER via ;
        RECT 1252.680 1687.800 1252.940 1688.060 ;
        RECT 1284.420 1687.800 1284.680 1688.060 ;
        RECT 1252.680 1683.380 1252.940 1683.640 ;
        RECT 1252.220 1635.440 1252.480 1635.700 ;
        RECT 1252.220 1586.820 1252.480 1587.080 ;
        RECT 1252.220 1538.880 1252.480 1539.140 ;
        RECT 1251.760 1110.820 1252.020 1111.080 ;
        RECT 1252.220 1110.820 1252.480 1111.080 ;
        RECT 1251.760 1062.540 1252.020 1062.800 ;
        RECT 1252.220 1062.540 1252.480 1062.800 ;
        RECT 496.440 72.120 496.700 72.380 ;
        RECT 1252.220 72.120 1252.480 72.380 ;
      LAYER met2 ;
        RECT 1284.410 1700.000 1284.690 1704.000 ;
        RECT 1284.480 1688.090 1284.620 1700.000 ;
        RECT 1252.680 1687.770 1252.940 1688.090 ;
        RECT 1284.420 1687.770 1284.680 1688.090 ;
        RECT 1252.740 1683.670 1252.880 1687.770 ;
        RECT 1252.680 1683.350 1252.940 1683.670 ;
        RECT 1252.220 1635.410 1252.480 1635.730 ;
        RECT 1252.280 1587.110 1252.420 1635.410 ;
        RECT 1252.220 1586.790 1252.480 1587.110 ;
        RECT 1252.220 1538.850 1252.480 1539.170 ;
        RECT 1252.280 1111.110 1252.420 1538.850 ;
        RECT 1251.760 1110.790 1252.020 1111.110 ;
        RECT 1252.220 1110.790 1252.480 1111.110 ;
        RECT 1251.820 1062.830 1251.960 1110.790 ;
        RECT 1251.760 1062.510 1252.020 1062.830 ;
        RECT 1252.220 1062.510 1252.480 1062.830 ;
        RECT 1252.280 72.410 1252.420 1062.510 ;
        RECT 496.440 72.090 496.700 72.410 ;
        RECT 1252.220 72.090 1252.480 72.410 ;
        RECT 496.500 2.400 496.640 72.090 ;
>>>>>>> re-updated local openlane
        RECT 496.290 -4.800 496.850 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 0.300 ;
=======
      LAYER met1 ;
        RECT 1283.930 1678.140 1284.250 1678.200 ;
        RECT 1288.070 1678.140 1288.390 1678.200 ;
        RECT 1283.930 1678.000 1288.390 1678.140 ;
        RECT 1283.930 1677.940 1284.250 1678.000 ;
        RECT 1288.070 1677.940 1288.390 1678.000 ;
        RECT 517.110 1493.860 517.430 1493.920 ;
        RECT 1283.930 1493.860 1284.250 1493.920 ;
        RECT 517.110 1493.720 1284.250 1493.860 ;
        RECT 517.110 1493.660 517.430 1493.720 ;
        RECT 1283.930 1493.660 1284.250 1493.720 ;
        RECT 513.890 15.540 514.210 15.600 ;
        RECT 517.110 15.540 517.430 15.600 ;
        RECT 513.890 15.400 517.430 15.540 ;
        RECT 513.890 15.340 514.210 15.400 ;
        RECT 517.110 15.340 517.430 15.400 ;
      LAYER via ;
        RECT 1283.960 1677.940 1284.220 1678.200 ;
        RECT 1288.100 1677.940 1288.360 1678.200 ;
        RECT 517.140 1493.660 517.400 1493.920 ;
        RECT 1283.960 1493.660 1284.220 1493.920 ;
        RECT 513.920 15.340 514.180 15.600 ;
        RECT 517.140 15.340 517.400 15.600 ;
      LAYER met2 ;
        RECT 1289.010 1700.410 1289.290 1704.000 ;
        RECT 1288.160 1700.270 1289.290 1700.410 ;
        RECT 1288.160 1678.230 1288.300 1700.270 ;
        RECT 1289.010 1700.000 1289.290 1700.270 ;
        RECT 1283.960 1677.910 1284.220 1678.230 ;
        RECT 1288.100 1677.910 1288.360 1678.230 ;
        RECT 1284.020 1493.950 1284.160 1677.910 ;
        RECT 517.140 1493.630 517.400 1493.950 ;
        RECT 1283.960 1493.630 1284.220 1493.950 ;
        RECT 517.200 15.630 517.340 1493.630 ;
        RECT 513.920 15.310 514.180 15.630 ;
        RECT 517.140 15.310 517.400 15.630 ;
        RECT 513.980 2.400 514.120 15.310 ;
        RECT 513.770 -4.800 514.330 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 0.300 ;
=======
      LAYER met1 ;
        RECT 1291.290 1677.120 1291.610 1677.180 ;
        RECT 1292.670 1677.120 1292.990 1677.180 ;
        RECT 1291.290 1676.980 1292.990 1677.120 ;
        RECT 1291.290 1676.920 1291.610 1676.980 ;
        RECT 1292.670 1676.920 1292.990 1676.980 ;
        RECT 537.350 1507.460 537.670 1507.520 ;
        RECT 1291.290 1507.460 1291.610 1507.520 ;
        RECT 537.350 1507.320 1291.610 1507.460 ;
        RECT 537.350 1507.260 537.670 1507.320 ;
        RECT 1291.290 1507.260 1291.610 1507.320 ;
        RECT 531.830 15.540 532.150 15.600 ;
        RECT 537.350 15.540 537.670 15.600 ;
        RECT 531.830 15.400 537.670 15.540 ;
        RECT 531.830 15.340 532.150 15.400 ;
        RECT 537.350 15.340 537.670 15.400 ;
      LAYER via ;
        RECT 1291.320 1676.920 1291.580 1677.180 ;
        RECT 1292.700 1676.920 1292.960 1677.180 ;
        RECT 537.380 1507.260 537.640 1507.520 ;
        RECT 1291.320 1507.260 1291.580 1507.520 ;
        RECT 531.860 15.340 532.120 15.600 ;
        RECT 537.380 15.340 537.640 15.600 ;
      LAYER met2 ;
        RECT 1294.070 1700.410 1294.350 1704.000 ;
        RECT 1292.760 1700.270 1294.350 1700.410 ;
        RECT 1292.760 1677.210 1292.900 1700.270 ;
        RECT 1294.070 1700.000 1294.350 1700.270 ;
        RECT 1291.320 1676.890 1291.580 1677.210 ;
        RECT 1292.700 1676.890 1292.960 1677.210 ;
        RECT 1291.380 1507.550 1291.520 1676.890 ;
        RECT 537.380 1507.230 537.640 1507.550 ;
        RECT 1291.320 1507.230 1291.580 1507.550 ;
        RECT 537.440 15.630 537.580 1507.230 ;
        RECT 531.860 15.310 532.120 15.630 ;
        RECT 537.380 15.310 537.640 15.630 ;
        RECT 531.920 2.400 532.060 15.310 ;
        RECT 531.710 -4.800 532.270 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 0.300 ;
=======
      LAYER met1 ;
        RECT 1286.690 1684.260 1287.010 1684.320 ;
        RECT 1298.650 1684.260 1298.970 1684.320 ;
        RECT 1286.690 1684.120 1298.970 1684.260 ;
        RECT 1286.690 1684.060 1287.010 1684.120 ;
        RECT 1298.650 1684.060 1298.970 1684.120 ;
        RECT 551.610 1052.200 551.930 1052.260 ;
        RECT 1286.690 1052.200 1287.010 1052.260 ;
        RECT 551.610 1052.060 1287.010 1052.200 ;
        RECT 551.610 1052.000 551.930 1052.060 ;
        RECT 1286.690 1052.000 1287.010 1052.060 ;
      LAYER via ;
        RECT 1286.720 1684.060 1286.980 1684.320 ;
        RECT 1298.680 1684.060 1298.940 1684.320 ;
        RECT 551.640 1052.000 551.900 1052.260 ;
        RECT 1286.720 1052.000 1286.980 1052.260 ;
      LAYER met2 ;
        RECT 1298.670 1700.000 1298.950 1704.000 ;
        RECT 1298.740 1684.350 1298.880 1700.000 ;
        RECT 1286.720 1684.030 1286.980 1684.350 ;
        RECT 1298.680 1684.030 1298.940 1684.350 ;
        RECT 1286.780 1052.290 1286.920 1684.030 ;
        RECT 551.640 1051.970 551.900 1052.290 ;
        RECT 1286.720 1051.970 1286.980 1052.290 ;
        RECT 551.700 17.410 551.840 1051.970 ;
        RECT 549.860 17.270 551.840 17.410 ;
        RECT 549.860 2.400 550.000 17.270 ;
        RECT 549.650 -4.800 550.210 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 0.300 ;
=======
      LAYER li1 ;
        RECT 1298.265 1338.665 1298.435 1345.975 ;
        RECT 1298.265 655.605 1298.435 703.375 ;
        RECT 1298.265 559.045 1298.435 607.155 ;
        RECT 1298.265 493.425 1298.435 517.395 ;
        RECT 1298.265 372.725 1298.435 380.035 ;
        RECT 1298.265 324.445 1298.435 331.415 ;
        RECT 600.905 15.045 601.075 17.935 ;
      LAYER mcon ;
        RECT 1298.265 1345.805 1298.435 1345.975 ;
        RECT 1298.265 703.205 1298.435 703.375 ;
        RECT 1298.265 606.985 1298.435 607.155 ;
        RECT 1298.265 517.225 1298.435 517.395 ;
        RECT 1298.265 379.865 1298.435 380.035 ;
        RECT 1298.265 331.245 1298.435 331.415 ;
        RECT 600.905 17.765 601.075 17.935 ;
      LAYER met1 ;
        RECT 1298.650 1387.100 1298.970 1387.160 ;
        RECT 1299.570 1387.100 1299.890 1387.160 ;
        RECT 1298.650 1386.960 1299.890 1387.100 ;
        RECT 1298.650 1386.900 1298.970 1386.960 ;
        RECT 1299.570 1386.900 1299.890 1386.960 ;
        RECT 1298.205 1345.960 1298.495 1346.005 ;
        RECT 1298.650 1345.960 1298.970 1346.020 ;
        RECT 1298.205 1345.820 1298.970 1345.960 ;
        RECT 1298.205 1345.775 1298.495 1345.820 ;
        RECT 1298.650 1345.760 1298.970 1345.820 ;
        RECT 1298.190 1338.820 1298.510 1338.880 ;
        RECT 1297.995 1338.680 1298.510 1338.820 ;
        RECT 1298.190 1338.620 1298.510 1338.680 ;
        RECT 1298.190 1152.500 1298.510 1152.560 ;
        RECT 1298.650 1152.500 1298.970 1152.560 ;
        RECT 1298.190 1152.360 1298.970 1152.500 ;
        RECT 1298.190 1152.300 1298.510 1152.360 ;
        RECT 1298.650 1152.300 1298.970 1152.360 ;
        RECT 1298.650 1125.300 1298.970 1125.360 ;
        RECT 1298.280 1125.160 1298.970 1125.300 ;
        RECT 1298.280 1124.680 1298.420 1125.160 ;
        RECT 1298.650 1125.100 1298.970 1125.160 ;
        RECT 1298.190 1124.420 1298.510 1124.680 ;
        RECT 1298.190 959.380 1298.510 959.440 ;
        RECT 1298.650 959.380 1298.970 959.440 ;
        RECT 1298.190 959.240 1298.970 959.380 ;
        RECT 1298.190 959.180 1298.510 959.240 ;
        RECT 1298.650 959.180 1298.970 959.240 ;
        RECT 1297.270 958.700 1297.590 958.760 ;
        RECT 1298.190 958.700 1298.510 958.760 ;
        RECT 1297.270 958.560 1298.510 958.700 ;
        RECT 1297.270 958.500 1297.590 958.560 ;
        RECT 1298.190 958.500 1298.510 958.560 ;
        RECT 1298.650 710.500 1298.970 710.560 ;
        RECT 1299.110 710.500 1299.430 710.560 ;
        RECT 1298.650 710.360 1299.430 710.500 ;
        RECT 1298.650 710.300 1298.970 710.360 ;
        RECT 1299.110 710.300 1299.430 710.360 ;
        RECT 1298.650 703.500 1298.970 703.760 ;
        RECT 1298.205 703.360 1298.495 703.405 ;
        RECT 1298.740 703.360 1298.880 703.500 ;
        RECT 1298.205 703.220 1298.880 703.360 ;
        RECT 1298.205 703.175 1298.495 703.220 ;
        RECT 1298.190 655.760 1298.510 655.820 ;
        RECT 1297.995 655.620 1298.510 655.760 ;
        RECT 1298.190 655.560 1298.510 655.620 ;
        RECT 1297.270 638.420 1297.590 638.480 ;
        RECT 1298.190 638.420 1298.510 638.480 ;
        RECT 1297.270 638.280 1298.510 638.420 ;
        RECT 1297.270 638.220 1297.590 638.280 ;
        RECT 1298.190 638.220 1298.510 638.280 ;
        RECT 1298.190 607.140 1298.510 607.200 ;
        RECT 1297.995 607.000 1298.510 607.140 ;
        RECT 1298.190 606.940 1298.510 607.000 ;
        RECT 1298.205 559.200 1298.495 559.245 ;
        RECT 1299.110 559.200 1299.430 559.260 ;
        RECT 1298.205 559.060 1299.430 559.200 ;
        RECT 1298.205 559.015 1298.495 559.060 ;
        RECT 1299.110 559.000 1299.430 559.060 ;
        RECT 1298.190 542.540 1298.510 542.600 ;
        RECT 1299.110 542.540 1299.430 542.600 ;
        RECT 1298.190 542.400 1299.430 542.540 ;
        RECT 1298.190 542.340 1298.510 542.400 ;
        RECT 1299.110 542.340 1299.430 542.400 ;
        RECT 1298.190 517.380 1298.510 517.440 ;
        RECT 1297.995 517.240 1298.510 517.380 ;
        RECT 1298.190 517.180 1298.510 517.240 ;
        RECT 1298.190 493.580 1298.510 493.640 ;
        RECT 1297.995 493.440 1298.510 493.580 ;
        RECT 1298.190 493.380 1298.510 493.440 ;
        RECT 1298.190 434.760 1298.510 434.820 ;
        RECT 1298.650 434.760 1298.970 434.820 ;
        RECT 1298.190 434.620 1298.970 434.760 ;
        RECT 1298.190 434.560 1298.510 434.620 ;
        RECT 1298.650 434.560 1298.970 434.620 ;
        RECT 1298.205 380.020 1298.495 380.065 ;
        RECT 1298.650 380.020 1298.970 380.080 ;
        RECT 1298.205 379.880 1298.970 380.020 ;
        RECT 1298.205 379.835 1298.495 379.880 ;
        RECT 1298.650 379.820 1298.970 379.880 ;
        RECT 1298.190 372.880 1298.510 372.940 ;
        RECT 1297.995 372.740 1298.510 372.880 ;
        RECT 1298.190 372.680 1298.510 372.740 ;
        RECT 1298.190 331.400 1298.510 331.460 ;
        RECT 1297.995 331.260 1298.510 331.400 ;
        RECT 1298.190 331.200 1298.510 331.260 ;
        RECT 1298.190 324.600 1298.510 324.660 ;
        RECT 1297.995 324.460 1298.510 324.600 ;
        RECT 1298.190 324.400 1298.510 324.460 ;
        RECT 1298.650 145.080 1298.970 145.140 ;
        RECT 1299.110 145.080 1299.430 145.140 ;
        RECT 1298.650 144.940 1299.430 145.080 ;
        RECT 1298.650 144.880 1298.970 144.940 ;
        RECT 1299.110 144.880 1299.430 144.940 ;
        RECT 567.710 17.920 568.030 17.980 ;
        RECT 600.845 17.920 601.135 17.965 ;
        RECT 567.710 17.780 601.135 17.920 ;
        RECT 567.710 17.720 568.030 17.780 ;
        RECT 600.845 17.735 601.135 17.780 ;
        RECT 600.845 15.200 601.135 15.245 ;
        RECT 1298.190 15.200 1298.510 15.260 ;
        RECT 600.845 15.060 1298.510 15.200 ;
        RECT 600.845 15.015 601.135 15.060 ;
        RECT 1298.190 15.000 1298.510 15.060 ;
      LAYER via ;
        RECT 1298.680 1386.900 1298.940 1387.160 ;
        RECT 1299.600 1386.900 1299.860 1387.160 ;
        RECT 1298.680 1345.760 1298.940 1346.020 ;
        RECT 1298.220 1338.620 1298.480 1338.880 ;
        RECT 1298.220 1152.300 1298.480 1152.560 ;
        RECT 1298.680 1152.300 1298.940 1152.560 ;
        RECT 1298.680 1125.100 1298.940 1125.360 ;
        RECT 1298.220 1124.420 1298.480 1124.680 ;
        RECT 1298.220 959.180 1298.480 959.440 ;
        RECT 1298.680 959.180 1298.940 959.440 ;
        RECT 1297.300 958.500 1297.560 958.760 ;
        RECT 1298.220 958.500 1298.480 958.760 ;
        RECT 1298.680 710.300 1298.940 710.560 ;
        RECT 1299.140 710.300 1299.400 710.560 ;
        RECT 1298.680 703.500 1298.940 703.760 ;
        RECT 1298.220 655.560 1298.480 655.820 ;
        RECT 1297.300 638.220 1297.560 638.480 ;
        RECT 1298.220 638.220 1298.480 638.480 ;
        RECT 1298.220 606.940 1298.480 607.200 ;
        RECT 1299.140 559.000 1299.400 559.260 ;
        RECT 1298.220 542.340 1298.480 542.600 ;
        RECT 1299.140 542.340 1299.400 542.600 ;
        RECT 1298.220 517.180 1298.480 517.440 ;
        RECT 1298.220 493.380 1298.480 493.640 ;
        RECT 1298.220 434.560 1298.480 434.820 ;
        RECT 1298.680 434.560 1298.940 434.820 ;
        RECT 1298.680 379.820 1298.940 380.080 ;
        RECT 1298.220 372.680 1298.480 372.940 ;
        RECT 1298.220 331.200 1298.480 331.460 ;
        RECT 1298.220 324.400 1298.480 324.660 ;
        RECT 1298.680 144.880 1298.940 145.140 ;
        RECT 1299.140 144.880 1299.400 145.140 ;
        RECT 567.740 17.720 568.000 17.980 ;
        RECT 1298.220 15.000 1298.480 15.260 ;
      LAYER met2 ;
        RECT 1302.810 1700.410 1303.090 1704.000 ;
        RECT 1302.420 1700.270 1303.090 1700.410 ;
        RECT 1302.420 1656.210 1302.560 1700.270 ;
        RECT 1302.810 1700.000 1303.090 1700.270 ;
        RECT 1298.740 1656.070 1302.560 1656.210 ;
        RECT 1298.740 1435.325 1298.880 1656.070 ;
        RECT 1298.670 1434.955 1298.950 1435.325 ;
        RECT 1299.590 1434.955 1299.870 1435.325 ;
        RECT 1299.660 1387.190 1299.800 1434.955 ;
        RECT 1298.680 1386.870 1298.940 1387.190 ;
        RECT 1299.600 1386.870 1299.860 1387.190 ;
        RECT 1298.740 1346.050 1298.880 1386.870 ;
        RECT 1298.680 1345.730 1298.940 1346.050 ;
        RECT 1298.220 1338.590 1298.480 1338.910 ;
        RECT 1298.280 1152.590 1298.420 1338.590 ;
        RECT 1298.220 1152.270 1298.480 1152.590 ;
        RECT 1298.680 1152.270 1298.940 1152.590 ;
        RECT 1298.740 1125.390 1298.880 1152.270 ;
        RECT 1298.680 1125.070 1298.940 1125.390 ;
        RECT 1298.220 1124.390 1298.480 1124.710 ;
        RECT 1298.280 1007.490 1298.420 1124.390 ;
        RECT 1298.280 1007.350 1298.880 1007.490 ;
        RECT 1298.740 959.470 1298.880 1007.350 ;
        RECT 1298.220 959.150 1298.480 959.470 ;
        RECT 1298.680 959.150 1298.940 959.470 ;
        RECT 1298.280 958.790 1298.420 959.150 ;
        RECT 1297.300 958.470 1297.560 958.790 ;
        RECT 1298.220 958.470 1298.480 958.790 ;
        RECT 1297.360 911.045 1297.500 958.470 ;
        RECT 1297.290 910.675 1297.570 911.045 ;
        RECT 1298.670 910.675 1298.950 911.045 ;
        RECT 1298.740 886.450 1298.880 910.675 ;
        RECT 1298.740 886.310 1299.340 886.450 ;
        RECT 1299.200 821.285 1299.340 886.310 ;
        RECT 1298.210 820.915 1298.490 821.285 ;
        RECT 1299.130 820.915 1299.410 821.285 ;
        RECT 1298.280 766.090 1298.420 820.915 ;
        RECT 1298.280 765.950 1298.880 766.090 ;
        RECT 1298.740 741.610 1298.880 765.950 ;
        RECT 1298.740 741.470 1299.340 741.610 ;
        RECT 1299.200 710.590 1299.340 741.470 ;
        RECT 1298.680 710.270 1298.940 710.590 ;
        RECT 1299.140 710.270 1299.400 710.590 ;
        RECT 1298.740 703.790 1298.880 710.270 ;
        RECT 1298.680 703.470 1298.940 703.790 ;
        RECT 1298.220 655.530 1298.480 655.850 ;
        RECT 1298.280 638.510 1298.420 655.530 ;
        RECT 1297.300 638.190 1297.560 638.510 ;
        RECT 1298.220 638.190 1298.480 638.510 ;
        RECT 1297.360 614.565 1297.500 638.190 ;
        RECT 1297.290 614.195 1297.570 614.565 ;
        RECT 1298.210 614.195 1298.490 614.565 ;
        RECT 1298.280 607.230 1298.420 614.195 ;
        RECT 1298.220 606.910 1298.480 607.230 ;
        RECT 1299.140 558.970 1299.400 559.290 ;
        RECT 1299.200 542.630 1299.340 558.970 ;
        RECT 1298.220 542.310 1298.480 542.630 ;
        RECT 1299.140 542.310 1299.400 542.630 ;
        RECT 1298.280 517.470 1298.420 542.310 ;
        RECT 1298.220 517.150 1298.480 517.470 ;
        RECT 1298.220 493.350 1298.480 493.670 ;
        RECT 1298.280 434.850 1298.420 493.350 ;
        RECT 1298.220 434.530 1298.480 434.850 ;
        RECT 1298.680 434.530 1298.940 434.850 ;
        RECT 1298.740 380.110 1298.880 434.530 ;
        RECT 1298.680 379.790 1298.940 380.110 ;
        RECT 1298.220 372.650 1298.480 372.970 ;
        RECT 1298.280 331.490 1298.420 372.650 ;
        RECT 1298.220 331.170 1298.480 331.490 ;
        RECT 1298.220 324.370 1298.480 324.690 ;
        RECT 1298.280 269.010 1298.420 324.370 ;
        RECT 1298.280 268.870 1298.880 269.010 ;
        RECT 1298.740 210.530 1298.880 268.870 ;
        RECT 1298.740 210.390 1299.800 210.530 ;
        RECT 1299.660 192.850 1299.800 210.390 ;
        RECT 1299.200 192.710 1299.800 192.850 ;
        RECT 1299.200 145.170 1299.340 192.710 ;
        RECT 1298.680 144.850 1298.940 145.170 ;
        RECT 1299.140 144.850 1299.400 145.170 ;
        RECT 1298.740 62.290 1298.880 144.850 ;
        RECT 1298.280 62.150 1298.880 62.290 ;
        RECT 567.740 17.690 568.000 18.010 ;
        RECT 567.800 2.400 567.940 17.690 ;
        RECT 1298.280 15.290 1298.420 62.150 ;
        RECT 1298.220 14.970 1298.480 15.290 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 1298.670 1435.000 1298.950 1435.280 ;
        RECT 1299.590 1435.000 1299.870 1435.280 ;
        RECT 1297.290 910.720 1297.570 911.000 ;
        RECT 1298.670 910.720 1298.950 911.000 ;
        RECT 1298.210 820.960 1298.490 821.240 ;
        RECT 1299.130 820.960 1299.410 821.240 ;
        RECT 1297.290 614.240 1297.570 614.520 ;
        RECT 1298.210 614.240 1298.490 614.520 ;
      LAYER met3 ;
        RECT 1298.645 1435.290 1298.975 1435.305 ;
        RECT 1299.565 1435.290 1299.895 1435.305 ;
        RECT 1298.645 1434.990 1299.895 1435.290 ;
        RECT 1298.645 1434.975 1298.975 1434.990 ;
        RECT 1299.565 1434.975 1299.895 1434.990 ;
        RECT 1297.265 911.010 1297.595 911.025 ;
        RECT 1298.645 911.010 1298.975 911.025 ;
        RECT 1297.265 910.710 1298.975 911.010 ;
        RECT 1297.265 910.695 1297.595 910.710 ;
        RECT 1298.645 910.695 1298.975 910.710 ;
        RECT 1298.185 821.250 1298.515 821.265 ;
        RECT 1299.105 821.250 1299.435 821.265 ;
        RECT 1298.185 820.950 1299.435 821.250 ;
        RECT 1298.185 820.935 1298.515 820.950 ;
        RECT 1299.105 820.935 1299.435 820.950 ;
        RECT 1297.265 614.530 1297.595 614.545 ;
        RECT 1298.185 614.530 1298.515 614.545 ;
        RECT 1297.265 614.230 1298.515 614.530 ;
        RECT 1297.265 614.215 1297.595 614.230 ;
        RECT 1298.185 614.215 1298.515 614.230 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1294.050 1683.920 1294.370 1683.980 ;
        RECT 1303.710 1683.920 1304.030 1683.980 ;
        RECT 1294.050 1683.780 1304.030 1683.920 ;
        RECT 1294.050 1683.720 1294.370 1683.780 ;
        RECT 1303.710 1683.720 1304.030 1683.780 ;
        RECT 572.310 1624.760 572.630 1624.820 ;
        RECT 1294.050 1624.760 1294.370 1624.820 ;
        RECT 572.310 1624.620 1294.370 1624.760 ;
        RECT 572.310 1624.560 572.630 1624.620 ;
        RECT 1294.050 1624.560 1294.370 1624.620 ;
        RECT 567.710 14.860 568.030 14.920 ;
        RECT 572.310 14.860 572.630 14.920 ;
        RECT 567.710 14.720 572.630 14.860 ;
        RECT 567.710 14.660 568.030 14.720 ;
        RECT 572.310 14.660 572.630 14.720 ;
      LAYER via ;
        RECT 1294.080 1683.720 1294.340 1683.980 ;
        RECT 1303.740 1683.720 1304.000 1683.980 ;
        RECT 572.340 1624.560 572.600 1624.820 ;
        RECT 1294.080 1624.560 1294.340 1624.820 ;
        RECT 567.740 14.660 568.000 14.920 ;
        RECT 572.340 14.660 572.600 14.920 ;
      LAYER met2 ;
        RECT 1303.730 1700.000 1304.010 1704.000 ;
        RECT 1303.800 1684.010 1303.940 1700.000 ;
        RECT 1294.080 1683.690 1294.340 1684.010 ;
        RECT 1303.740 1683.690 1304.000 1684.010 ;
        RECT 1294.140 1624.850 1294.280 1683.690 ;
        RECT 572.340 1624.530 572.600 1624.850 ;
        RECT 1294.080 1624.530 1294.340 1624.850 ;
        RECT 572.400 14.950 572.540 1624.530 ;
        RECT 567.740 14.630 568.000 14.950 ;
        RECT 572.340 14.630 572.600 14.950 ;
        RECT 567.800 2.400 567.940 14.630 ;
        RECT 567.590 -4.800 568.150 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 0.300 ;
=======
      LAYER met1 ;
        RECT 927.890 1684.600 928.210 1684.660 ;
        RECT 1307.850 1684.600 1308.170 1684.660 ;
        RECT 927.890 1684.460 1308.170 1684.600 ;
        RECT 927.890 1684.400 928.210 1684.460 ;
        RECT 1307.850 1684.400 1308.170 1684.460 ;
        RECT 586.110 27.100 586.430 27.160 ;
        RECT 927.890 27.100 928.210 27.160 ;
        RECT 586.110 26.960 928.210 27.100 ;
        RECT 586.110 26.900 586.430 26.960 ;
        RECT 927.890 26.900 928.210 26.960 ;
      LAYER via ;
        RECT 927.920 1684.400 928.180 1684.660 ;
        RECT 1307.880 1684.400 1308.140 1684.660 ;
        RECT 586.140 26.900 586.400 27.160 ;
        RECT 927.920 26.900 928.180 27.160 ;
      LAYER met2 ;
        RECT 1307.870 1700.000 1308.150 1704.000 ;
        RECT 1307.940 1684.690 1308.080 1700.000 ;
        RECT 927.920 1684.370 928.180 1684.690 ;
        RECT 1307.880 1684.370 1308.140 1684.690 ;
        RECT 927.980 27.190 928.120 1684.370 ;
        RECT 586.140 26.870 586.400 27.190 ;
        RECT 927.920 26.870 928.180 27.190 ;
        RECT 586.200 14.010 586.340 26.870 ;
        RECT 585.740 13.870 586.340 14.010 ;
        RECT 585.740 2.400 585.880 13.870 ;
        RECT 585.530 -4.800 586.090 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1306.545 1110.525 1306.715 1152.175 ;
        RECT 1306.545 1007.165 1306.715 1048.815 ;
        RECT 1306.545 931.345 1306.715 1000.535 ;
        RECT 1306.545 766.105 1306.715 813.875 ;
        RECT 1306.545 641.325 1306.715 710.515 ;
        RECT 1307.005 591.685 1307.175 620.755 ;
        RECT 1307.005 113.645 1307.175 144.755 ;
      LAYER mcon ;
        RECT 1306.545 1152.005 1306.715 1152.175 ;
        RECT 1306.545 1048.645 1306.715 1048.815 ;
        RECT 1306.545 1000.365 1306.715 1000.535 ;
        RECT 1306.545 813.705 1306.715 813.875 ;
        RECT 1306.545 710.345 1306.715 710.515 ;
        RECT 1307.005 620.585 1307.175 620.755 ;
        RECT 1307.005 144.585 1307.175 144.755 ;
      LAYER met1 ;
        RECT 1306.930 1642.440 1307.250 1642.500 ;
        RECT 1307.850 1642.440 1308.170 1642.500 ;
        RECT 1306.930 1642.300 1308.170 1642.440 ;
        RECT 1306.930 1642.240 1307.250 1642.300 ;
        RECT 1307.850 1642.240 1308.170 1642.300 ;
        RECT 1306.470 1594.160 1306.790 1594.220 ;
        RECT 1306.930 1594.160 1307.250 1594.220 ;
        RECT 1306.470 1594.020 1307.250 1594.160 ;
        RECT 1306.470 1593.960 1306.790 1594.020 ;
        RECT 1306.930 1593.960 1307.250 1594.020 ;
        RECT 1306.930 1366.500 1307.250 1366.760 ;
        RECT 1307.020 1366.080 1307.160 1366.500 ;
        RECT 1306.930 1365.820 1307.250 1366.080 ;
        RECT 1306.470 1152.160 1306.790 1152.220 ;
        RECT 1306.275 1152.020 1306.790 1152.160 ;
        RECT 1306.470 1151.960 1306.790 1152.020 ;
        RECT 1306.485 1110.680 1306.775 1110.725 ;
        RECT 1306.930 1110.680 1307.250 1110.740 ;
        RECT 1306.485 1110.540 1307.250 1110.680 ;
        RECT 1306.485 1110.495 1306.775 1110.540 ;
        RECT 1306.930 1110.480 1307.250 1110.540 ;
        RECT 1306.470 1048.800 1306.790 1048.860 ;
        RECT 1306.275 1048.660 1306.790 1048.800 ;
        RECT 1306.470 1048.600 1306.790 1048.660 ;
        RECT 1306.470 1007.320 1306.790 1007.380 ;
        RECT 1306.275 1007.180 1306.790 1007.320 ;
        RECT 1306.470 1007.120 1306.790 1007.180 ;
        RECT 1306.470 1000.520 1306.790 1000.580 ;
        RECT 1306.275 1000.380 1306.790 1000.520 ;
        RECT 1306.470 1000.320 1306.790 1000.380 ;
        RECT 1306.470 931.500 1306.790 931.560 ;
        RECT 1306.275 931.360 1306.790 931.500 ;
        RECT 1306.470 931.300 1306.790 931.360 ;
        RECT 1306.930 883.900 1307.250 883.960 ;
        RECT 1306.100 883.760 1307.250 883.900 ;
        RECT 1306.100 883.620 1306.240 883.760 ;
        RECT 1306.930 883.700 1307.250 883.760 ;
        RECT 1306.010 883.360 1306.330 883.620 ;
        RECT 1305.090 862.480 1305.410 862.540 ;
        RECT 1306.010 862.480 1306.330 862.540 ;
        RECT 1305.090 862.340 1306.330 862.480 ;
        RECT 1305.090 862.280 1305.410 862.340 ;
        RECT 1306.010 862.280 1306.330 862.340 ;
        RECT 1306.470 813.860 1306.790 813.920 ;
        RECT 1306.275 813.720 1306.790 813.860 ;
        RECT 1306.470 813.660 1306.790 813.720 ;
        RECT 1306.470 766.260 1306.790 766.320 ;
        RECT 1306.275 766.120 1306.790 766.260 ;
        RECT 1306.470 766.060 1306.790 766.120 ;
        RECT 1306.470 710.500 1306.790 710.560 ;
        RECT 1306.275 710.360 1306.790 710.500 ;
        RECT 1306.470 710.300 1306.790 710.360 ;
        RECT 1306.470 641.480 1306.790 641.540 ;
        RECT 1306.275 641.340 1306.790 641.480 ;
        RECT 1306.470 641.280 1306.790 641.340 ;
        RECT 1306.930 620.740 1307.250 620.800 ;
        RECT 1306.735 620.600 1307.250 620.740 ;
        RECT 1306.930 620.540 1307.250 620.600 ;
        RECT 1306.930 591.840 1307.250 591.900 ;
        RECT 1306.735 591.700 1307.250 591.840 ;
        RECT 1306.930 591.640 1307.250 591.700 ;
        RECT 1306.470 337.860 1306.790 337.920 ;
        RECT 1306.930 337.860 1307.250 337.920 ;
        RECT 1306.470 337.720 1307.250 337.860 ;
        RECT 1306.470 337.660 1306.790 337.720 ;
        RECT 1306.930 337.660 1307.250 337.720 ;
        RECT 1306.930 144.740 1307.250 144.800 ;
        RECT 1306.735 144.600 1307.250 144.740 ;
        RECT 1306.930 144.540 1307.250 144.600 ;
        RECT 586.110 113.800 586.430 113.860 ;
        RECT 1306.945 113.800 1307.235 113.845 ;
        RECT 586.110 113.660 1307.235 113.800 ;
        RECT 586.110 113.600 586.430 113.660 ;
        RECT 1306.945 113.615 1307.235 113.660 ;
      LAYER via ;
        RECT 1306.960 1642.240 1307.220 1642.500 ;
        RECT 1307.880 1642.240 1308.140 1642.500 ;
        RECT 1306.500 1593.960 1306.760 1594.220 ;
        RECT 1306.960 1593.960 1307.220 1594.220 ;
        RECT 1306.960 1366.500 1307.220 1366.760 ;
        RECT 1306.960 1365.820 1307.220 1366.080 ;
        RECT 1306.500 1151.960 1306.760 1152.220 ;
        RECT 1306.960 1110.480 1307.220 1110.740 ;
        RECT 1306.500 1048.600 1306.760 1048.860 ;
        RECT 1306.500 1007.120 1306.760 1007.380 ;
        RECT 1306.500 1000.320 1306.760 1000.580 ;
        RECT 1306.500 931.300 1306.760 931.560 ;
        RECT 1306.960 883.700 1307.220 883.960 ;
        RECT 1306.040 883.360 1306.300 883.620 ;
        RECT 1305.120 862.280 1305.380 862.540 ;
        RECT 1306.040 862.280 1306.300 862.540 ;
        RECT 1306.500 813.660 1306.760 813.920 ;
        RECT 1306.500 766.060 1306.760 766.320 ;
        RECT 1306.500 710.300 1306.760 710.560 ;
        RECT 1306.500 641.280 1306.760 641.540 ;
        RECT 1306.960 620.540 1307.220 620.800 ;
        RECT 1306.960 591.640 1307.220 591.900 ;
        RECT 1306.500 337.660 1306.760 337.920 ;
        RECT 1306.960 337.660 1307.220 337.920 ;
        RECT 1306.960 144.540 1307.220 144.800 ;
        RECT 586.140 113.600 586.400 113.860 ;
      LAYER met2 ;
        RECT 1308.330 1700.410 1308.610 1704.000 ;
        RECT 1307.940 1700.270 1308.610 1700.410 ;
        RECT 1307.940 1642.530 1308.080 1700.270 ;
        RECT 1308.330 1700.000 1308.610 1700.270 ;
        RECT 1306.960 1642.210 1307.220 1642.530 ;
        RECT 1307.880 1642.210 1308.140 1642.530 ;
        RECT 1307.020 1594.250 1307.160 1642.210 ;
        RECT 1306.500 1593.930 1306.760 1594.250 ;
        RECT 1306.960 1593.930 1307.220 1594.250 ;
        RECT 1306.560 1593.650 1306.700 1593.930 ;
        RECT 1306.560 1593.510 1307.160 1593.650 ;
        RECT 1307.020 1463.090 1307.160 1593.510 ;
        RECT 1306.560 1462.950 1307.160 1463.090 ;
        RECT 1306.560 1462.410 1306.700 1462.950 ;
        RECT 1306.560 1462.270 1307.160 1462.410 ;
        RECT 1307.020 1366.790 1307.160 1462.270 ;
        RECT 1306.960 1366.470 1307.220 1366.790 ;
        RECT 1306.960 1365.790 1307.220 1366.110 ;
        RECT 1307.020 1269.970 1307.160 1365.790 ;
        RECT 1306.560 1269.830 1307.160 1269.970 ;
        RECT 1306.560 1269.290 1306.700 1269.830 ;
        RECT 1306.560 1269.150 1307.160 1269.290 ;
        RECT 1307.020 1173.410 1307.160 1269.150 ;
        RECT 1306.560 1173.270 1307.160 1173.410 ;
        RECT 1306.560 1152.250 1306.700 1173.270 ;
        RECT 1306.500 1151.930 1306.760 1152.250 ;
        RECT 1306.960 1110.450 1307.220 1110.770 ;
        RECT 1307.020 1055.770 1307.160 1110.450 ;
        RECT 1306.560 1055.630 1307.160 1055.770 ;
        RECT 1306.560 1048.890 1306.700 1055.630 ;
        RECT 1306.500 1048.570 1306.760 1048.890 ;
        RECT 1306.500 1007.090 1306.760 1007.410 ;
        RECT 1306.560 1000.610 1306.700 1007.090 ;
        RECT 1306.500 1000.290 1306.760 1000.610 ;
        RECT 1306.500 931.270 1306.760 931.590 ;
        RECT 1306.560 910.930 1306.700 931.270 ;
        RECT 1306.560 910.790 1307.160 910.930 ;
        RECT 1307.020 883.990 1307.160 910.790 ;
        RECT 1306.960 883.670 1307.220 883.990 ;
        RECT 1306.040 883.330 1306.300 883.650 ;
        RECT 1306.100 862.570 1306.240 883.330 ;
        RECT 1305.120 862.250 1305.380 862.570 ;
        RECT 1306.040 862.250 1306.300 862.570 ;
        RECT 1305.180 814.485 1305.320 862.250 ;
        RECT 1305.110 814.115 1305.390 814.485 ;
        RECT 1306.490 814.115 1306.770 814.485 ;
        RECT 1306.560 813.950 1306.700 814.115 ;
        RECT 1306.500 813.630 1306.760 813.950 ;
        RECT 1306.500 766.030 1306.760 766.350 ;
        RECT 1306.560 719.285 1306.700 766.030 ;
        RECT 1306.490 718.915 1306.770 719.285 ;
        RECT 1306.490 717.555 1306.770 717.925 ;
        RECT 1306.560 710.590 1306.700 717.555 ;
        RECT 1306.500 710.270 1306.760 710.590 ;
        RECT 1306.500 641.250 1306.760 641.570 ;
        RECT 1306.560 621.250 1306.700 641.250 ;
        RECT 1306.560 621.110 1307.160 621.250 ;
        RECT 1307.020 620.830 1307.160 621.110 ;
        RECT 1306.960 620.510 1307.220 620.830 ;
        RECT 1306.960 591.610 1307.220 591.930 ;
        RECT 1307.020 337.950 1307.160 591.610 ;
        RECT 1306.500 337.630 1306.760 337.950 ;
        RECT 1306.960 337.630 1307.220 337.950 ;
        RECT 1306.560 290.090 1306.700 337.630 ;
        RECT 1306.560 289.950 1307.160 290.090 ;
        RECT 1307.020 256.090 1307.160 289.950 ;
        RECT 1306.100 255.950 1307.160 256.090 ;
        RECT 1306.100 241.925 1306.240 255.950 ;
        RECT 1306.030 241.555 1306.310 241.925 ;
        RECT 1306.950 240.195 1307.230 240.565 ;
        RECT 1307.020 144.830 1307.160 240.195 ;
        RECT 1306.960 144.510 1307.220 144.830 ;
        RECT 586.140 113.570 586.400 113.890 ;
        RECT 586.200 17.410 586.340 113.570 ;
        RECT 585.740 17.270 586.340 17.410 ;
        RECT 585.740 2.400 585.880 17.270 ;
        RECT 585.530 -4.800 586.090 2.400 ;
      LAYER via2 ;
        RECT 1305.110 814.160 1305.390 814.440 ;
        RECT 1306.490 814.160 1306.770 814.440 ;
        RECT 1306.490 718.960 1306.770 719.240 ;
        RECT 1306.490 717.600 1306.770 717.880 ;
        RECT 1306.030 241.600 1306.310 241.880 ;
        RECT 1306.950 240.240 1307.230 240.520 ;
      LAYER met3 ;
        RECT 1305.085 814.450 1305.415 814.465 ;
        RECT 1306.465 814.450 1306.795 814.465 ;
        RECT 1305.085 814.150 1306.795 814.450 ;
        RECT 1305.085 814.135 1305.415 814.150 ;
        RECT 1306.465 814.135 1306.795 814.150 ;
        RECT 1306.465 719.250 1306.795 719.265 ;
        RECT 1306.465 718.935 1307.010 719.250 ;
        RECT 1306.710 717.905 1307.010 718.935 ;
        RECT 1306.465 717.590 1307.010 717.905 ;
        RECT 1306.465 717.575 1306.795 717.590 ;
        RECT 1306.005 241.890 1306.335 241.905 ;
        RECT 1305.790 241.575 1306.335 241.890 ;
        RECT 1305.790 240.530 1306.090 241.575 ;
        RECT 1306.925 240.530 1307.255 240.545 ;
        RECT 1305.790 240.230 1307.255 240.530 ;
        RECT 1306.925 240.215 1307.255 240.230 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 91.490 -4.800 92.050 0.300 ;
=======
        RECT 1174.470 1700.410 1174.750 1704.000 ;
        RECT 1173.160 1700.270 1174.750 1700.410 ;
        RECT 1173.160 19.565 1173.300 1700.270 ;
        RECT 1174.470 1700.000 1174.750 1700.270 ;
        RECT 91.630 19.195 91.910 19.565 ;
        RECT 1173.090 19.195 1173.370 19.565 ;
        RECT 91.700 2.400 91.840 19.195 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 91.630 19.240 91.910 19.520 ;
        RECT 1173.090 19.240 1173.370 19.520 ;
      LAYER met3 ;
        RECT 91.605 19.530 91.935 19.545 ;
        RECT 1173.065 19.530 1173.395 19.545 ;
        RECT 91.605 19.230 1173.395 19.530 ;
        RECT 91.605 19.215 91.935 19.230 ;
        RECT 1173.065 19.215 1173.395 19.230 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 99.890 1666.240 100.210 1666.300 ;
        RECT 1174.450 1666.240 1174.770 1666.300 ;
        RECT 99.890 1666.100 1174.770 1666.240 ;
        RECT 99.890 1666.040 100.210 1666.100 ;
        RECT 1174.450 1666.040 1174.770 1666.100 ;
        RECT 91.610 17.580 91.930 17.640 ;
        RECT 99.890 17.580 100.210 17.640 ;
        RECT 91.610 17.440 100.210 17.580 ;
        RECT 91.610 17.380 91.930 17.440 ;
        RECT 99.890 17.380 100.210 17.440 ;
      LAYER via ;
        RECT 99.920 1666.040 100.180 1666.300 ;
        RECT 1174.480 1666.040 1174.740 1666.300 ;
        RECT 91.640 17.380 91.900 17.640 ;
        RECT 99.920 17.380 100.180 17.640 ;
      LAYER met2 ;
        RECT 1174.470 1700.000 1174.750 1704.000 ;
        RECT 1174.540 1666.330 1174.680 1700.000 ;
        RECT 99.920 1666.010 100.180 1666.330 ;
        RECT 1174.480 1666.010 1174.740 1666.330 ;
        RECT 99.980 17.670 100.120 1666.010 ;
        RECT 91.640 17.350 91.900 17.670 ;
        RECT 99.920 17.350 100.180 17.670 ;
        RECT 91.700 2.400 91.840 17.350 ;
        RECT 91.490 -4.800 92.050 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 0.300 ;
=======
      LAYER met1 ;
        RECT 606.810 1500.660 607.130 1500.720 ;
        RECT 1312.450 1500.660 1312.770 1500.720 ;
        RECT 606.810 1500.520 1312.770 1500.660 ;
        RECT 606.810 1500.460 607.130 1500.520 ;
        RECT 1312.450 1500.460 1312.770 1500.520 ;
        RECT 603.130 14.860 603.450 14.920 ;
        RECT 606.810 14.860 607.130 14.920 ;
        RECT 603.130 14.720 607.130 14.860 ;
        RECT 603.130 14.660 603.450 14.720 ;
        RECT 606.810 14.660 607.130 14.720 ;
      LAYER via ;
        RECT 606.840 1500.460 607.100 1500.720 ;
        RECT 1312.480 1500.460 1312.740 1500.720 ;
        RECT 603.160 14.660 603.420 14.920 ;
        RECT 606.840 14.660 607.100 14.920 ;
      LAYER met2 ;
        RECT 1313.390 1700.410 1313.670 1704.000 ;
        RECT 1312.540 1700.270 1313.670 1700.410 ;
        RECT 1312.540 1500.750 1312.680 1700.270 ;
        RECT 1313.390 1700.000 1313.670 1700.270 ;
        RECT 606.840 1500.430 607.100 1500.750 ;
        RECT 1312.480 1500.430 1312.740 1500.750 ;
        RECT 606.900 14.950 607.040 1500.430 ;
        RECT 603.160 14.630 603.420 14.950 ;
        RECT 606.840 14.630 607.100 14.950 ;
        RECT 603.220 2.400 603.360 14.630 ;
        RECT 603.010 -4.800 603.570 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 0.300 ;
=======
      LAYER met1 ;
        RECT 627.050 1604.360 627.370 1604.420 ;
        RECT 1319.350 1604.360 1319.670 1604.420 ;
        RECT 627.050 1604.220 1319.670 1604.360 ;
        RECT 627.050 1604.160 627.370 1604.220 ;
        RECT 1319.350 1604.160 1319.670 1604.220 ;
        RECT 621.070 20.980 621.390 21.040 ;
        RECT 627.050 20.980 627.370 21.040 ;
        RECT 621.070 20.840 627.370 20.980 ;
        RECT 621.070 20.780 621.390 20.840 ;
        RECT 627.050 20.780 627.370 20.840 ;
      LAYER via ;
        RECT 627.080 1604.160 627.340 1604.420 ;
        RECT 1319.380 1604.160 1319.640 1604.420 ;
        RECT 621.100 20.780 621.360 21.040 ;
        RECT 627.080 20.780 627.340 21.040 ;
      LAYER met2 ;
        RECT 1317.990 1700.410 1318.270 1704.000 ;
        RECT 1317.990 1700.270 1319.580 1700.410 ;
        RECT 1317.990 1700.000 1318.270 1700.270 ;
        RECT 1319.440 1604.450 1319.580 1700.270 ;
        RECT 627.080 1604.130 627.340 1604.450 ;
        RECT 1319.380 1604.130 1319.640 1604.450 ;
        RECT 627.140 21.070 627.280 1604.130 ;
        RECT 621.100 20.750 621.360 21.070 ;
        RECT 627.080 20.750 627.340 21.070 ;
        RECT 621.160 2.400 621.300 20.750 ;
        RECT 620.950 -4.800 621.510 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 0.300 ;
=======
      LAYER met1 ;
        RECT 120.590 1617.960 120.910 1618.020 ;
        RECT 1181.350 1617.960 1181.670 1618.020 ;
        RECT 120.590 1617.820 1181.670 1617.960 ;
        RECT 120.590 1617.760 120.910 1617.820 ;
        RECT 1181.350 1617.760 1181.670 1617.820 ;
        RECT 115.530 17.580 115.850 17.640 ;
        RECT 120.590 17.580 120.910 17.640 ;
        RECT 115.530 17.440 120.910 17.580 ;
        RECT 115.530 17.380 115.850 17.440 ;
        RECT 120.590 17.380 120.910 17.440 ;
      LAYER via ;
        RECT 120.620 1617.760 120.880 1618.020 ;
        RECT 1181.380 1617.760 1181.640 1618.020 ;
        RECT 115.560 17.380 115.820 17.640 ;
        RECT 120.620 17.380 120.880 17.640 ;
      LAYER met2 ;
        RECT 1180.910 1700.000 1181.190 1704.000 ;
        RECT 1180.980 1666.410 1181.120 1700.000 ;
        RECT 1180.980 1666.270 1181.580 1666.410 ;
        RECT 1181.440 1618.050 1181.580 1666.270 ;
        RECT 120.620 1617.730 120.880 1618.050 ;
        RECT 1181.380 1617.730 1181.640 1618.050 ;
        RECT 120.680 17.670 120.820 1617.730 ;
        RECT 115.560 17.350 115.820 17.670 ;
        RECT 120.620 17.350 120.880 17.670 ;
        RECT 115.620 2.400 115.760 17.350 ;
        RECT 115.410 -4.800 115.970 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 0.300 ;
=======
      LAYER li1 ;
        RECT 276.145 16.405 276.315 18.275 ;
        RECT 323.985 16.405 324.155 18.275 ;
        RECT 372.745 15.385 372.915 18.275 ;
        RECT 420.585 15.385 420.755 18.275 ;
        RECT 469.345 15.045 469.515 18.275 ;
        RECT 517.185 15.045 517.355 18.275 ;
        RECT 565.945 15.045 566.115 18.275 ;
        RECT 599.525 14.875 599.695 15.215 ;
        RECT 599.525 14.705 601.535 14.875 ;
        RECT 613.785 14.705 613.955 18.275 ;
        RECT 662.545 18.105 662.715 21.335 ;
        RECT 709.925 20.995 710.095 21.335 ;
        RECT 709.925 20.825 710.555 20.995 ;
        RECT 710.385 18.105 710.555 20.825 ;
        RECT 759.145 18.105 759.315 21.335 ;
        RECT 806.985 18.105 807.155 21.335 ;
        RECT 855.745 18.105 855.915 20.995 ;
        RECT 903.585 18.105 903.755 20.995 ;
        RECT 952.345 18.105 952.515 20.995 ;
        RECT 1000.185 18.105 1000.355 20.995 ;
        RECT 1048.945 18.105 1049.115 20.995 ;
        RECT 1096.785 18.105 1096.955 20.995 ;
      LAYER mcon ;
        RECT 662.545 21.165 662.715 21.335 ;
        RECT 709.925 21.165 710.095 21.335 ;
        RECT 759.145 21.165 759.315 21.335 ;
        RECT 276.145 18.105 276.315 18.275 ;
        RECT 323.985 18.105 324.155 18.275 ;
        RECT 372.745 18.105 372.915 18.275 ;
        RECT 420.585 18.105 420.755 18.275 ;
        RECT 469.345 18.105 469.515 18.275 ;
        RECT 517.185 18.105 517.355 18.275 ;
        RECT 565.945 18.105 566.115 18.275 ;
        RECT 613.785 18.105 613.955 18.275 ;
        RECT 806.985 21.165 807.155 21.335 ;
        RECT 855.745 20.825 855.915 20.995 ;
        RECT 903.585 20.825 903.755 20.995 ;
        RECT 952.345 20.825 952.515 20.995 ;
        RECT 1000.185 20.825 1000.355 20.995 ;
        RECT 1048.945 20.825 1049.115 20.995 ;
        RECT 1096.785 20.825 1096.955 20.995 ;
        RECT 599.525 15.045 599.695 15.215 ;
        RECT 601.365 14.705 601.535 14.875 ;
      LAYER met1 ;
        RECT 662.485 21.320 662.775 21.365 ;
        RECT 709.865 21.320 710.155 21.365 ;
        RECT 662.485 21.180 710.155 21.320 ;
        RECT 662.485 21.135 662.775 21.180 ;
        RECT 709.865 21.135 710.155 21.180 ;
        RECT 759.085 21.320 759.375 21.365 ;
        RECT 806.925 21.320 807.215 21.365 ;
        RECT 759.085 21.180 807.215 21.320 ;
        RECT 759.085 21.135 759.375 21.180 ;
        RECT 806.925 21.135 807.215 21.180 ;
        RECT 855.685 20.980 855.975 21.025 ;
        RECT 903.525 20.980 903.815 21.025 ;
        RECT 855.685 20.840 903.815 20.980 ;
        RECT 855.685 20.795 855.975 20.840 ;
        RECT 903.525 20.795 903.815 20.840 ;
        RECT 952.285 20.980 952.575 21.025 ;
        RECT 1000.125 20.980 1000.415 21.025 ;
        RECT 952.285 20.840 1000.415 20.980 ;
        RECT 952.285 20.795 952.575 20.840 ;
        RECT 1000.125 20.795 1000.415 20.840 ;
        RECT 1048.885 20.980 1049.175 21.025 ;
        RECT 1096.725 20.980 1097.015 21.025 ;
        RECT 1048.885 20.840 1097.015 20.980 ;
        RECT 1048.885 20.795 1049.175 20.840 ;
        RECT 1096.725 20.795 1097.015 20.840 ;
        RECT 139.450 18.260 139.770 18.320 ;
        RECT 276.085 18.260 276.375 18.305 ;
        RECT 139.450 18.120 276.375 18.260 ;
        RECT 139.450 18.060 139.770 18.120 ;
        RECT 276.085 18.075 276.375 18.120 ;
        RECT 323.925 18.260 324.215 18.305 ;
        RECT 372.685 18.260 372.975 18.305 ;
        RECT 323.925 18.120 372.975 18.260 ;
        RECT 323.925 18.075 324.215 18.120 ;
        RECT 372.685 18.075 372.975 18.120 ;
        RECT 420.525 18.260 420.815 18.305 ;
        RECT 469.285 18.260 469.575 18.305 ;
        RECT 420.525 18.120 469.575 18.260 ;
        RECT 420.525 18.075 420.815 18.120 ;
        RECT 469.285 18.075 469.575 18.120 ;
        RECT 517.125 18.260 517.415 18.305 ;
        RECT 565.885 18.260 566.175 18.305 ;
        RECT 517.125 18.120 566.175 18.260 ;
        RECT 517.125 18.075 517.415 18.120 ;
        RECT 565.885 18.075 566.175 18.120 ;
        RECT 613.725 18.260 614.015 18.305 ;
        RECT 662.485 18.260 662.775 18.305 ;
        RECT 613.725 18.120 662.775 18.260 ;
        RECT 613.725 18.075 614.015 18.120 ;
        RECT 662.485 18.075 662.775 18.120 ;
        RECT 710.325 18.260 710.615 18.305 ;
        RECT 759.085 18.260 759.375 18.305 ;
        RECT 710.325 18.120 759.375 18.260 ;
        RECT 710.325 18.075 710.615 18.120 ;
        RECT 759.085 18.075 759.375 18.120 ;
        RECT 806.925 18.260 807.215 18.305 ;
        RECT 855.685 18.260 855.975 18.305 ;
        RECT 806.925 18.120 855.975 18.260 ;
        RECT 806.925 18.075 807.215 18.120 ;
        RECT 855.685 18.075 855.975 18.120 ;
        RECT 903.525 18.260 903.815 18.305 ;
        RECT 952.285 18.260 952.575 18.305 ;
        RECT 903.525 18.120 952.575 18.260 ;
        RECT 903.525 18.075 903.815 18.120 ;
        RECT 952.285 18.075 952.575 18.120 ;
        RECT 1000.125 18.260 1000.415 18.305 ;
        RECT 1048.885 18.260 1049.175 18.305 ;
        RECT 1000.125 18.120 1049.175 18.260 ;
        RECT 1000.125 18.075 1000.415 18.120 ;
        RECT 1048.885 18.075 1049.175 18.120 ;
        RECT 1096.725 18.260 1097.015 18.305 ;
        RECT 1186.870 18.260 1187.190 18.320 ;
        RECT 1096.725 18.120 1187.190 18.260 ;
        RECT 1096.725 18.075 1097.015 18.120 ;
        RECT 1186.870 18.060 1187.190 18.120 ;
        RECT 276.085 16.560 276.375 16.605 ;
        RECT 323.925 16.560 324.215 16.605 ;
        RECT 276.085 16.420 324.215 16.560 ;
        RECT 276.085 16.375 276.375 16.420 ;
        RECT 323.925 16.375 324.215 16.420 ;
        RECT 372.685 15.540 372.975 15.585 ;
        RECT 420.525 15.540 420.815 15.585 ;
        RECT 372.685 15.400 420.815 15.540 ;
        RECT 372.685 15.355 372.975 15.400 ;
        RECT 420.525 15.355 420.815 15.400 ;
        RECT 469.285 15.200 469.575 15.245 ;
        RECT 517.125 15.200 517.415 15.245 ;
        RECT 469.285 15.060 517.415 15.200 ;
        RECT 469.285 15.015 469.575 15.060 ;
        RECT 517.125 15.015 517.415 15.060 ;
        RECT 565.885 15.200 566.175 15.245 ;
        RECT 599.465 15.200 599.755 15.245 ;
        RECT 565.885 15.060 599.755 15.200 ;
        RECT 565.885 15.015 566.175 15.060 ;
        RECT 599.465 15.015 599.755 15.060 ;
        RECT 601.305 14.860 601.595 14.905 ;
        RECT 613.725 14.860 614.015 14.905 ;
        RECT 601.305 14.720 614.015 14.860 ;
        RECT 601.305 14.675 601.595 14.720 ;
        RECT 613.725 14.675 614.015 14.720 ;
      LAYER via ;
        RECT 139.480 18.060 139.740 18.320 ;
        RECT 1186.900 18.060 1187.160 18.320 ;
      LAYER met2 ;
        RECT 1187.350 1700.410 1187.630 1704.000 ;
        RECT 1186.960 1700.270 1187.630 1700.410 ;
        RECT 1186.960 18.350 1187.100 1700.270 ;
        RECT 1187.350 1700.000 1187.630 1700.270 ;
        RECT 139.480 18.030 139.740 18.350 ;
        RECT 1186.900 18.030 1187.160 18.350 ;
        RECT 139.540 2.400 139.680 18.030 ;
=======
      LAYER met1 ;
        RECT 155.090 1569.680 155.410 1569.740 ;
        RECT 1187.330 1569.680 1187.650 1569.740 ;
        RECT 155.090 1569.540 1187.650 1569.680 ;
        RECT 155.090 1569.480 155.410 1569.540 ;
        RECT 1187.330 1569.480 1187.650 1569.540 ;
        RECT 139.450 16.220 139.770 16.280 ;
        RECT 155.090 16.220 155.410 16.280 ;
        RECT 139.450 16.080 155.410 16.220 ;
        RECT 139.450 16.020 139.770 16.080 ;
        RECT 155.090 16.020 155.410 16.080 ;
      LAYER via ;
        RECT 155.120 1569.480 155.380 1569.740 ;
        RECT 1187.360 1569.480 1187.620 1569.740 ;
        RECT 139.480 16.020 139.740 16.280 ;
        RECT 155.120 16.020 155.380 16.280 ;
      LAYER met2 ;
        RECT 1187.350 1700.000 1187.630 1704.000 ;
        RECT 1187.420 1569.770 1187.560 1700.000 ;
        RECT 155.120 1569.450 155.380 1569.770 ;
        RECT 1187.360 1569.450 1187.620 1569.770 ;
        RECT 155.180 16.310 155.320 1569.450 ;
        RECT 139.480 15.990 139.740 16.310 ;
        RECT 155.120 15.990 155.380 16.310 ;
        RECT 139.540 2.400 139.680 15.990 ;
>>>>>>> re-updated local openlane
        RECT 139.330 -4.800 139.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 157.270 -4.800 157.830 0.300 ;
=======
        RECT 1191.950 1700.000 1192.230 1704.000 ;
        RECT 1192.020 1688.965 1192.160 1700.000 ;
        RECT 158.330 1688.595 158.610 1688.965 ;
        RECT 1191.950 1688.595 1192.230 1688.965 ;
        RECT 158.400 17.410 158.540 1688.595 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 158.330 1688.640 158.610 1688.920 ;
        RECT 1191.950 1688.640 1192.230 1688.920 ;
      LAYER met3 ;
        RECT 158.305 1688.930 158.635 1688.945 ;
        RECT 1191.925 1688.930 1192.255 1688.945 ;
        RECT 158.305 1688.630 1192.255 1688.930 ;
        RECT 158.305 1688.615 158.635 1688.630 ;
        RECT 1191.925 1688.615 1192.255 1688.630 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 1187.790 1656.380 1188.110 1656.440 ;
        RECT 1191.010 1656.380 1191.330 1656.440 ;
        RECT 1187.790 1656.240 1191.330 1656.380 ;
        RECT 1187.790 1656.180 1188.110 1656.240 ;
        RECT 1191.010 1656.180 1191.330 1656.240 ;
        RECT 162.450 1597.220 162.770 1597.280 ;
        RECT 1187.790 1597.220 1188.110 1597.280 ;
        RECT 162.450 1597.080 1188.110 1597.220 ;
        RECT 162.450 1597.020 162.770 1597.080 ;
        RECT 1187.790 1597.020 1188.110 1597.080 ;
        RECT 157.390 17.240 157.710 17.300 ;
        RECT 162.450 17.240 162.770 17.300 ;
        RECT 157.390 17.100 162.770 17.240 ;
        RECT 157.390 17.040 157.710 17.100 ;
        RECT 162.450 17.040 162.770 17.100 ;
      LAYER via ;
        RECT 1187.820 1656.180 1188.080 1656.440 ;
        RECT 1191.040 1656.180 1191.300 1656.440 ;
        RECT 162.480 1597.020 162.740 1597.280 ;
        RECT 1187.820 1597.020 1188.080 1597.280 ;
        RECT 157.420 17.040 157.680 17.300 ;
        RECT 162.480 17.040 162.740 17.300 ;
      LAYER met2 ;
        RECT 1192.410 1700.410 1192.690 1704.000 ;
        RECT 1191.100 1700.270 1192.690 1700.410 ;
        RECT 1191.100 1656.470 1191.240 1700.270 ;
        RECT 1192.410 1700.000 1192.690 1700.270 ;
        RECT 1187.820 1656.150 1188.080 1656.470 ;
        RECT 1191.040 1656.150 1191.300 1656.470 ;
        RECT 1187.880 1597.310 1188.020 1656.150 ;
        RECT 162.480 1596.990 162.740 1597.310 ;
        RECT 1187.820 1596.990 1188.080 1597.310 ;
        RECT 162.540 17.330 162.680 1596.990 ;
        RECT 157.420 17.010 157.680 17.330 ;
        RECT 162.480 17.010 162.740 17.330 ;
        RECT 157.480 2.400 157.620 17.010 ;
        RECT 157.270 -4.800 157.830 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 0.300 ;
=======
      LAYER met1 ;
        RECT 189.590 1645.500 189.910 1645.560 ;
        RECT 1195.150 1645.500 1195.470 1645.560 ;
        RECT 189.590 1645.360 1195.470 1645.500 ;
        RECT 189.590 1645.300 189.910 1645.360 ;
        RECT 1195.150 1645.300 1195.470 1645.360 ;
        RECT 174.870 20.300 175.190 20.360 ;
        RECT 189.590 20.300 189.910 20.360 ;
        RECT 174.870 20.160 189.910 20.300 ;
        RECT 174.870 20.100 175.190 20.160 ;
        RECT 189.590 20.100 189.910 20.160 ;
      LAYER via ;
        RECT 189.620 1645.300 189.880 1645.560 ;
        RECT 1195.180 1645.300 1195.440 1645.560 ;
        RECT 174.900 20.100 175.160 20.360 ;
        RECT 189.620 20.100 189.880 20.360 ;
      LAYER met2 ;
        RECT 1197.010 1700.410 1197.290 1704.000 ;
        RECT 1196.620 1700.270 1197.290 1700.410 ;
        RECT 1196.620 1667.090 1196.760 1700.270 ;
        RECT 1197.010 1700.000 1197.290 1700.270 ;
        RECT 1195.240 1666.950 1196.760 1667.090 ;
        RECT 1195.240 1645.590 1195.380 1666.950 ;
        RECT 189.620 1645.270 189.880 1645.590 ;
        RECT 1195.180 1645.270 1195.440 1645.590 ;
        RECT 189.680 20.390 189.820 1645.270 ;
        RECT 174.900 20.070 175.160 20.390 ;
        RECT 189.620 20.070 189.880 20.390 ;
        RECT 174.960 2.400 175.100 20.070 ;
        RECT 174.750 -4.800 175.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 0.300 ;
=======
      LAYER met1 ;
        RECT 192.810 1590.420 193.130 1590.480 ;
        RECT 1202.050 1590.420 1202.370 1590.480 ;
        RECT 192.810 1590.280 1202.370 1590.420 ;
        RECT 192.810 1590.220 193.130 1590.280 ;
        RECT 1202.050 1590.220 1202.370 1590.280 ;
      LAYER via ;
        RECT 192.840 1590.220 193.100 1590.480 ;
        RECT 1202.080 1590.220 1202.340 1590.480 ;
      LAYER met2 ;
        RECT 1202.070 1700.000 1202.350 1704.000 ;
        RECT 1202.140 1590.510 1202.280 1700.000 ;
        RECT 192.840 1590.190 193.100 1590.510 ;
        RECT 1202.080 1590.190 1202.340 1590.510 ;
        RECT 192.900 2.400 193.040 1590.190 ;
        RECT 192.690 -4.800 193.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 0.300 ;
=======
      LAYER li1 ;
        RECT 1201.665 786.505 1201.835 814.215 ;
        RECT 1201.665 524.365 1201.835 572.475 ;
        RECT 1202.125 276.165 1202.295 324.275 ;
        RECT 1202.125 179.605 1202.295 227.715 ;
        RECT 1202.125 65.365 1202.295 131.155 ;
      LAYER mcon ;
        RECT 1201.665 814.045 1201.835 814.215 ;
        RECT 1201.665 572.305 1201.835 572.475 ;
        RECT 1202.125 324.105 1202.295 324.275 ;
        RECT 1202.125 227.545 1202.295 227.715 ;
        RECT 1202.125 130.985 1202.295 131.155 ;
      LAYER met1 ;
        RECT 1202.050 1028.200 1202.370 1028.460 ;
        RECT 1202.140 1027.780 1202.280 1028.200 ;
        RECT 1202.050 1027.520 1202.370 1027.780 ;
        RECT 1202.510 1006.980 1202.830 1007.040 ;
        RECT 1204.350 1006.980 1204.670 1007.040 ;
        RECT 1202.510 1006.840 1204.670 1006.980 ;
        RECT 1202.510 1006.780 1202.830 1006.840 ;
        RECT 1204.350 1006.780 1204.670 1006.840 ;
        RECT 1202.050 869.420 1202.370 869.680 ;
        RECT 1202.140 868.940 1202.280 869.420 ;
        RECT 1202.510 868.940 1202.830 869.000 ;
        RECT 1202.140 868.800 1202.830 868.940 ;
        RECT 1202.510 868.740 1202.830 868.800 ;
        RECT 1201.590 845.480 1201.910 845.540 ;
        RECT 1202.510 845.480 1202.830 845.540 ;
        RECT 1201.590 845.340 1202.830 845.480 ;
        RECT 1201.590 845.280 1201.910 845.340 ;
        RECT 1202.510 845.280 1202.830 845.340 ;
        RECT 1201.590 814.200 1201.910 814.260 ;
        RECT 1201.395 814.060 1201.910 814.200 ;
        RECT 1201.590 814.000 1201.910 814.060 ;
        RECT 1201.590 786.660 1201.910 786.720 ;
        RECT 1201.395 786.520 1201.910 786.660 ;
        RECT 1201.590 786.460 1201.910 786.520 ;
        RECT 1201.605 572.460 1201.895 572.505 ;
        RECT 1202.050 572.460 1202.370 572.520 ;
        RECT 1201.605 572.320 1202.370 572.460 ;
        RECT 1201.605 572.275 1201.895 572.320 ;
        RECT 1202.050 572.260 1202.370 572.320 ;
        RECT 1201.590 524.520 1201.910 524.580 ;
        RECT 1201.395 524.380 1201.910 524.520 ;
        RECT 1201.590 524.320 1201.910 524.380 ;
        RECT 1201.590 427.620 1201.910 427.680 ;
        RECT 1202.050 427.620 1202.370 427.680 ;
        RECT 1201.590 427.480 1202.370 427.620 ;
        RECT 1201.590 427.420 1201.910 427.480 ;
        RECT 1202.050 427.420 1202.370 427.480 ;
        RECT 1201.590 331.060 1201.910 331.120 ;
        RECT 1202.050 331.060 1202.370 331.120 ;
        RECT 1201.590 330.920 1202.370 331.060 ;
        RECT 1201.590 330.860 1201.910 330.920 ;
        RECT 1202.050 330.860 1202.370 330.920 ;
        RECT 1202.050 324.260 1202.370 324.320 ;
        RECT 1201.855 324.120 1202.370 324.260 ;
        RECT 1202.050 324.060 1202.370 324.120 ;
        RECT 1202.050 276.320 1202.370 276.380 ;
        RECT 1201.855 276.180 1202.370 276.320 ;
        RECT 1202.050 276.120 1202.370 276.180 ;
        RECT 1201.590 234.300 1201.910 234.560 ;
        RECT 1201.680 234.160 1201.820 234.300 ;
        RECT 1202.050 234.160 1202.370 234.220 ;
        RECT 1201.680 234.020 1202.370 234.160 ;
        RECT 1202.050 233.960 1202.370 234.020 ;
        RECT 1202.050 227.700 1202.370 227.760 ;
        RECT 1201.855 227.560 1202.370 227.700 ;
        RECT 1202.050 227.500 1202.370 227.560 ;
        RECT 1202.050 179.760 1202.370 179.820 ;
        RECT 1201.855 179.620 1202.370 179.760 ;
        RECT 1202.050 179.560 1202.370 179.620 ;
        RECT 1201.590 131.140 1201.910 131.200 ;
        RECT 1202.065 131.140 1202.355 131.185 ;
        RECT 1201.590 131.000 1202.355 131.140 ;
        RECT 1201.590 130.940 1201.910 131.000 ;
        RECT 1202.065 130.955 1202.355 131.000 ;
        RECT 1202.065 65.520 1202.355 65.565 ;
        RECT 1202.970 65.520 1203.290 65.580 ;
        RECT 1202.065 65.380 1203.290 65.520 ;
        RECT 1202.065 65.335 1202.355 65.380 ;
        RECT 1202.970 65.320 1203.290 65.380 ;
        RECT 210.750 19.620 211.070 19.680 ;
        RECT 1201.590 19.620 1201.910 19.680 ;
        RECT 210.750 19.480 1201.910 19.620 ;
        RECT 210.750 19.420 211.070 19.480 ;
        RECT 1201.590 19.420 1201.910 19.480 ;
      LAYER via ;
        RECT 1202.080 1028.200 1202.340 1028.460 ;
        RECT 1202.080 1027.520 1202.340 1027.780 ;
        RECT 1202.540 1006.780 1202.800 1007.040 ;
        RECT 1204.380 1006.780 1204.640 1007.040 ;
        RECT 1202.080 869.420 1202.340 869.680 ;
        RECT 1202.540 868.740 1202.800 869.000 ;
        RECT 1201.620 845.280 1201.880 845.540 ;
        RECT 1202.540 845.280 1202.800 845.540 ;
        RECT 1201.620 814.000 1201.880 814.260 ;
        RECT 1201.620 786.460 1201.880 786.720 ;
        RECT 1202.080 572.260 1202.340 572.520 ;
        RECT 1201.620 524.320 1201.880 524.580 ;
        RECT 1201.620 427.420 1201.880 427.680 ;
        RECT 1202.080 427.420 1202.340 427.680 ;
        RECT 1201.620 330.860 1201.880 331.120 ;
        RECT 1202.080 330.860 1202.340 331.120 ;
        RECT 1202.080 324.060 1202.340 324.320 ;
        RECT 1202.080 276.120 1202.340 276.380 ;
        RECT 1201.620 234.300 1201.880 234.560 ;
        RECT 1202.080 233.960 1202.340 234.220 ;
        RECT 1202.080 227.500 1202.340 227.760 ;
        RECT 1202.080 179.560 1202.340 179.820 ;
        RECT 1201.620 130.940 1201.880 131.200 ;
        RECT 1203.000 65.320 1203.260 65.580 ;
        RECT 210.780 19.420 211.040 19.680 ;
        RECT 1201.620 19.420 1201.880 19.680 ;
=======
      LAYER met1 ;
        RECT 1201.590 1667.600 1201.910 1667.660 ;
        RECT 1205.730 1667.600 1206.050 1667.660 ;
        RECT 1201.590 1667.460 1206.050 1667.600 ;
        RECT 1201.590 1667.400 1201.910 1667.460 ;
        RECT 1205.730 1667.400 1206.050 1667.460 ;
        RECT 217.190 1479.920 217.510 1479.980 ;
        RECT 1201.590 1479.920 1201.910 1479.980 ;
        RECT 217.190 1479.780 1201.910 1479.920 ;
        RECT 217.190 1479.720 217.510 1479.780 ;
        RECT 1201.590 1479.720 1201.910 1479.780 ;
        RECT 210.750 17.580 211.070 17.640 ;
        RECT 217.190 17.580 217.510 17.640 ;
        RECT 210.750 17.440 217.510 17.580 ;
        RECT 210.750 17.380 211.070 17.440 ;
        RECT 217.190 17.380 217.510 17.440 ;
      LAYER via ;
        RECT 1201.620 1667.400 1201.880 1667.660 ;
        RECT 1205.760 1667.400 1206.020 1667.660 ;
        RECT 217.220 1479.720 217.480 1479.980 ;
        RECT 1201.620 1479.720 1201.880 1479.980 ;
        RECT 210.780 17.380 211.040 17.640 ;
        RECT 217.220 17.380 217.480 17.640 ;
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1206.670 1700.410 1206.950 1704.000 ;
        RECT 1205.820 1700.270 1206.950 1700.410 ;
        RECT 1205.820 1667.690 1205.960 1700.270 ;
        RECT 1206.670 1700.000 1206.950 1700.270 ;
        RECT 1201.620 1667.370 1201.880 1667.690 ;
        RECT 1205.760 1667.370 1206.020 1667.690 ;
        RECT 1201.680 1480.010 1201.820 1667.370 ;
        RECT 217.220 1479.690 217.480 1480.010 ;
        RECT 1201.620 1479.690 1201.880 1480.010 ;
        RECT 217.280 17.670 217.420 1479.690 ;
        RECT 210.780 17.350 211.040 17.670 ;
        RECT 217.220 17.350 217.480 17.670 ;
        RECT 210.840 2.400 210.980 17.350 ;
        RECT 210.630 -4.800 211.190 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 1203.450 959.000 1203.730 959.280 ;
        RECT 1204.370 959.000 1204.650 959.280 ;
        RECT 1202.070 910.720 1202.350 911.000 ;
        RECT 1203.450 910.720 1203.730 911.000 ;
        RECT 1202.070 628.520 1202.350 628.800 ;
        RECT 1201.610 627.840 1201.890 628.120 ;
        RECT 1202.070 435.400 1202.350 435.680 ;
        RECT 1201.610 434.720 1201.890 435.000 ;
        RECT 1202.070 41.680 1202.350 41.960 ;
        RECT 1202.990 41.680 1203.270 41.960 ;
      LAYER met3 ;
        RECT 1203.425 959.290 1203.755 959.305 ;
        RECT 1204.345 959.290 1204.675 959.305 ;
        RECT 1203.425 958.990 1204.675 959.290 ;
        RECT 1203.425 958.975 1203.755 958.990 ;
        RECT 1204.345 958.975 1204.675 958.990 ;
        RECT 1202.045 911.010 1202.375 911.025 ;
        RECT 1203.425 911.010 1203.755 911.025 ;
        RECT 1202.045 910.710 1203.755 911.010 ;
        RECT 1202.045 910.695 1202.375 910.710 ;
        RECT 1203.425 910.695 1203.755 910.710 ;
        RECT 1202.045 628.810 1202.375 628.825 ;
        RECT 1201.830 628.495 1202.375 628.810 ;
        RECT 1201.830 628.145 1202.130 628.495 ;
        RECT 1201.585 627.830 1202.130 628.145 ;
        RECT 1201.585 627.815 1201.915 627.830 ;
        RECT 1202.045 435.690 1202.375 435.705 ;
        RECT 1201.830 435.375 1202.375 435.690 ;
        RECT 1201.830 435.025 1202.130 435.375 ;
        RECT 1201.585 434.710 1202.130 435.025 ;
        RECT 1201.585 434.695 1201.915 434.710 ;
        RECT 1202.045 41.970 1202.375 41.985 ;
        RECT 1202.965 41.970 1203.295 41.985 ;
        RECT 1202.045 41.670 1203.295 41.970 ;
        RECT 1202.045 41.655 1202.375 41.670 ;
        RECT 1202.965 41.655 1203.295 41.670 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 0.300 ;
=======
      LAYER li1 ;
        RECT 1186.945 1687.165 1187.115 1689.035 ;
      LAYER mcon ;
        RECT 1186.945 1688.865 1187.115 1689.035 ;
      LAYER met1 ;
        RECT 1186.885 1689.020 1187.175 1689.065 ;
        RECT 1211.250 1689.020 1211.570 1689.080 ;
        RECT 1186.885 1688.880 1211.570 1689.020 ;
        RECT 1186.885 1688.835 1187.175 1688.880 ;
        RECT 1211.250 1688.820 1211.570 1688.880 ;
        RECT 234.210 1687.320 234.530 1687.380 ;
        RECT 1186.885 1687.320 1187.175 1687.365 ;
        RECT 234.210 1687.180 1187.175 1687.320 ;
        RECT 234.210 1687.120 234.530 1687.180 ;
        RECT 1186.885 1687.135 1187.175 1687.180 ;
        RECT 228.690 16.900 229.010 16.960 ;
        RECT 234.210 16.900 234.530 16.960 ;
        RECT 228.690 16.760 234.530 16.900 ;
        RECT 228.690 16.700 229.010 16.760 ;
        RECT 234.210 16.700 234.530 16.760 ;
      LAYER via ;
        RECT 1211.280 1688.820 1211.540 1689.080 ;
        RECT 234.240 1687.120 234.500 1687.380 ;
        RECT 228.720 16.700 228.980 16.960 ;
        RECT 234.240 16.700 234.500 16.960 ;
      LAYER met2 ;
        RECT 1211.270 1700.000 1211.550 1704.000 ;
        RECT 1211.340 1689.110 1211.480 1700.000 ;
        RECT 1211.280 1688.790 1211.540 1689.110 ;
        RECT 234.240 1687.090 234.500 1687.410 ;
        RECT 234.300 16.990 234.440 1687.090 ;
        RECT 228.720 16.670 228.980 16.990 ;
        RECT 234.240 16.670 234.500 16.990 ;
        RECT 228.780 2.400 228.920 16.670 ;
=======
      LAYER met1 ;
        RECT 1190.090 1683.920 1190.410 1683.980 ;
        RECT 1211.710 1683.920 1212.030 1683.980 ;
        RECT 1190.090 1683.780 1212.030 1683.920 ;
        RECT 1190.090 1683.720 1190.410 1683.780 ;
        RECT 1211.710 1683.720 1212.030 1683.780 ;
        RECT 234.210 1487.060 234.530 1487.120 ;
        RECT 1190.090 1487.060 1190.410 1487.120 ;
        RECT 234.210 1486.920 1190.410 1487.060 ;
        RECT 234.210 1486.860 234.530 1486.920 ;
        RECT 1190.090 1486.860 1190.410 1486.920 ;
        RECT 228.690 17.580 229.010 17.640 ;
        RECT 234.210 17.580 234.530 17.640 ;
        RECT 228.690 17.440 234.530 17.580 ;
        RECT 228.690 17.380 229.010 17.440 ;
        RECT 234.210 17.380 234.530 17.440 ;
      LAYER via ;
        RECT 1190.120 1683.720 1190.380 1683.980 ;
        RECT 1211.740 1683.720 1212.000 1683.980 ;
        RECT 234.240 1486.860 234.500 1487.120 ;
        RECT 1190.120 1486.860 1190.380 1487.120 ;
        RECT 228.720 17.380 228.980 17.640 ;
        RECT 234.240 17.380 234.500 17.640 ;
      LAYER met2 ;
        RECT 1211.730 1700.000 1212.010 1704.000 ;
        RECT 1211.800 1684.010 1211.940 1700.000 ;
        RECT 1190.120 1683.690 1190.380 1684.010 ;
        RECT 1211.740 1683.690 1212.000 1684.010 ;
        RECT 1190.180 1487.150 1190.320 1683.690 ;
        RECT 234.240 1486.830 234.500 1487.150 ;
        RECT 1190.120 1486.830 1190.380 1487.150 ;
        RECT 234.300 17.670 234.440 1486.830 ;
        RECT 228.720 17.350 228.980 17.670 ;
        RECT 234.240 17.350 234.500 17.670 ;
        RECT 228.780 2.400 228.920 17.350 ;
>>>>>>> re-updated local openlane
        RECT 228.570 -4.800 229.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 0.300 ;
=======
      LAYER li1 ;
        RECT 1162.105 1538.925 1162.275 1587.035 ;
        RECT 1161.185 1497.445 1161.355 1511.555 ;
        RECT 1161.185 1442.025 1161.355 1490.475 ;
        RECT 1161.645 966.365 1161.815 980.135 ;
        RECT 1161.645 303.365 1161.815 337.875 ;
      LAYER mcon ;
        RECT 1162.105 1586.865 1162.275 1587.035 ;
        RECT 1161.185 1511.385 1161.355 1511.555 ;
        RECT 1161.185 1490.305 1161.355 1490.475 ;
        RECT 1161.645 979.965 1161.815 980.135 ;
        RECT 1161.645 337.705 1161.815 337.875 ;
      LAYER met1 ;
        RECT 1161.570 1607.900 1161.890 1608.160 ;
        RECT 1161.660 1607.420 1161.800 1607.900 ;
        RECT 1162.030 1607.420 1162.350 1607.480 ;
        RECT 1161.660 1607.280 1162.350 1607.420 ;
        RECT 1162.030 1607.220 1162.350 1607.280 ;
        RECT 1162.045 1587.020 1162.335 1587.065 ;
        RECT 1162.490 1587.020 1162.810 1587.080 ;
        RECT 1162.045 1586.880 1162.810 1587.020 ;
        RECT 1162.045 1586.835 1162.335 1586.880 ;
        RECT 1162.490 1586.820 1162.810 1586.880 ;
        RECT 1162.030 1539.080 1162.350 1539.140 ;
        RECT 1161.835 1538.940 1162.350 1539.080 ;
        RECT 1162.030 1538.880 1162.350 1538.940 ;
        RECT 1161.125 1511.540 1161.415 1511.585 ;
        RECT 1162.030 1511.540 1162.350 1511.600 ;
        RECT 1161.125 1511.400 1162.350 1511.540 ;
        RECT 1161.125 1511.355 1161.415 1511.400 ;
        RECT 1162.030 1511.340 1162.350 1511.400 ;
        RECT 1161.110 1497.600 1161.430 1497.660 ;
        RECT 1160.915 1497.460 1161.430 1497.600 ;
        RECT 1161.110 1497.400 1161.430 1497.460 ;
        RECT 1161.110 1490.460 1161.430 1490.520 ;
        RECT 1160.915 1490.320 1161.430 1490.460 ;
        RECT 1161.110 1490.260 1161.430 1490.320 ;
        RECT 1161.125 1442.180 1161.415 1442.225 ;
        RECT 1162.490 1442.180 1162.810 1442.240 ;
        RECT 1161.125 1442.040 1162.810 1442.180 ;
        RECT 1161.125 1441.995 1161.415 1442.040 ;
        RECT 1162.490 1441.980 1162.810 1442.040 ;
        RECT 1162.030 1345.620 1162.350 1345.680 ;
        RECT 1162.490 1345.620 1162.810 1345.680 ;
        RECT 1162.030 1345.480 1162.810 1345.620 ;
        RECT 1162.030 1345.420 1162.350 1345.480 ;
        RECT 1162.490 1345.420 1162.810 1345.480 ;
        RECT 1161.570 1304.820 1161.890 1304.880 ;
        RECT 1162.030 1304.820 1162.350 1304.880 ;
        RECT 1161.570 1304.680 1162.350 1304.820 ;
        RECT 1161.570 1304.620 1161.890 1304.680 ;
        RECT 1162.030 1304.620 1162.350 1304.680 ;
        RECT 1161.570 1304.140 1161.890 1304.200 ;
        RECT 1162.030 1304.140 1162.350 1304.200 ;
        RECT 1161.570 1304.000 1162.350 1304.140 ;
        RECT 1161.570 1303.940 1161.890 1304.000 ;
        RECT 1162.030 1303.940 1162.350 1304.000 ;
        RECT 1161.570 1159.300 1161.890 1159.360 ;
        RECT 1162.030 1159.300 1162.350 1159.360 ;
        RECT 1161.570 1159.160 1162.350 1159.300 ;
        RECT 1161.570 1159.100 1161.890 1159.160 ;
        RECT 1162.030 1159.100 1162.350 1159.160 ;
        RECT 1161.570 1062.740 1161.890 1062.800 ;
        RECT 1162.030 1062.740 1162.350 1062.800 ;
        RECT 1161.570 1062.600 1162.350 1062.740 ;
        RECT 1161.570 1062.540 1161.890 1062.600 ;
        RECT 1162.030 1062.540 1162.350 1062.600 ;
        RECT 1161.570 980.120 1161.890 980.180 ;
        RECT 1161.375 979.980 1161.890 980.120 ;
        RECT 1161.570 979.920 1161.890 979.980 ;
        RECT 1161.570 966.520 1161.890 966.580 ;
        RECT 1161.375 966.380 1161.890 966.520 ;
        RECT 1161.570 966.320 1161.890 966.380 ;
        RECT 1161.570 931.980 1161.890 932.240 ;
        RECT 1161.660 931.560 1161.800 931.980 ;
        RECT 1161.570 931.300 1161.890 931.560 ;
        RECT 1161.570 869.620 1161.890 869.680 ;
        RECT 1162.030 869.620 1162.350 869.680 ;
        RECT 1161.570 869.480 1162.350 869.620 ;
        RECT 1161.570 869.420 1161.890 869.480 ;
        RECT 1162.030 869.420 1162.350 869.480 ;
        RECT 1161.110 786.660 1161.430 786.720 ;
        RECT 1162.030 786.660 1162.350 786.720 ;
        RECT 1161.110 786.520 1162.350 786.660 ;
        RECT 1161.110 786.460 1161.430 786.520 ;
        RECT 1162.030 786.460 1162.350 786.520 ;
        RECT 1161.570 689.900 1161.890 690.160 ;
        RECT 1161.660 689.760 1161.800 689.900 ;
        RECT 1162.030 689.760 1162.350 689.820 ;
        RECT 1161.660 689.620 1162.350 689.760 ;
        RECT 1162.030 689.560 1162.350 689.620 ;
        RECT 1161.570 593.340 1161.890 593.600 ;
        RECT 1161.660 593.200 1161.800 593.340 ;
        RECT 1162.030 593.200 1162.350 593.260 ;
        RECT 1161.660 593.060 1162.350 593.200 ;
        RECT 1162.030 593.000 1162.350 593.060 ;
        RECT 1161.570 517.380 1161.890 517.440 ;
        RECT 1162.030 517.380 1162.350 517.440 ;
        RECT 1161.570 517.240 1162.350 517.380 ;
        RECT 1161.570 517.180 1161.890 517.240 ;
        RECT 1162.030 517.180 1162.350 517.240 ;
        RECT 1161.570 337.860 1161.890 337.920 ;
        RECT 1161.375 337.720 1161.890 337.860 ;
        RECT 1161.570 337.660 1161.890 337.720 ;
        RECT 1161.570 303.520 1161.890 303.580 ;
        RECT 1161.375 303.380 1161.890 303.520 ;
        RECT 1161.570 303.320 1161.890 303.380 ;
      LAYER via ;
        RECT 1161.600 1607.900 1161.860 1608.160 ;
        RECT 1162.060 1607.220 1162.320 1607.480 ;
        RECT 1162.520 1586.820 1162.780 1587.080 ;
        RECT 1162.060 1538.880 1162.320 1539.140 ;
        RECT 1162.060 1511.340 1162.320 1511.600 ;
        RECT 1161.140 1497.400 1161.400 1497.660 ;
        RECT 1161.140 1490.260 1161.400 1490.520 ;
        RECT 1162.520 1441.980 1162.780 1442.240 ;
        RECT 1162.060 1345.420 1162.320 1345.680 ;
        RECT 1162.520 1345.420 1162.780 1345.680 ;
        RECT 1161.600 1304.620 1161.860 1304.880 ;
        RECT 1162.060 1304.620 1162.320 1304.880 ;
        RECT 1161.600 1303.940 1161.860 1304.200 ;
        RECT 1162.060 1303.940 1162.320 1304.200 ;
        RECT 1161.600 1159.100 1161.860 1159.360 ;
        RECT 1162.060 1159.100 1162.320 1159.360 ;
        RECT 1161.600 1062.540 1161.860 1062.800 ;
        RECT 1162.060 1062.540 1162.320 1062.800 ;
        RECT 1161.600 979.920 1161.860 980.180 ;
        RECT 1161.600 966.320 1161.860 966.580 ;
        RECT 1161.600 931.980 1161.860 932.240 ;
        RECT 1161.600 931.300 1161.860 931.560 ;
        RECT 1161.600 869.420 1161.860 869.680 ;
        RECT 1162.060 869.420 1162.320 869.680 ;
        RECT 1161.140 786.460 1161.400 786.720 ;
        RECT 1162.060 786.460 1162.320 786.720 ;
        RECT 1161.600 689.900 1161.860 690.160 ;
        RECT 1162.060 689.560 1162.320 689.820 ;
        RECT 1161.600 593.340 1161.860 593.600 ;
        RECT 1162.060 593.000 1162.320 593.260 ;
        RECT 1161.600 517.180 1161.860 517.440 ;
        RECT 1162.060 517.180 1162.320 517.440 ;
        RECT 1161.600 337.660 1161.860 337.920 ;
        RECT 1161.600 303.320 1161.860 303.580 ;
      LAYER met2 ;
        RECT 1162.970 1700.410 1163.250 1704.000 ;
        RECT 1162.580 1700.270 1163.250 1700.410 ;
        RECT 1162.580 1688.850 1162.720 1700.270 ;
        RECT 1162.970 1700.000 1163.250 1700.270 ;
        RECT 1161.660 1688.710 1162.720 1688.850 ;
        RECT 1161.660 1608.190 1161.800 1688.710 ;
        RECT 1161.600 1607.870 1161.860 1608.190 ;
        RECT 1162.060 1607.190 1162.320 1607.510 ;
        RECT 1162.120 1594.330 1162.260 1607.190 ;
        RECT 1162.120 1594.190 1162.720 1594.330 ;
        RECT 1162.580 1587.110 1162.720 1594.190 ;
        RECT 1162.520 1586.790 1162.780 1587.110 ;
        RECT 1162.060 1538.850 1162.320 1539.170 ;
        RECT 1162.120 1511.630 1162.260 1538.850 ;
        RECT 1162.060 1511.310 1162.320 1511.630 ;
        RECT 1161.140 1497.370 1161.400 1497.690 ;
        RECT 1161.200 1490.550 1161.340 1497.370 ;
        RECT 1161.140 1490.230 1161.400 1490.550 ;
        RECT 1162.520 1441.950 1162.780 1442.270 ;
        RECT 1162.580 1345.710 1162.720 1441.950 ;
        RECT 1162.060 1345.390 1162.320 1345.710 ;
        RECT 1162.520 1345.390 1162.780 1345.710 ;
        RECT 1162.120 1304.910 1162.260 1345.390 ;
        RECT 1161.600 1304.590 1161.860 1304.910 ;
        RECT 1162.060 1304.590 1162.320 1304.910 ;
        RECT 1161.660 1304.230 1161.800 1304.590 ;
        RECT 1161.600 1303.910 1161.860 1304.230 ;
        RECT 1162.060 1303.910 1162.320 1304.230 ;
        RECT 1162.120 1221.010 1162.260 1303.910 ;
        RECT 1161.660 1220.870 1162.260 1221.010 ;
        RECT 1161.660 1159.390 1161.800 1220.870 ;
        RECT 1161.600 1159.070 1161.860 1159.390 ;
        RECT 1162.060 1159.070 1162.320 1159.390 ;
        RECT 1162.120 1124.450 1162.260 1159.070 ;
        RECT 1161.660 1124.310 1162.260 1124.450 ;
        RECT 1161.660 1062.830 1161.800 1124.310 ;
        RECT 1161.600 1062.510 1161.860 1062.830 ;
        RECT 1162.060 1062.510 1162.320 1062.830 ;
        RECT 1162.120 1027.890 1162.260 1062.510 ;
        RECT 1161.660 1027.750 1162.260 1027.890 ;
        RECT 1161.660 980.210 1161.800 1027.750 ;
        RECT 1161.600 979.890 1161.860 980.210 ;
        RECT 1161.600 966.290 1161.860 966.610 ;
        RECT 1161.660 932.270 1161.800 966.290 ;
        RECT 1161.600 931.950 1161.860 932.270 ;
        RECT 1161.600 931.270 1161.860 931.590 ;
        RECT 1161.660 869.710 1161.800 931.270 ;
        RECT 1161.600 869.390 1161.860 869.710 ;
        RECT 1162.060 869.390 1162.320 869.710 ;
        RECT 1162.120 845.650 1162.260 869.390 ;
        RECT 1161.660 845.510 1162.260 845.650 ;
        RECT 1161.660 787.170 1161.800 845.510 ;
        RECT 1161.200 787.030 1161.800 787.170 ;
        RECT 1161.200 786.750 1161.340 787.030 ;
        RECT 1161.140 786.430 1161.400 786.750 ;
        RECT 1162.060 786.430 1162.320 786.750 ;
        RECT 1162.120 725.405 1162.260 786.430 ;
        RECT 1162.050 725.035 1162.330 725.405 ;
        RECT 1161.590 724.355 1161.870 724.725 ;
        RECT 1161.660 690.190 1161.800 724.355 ;
        RECT 1161.600 689.870 1161.860 690.190 ;
        RECT 1162.060 689.530 1162.320 689.850 ;
        RECT 1162.120 641.650 1162.260 689.530 ;
        RECT 1161.660 641.510 1162.260 641.650 ;
        RECT 1161.660 593.630 1161.800 641.510 ;
        RECT 1161.600 593.310 1161.860 593.630 ;
        RECT 1162.060 592.970 1162.320 593.290 ;
        RECT 1162.120 545.090 1162.260 592.970 ;
        RECT 1161.660 544.950 1162.260 545.090 ;
        RECT 1161.660 517.470 1161.800 544.950 ;
        RECT 1161.600 517.150 1161.860 517.470 ;
        RECT 1162.060 517.150 1162.320 517.470 ;
        RECT 1162.120 362.170 1162.260 517.150 ;
        RECT 1161.660 362.030 1162.260 362.170 ;
        RECT 1161.660 337.950 1161.800 362.030 ;
        RECT 1161.600 337.630 1161.860 337.950 ;
        RECT 1161.600 303.290 1161.860 303.610 ;
        RECT 1161.660 265.610 1161.800 303.290 ;
        RECT 1161.200 265.470 1161.800 265.610 ;
        RECT 1161.200 254.730 1161.340 265.470 ;
        RECT 1161.200 254.590 1162.260 254.730 ;
        RECT 1162.120 207.130 1162.260 254.590 ;
        RECT 1161.200 206.990 1162.260 207.130 ;
        RECT 1161.200 206.450 1161.340 206.990 ;
        RECT 1161.200 206.310 1161.800 206.450 ;
        RECT 1161.660 72.490 1161.800 206.310 ;
        RECT 1161.660 72.350 1162.260 72.490 ;
        RECT 1162.120 17.525 1162.260 72.350 ;
        RECT 50.230 17.155 50.510 17.525 ;
        RECT 1162.050 17.155 1162.330 17.525 ;
        RECT 50.300 2.400 50.440 17.155 ;
        RECT 50.090 -4.800 50.650 2.400 ;
      LAYER via2 ;
        RECT 1162.050 725.080 1162.330 725.360 ;
        RECT 1161.590 724.400 1161.870 724.680 ;
        RECT 50.230 17.200 50.510 17.480 ;
        RECT 1162.050 17.200 1162.330 17.480 ;
      LAYER met3 ;
        RECT 1162.025 725.370 1162.355 725.385 ;
        RECT 1161.350 725.070 1162.355 725.370 ;
        RECT 1161.350 724.705 1161.650 725.070 ;
        RECT 1162.025 725.055 1162.355 725.070 ;
        RECT 1161.350 724.390 1161.895 724.705 ;
        RECT 1161.565 724.375 1161.895 724.390 ;
        RECT 50.205 17.490 50.535 17.505 ;
        RECT 1162.025 17.490 1162.355 17.505 ;
        RECT 50.205 17.190 1162.355 17.490 ;
        RECT 50.205 17.175 50.535 17.190 ;
        RECT 1162.025 17.175 1162.355 17.190 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 72.290 1687.320 72.610 1687.380 ;
        RECT 1163.410 1687.320 1163.730 1687.380 ;
        RECT 72.290 1687.180 1163.730 1687.320 ;
        RECT 72.290 1687.120 72.610 1687.180 ;
        RECT 1163.410 1687.120 1163.730 1687.180 ;
        RECT 50.210 14.520 50.530 14.580 ;
        RECT 72.290 14.520 72.610 14.580 ;
        RECT 50.210 14.380 72.610 14.520 ;
        RECT 50.210 14.320 50.530 14.380 ;
        RECT 72.290 14.320 72.610 14.380 ;
      LAYER via ;
        RECT 72.320 1687.120 72.580 1687.380 ;
        RECT 1163.440 1687.120 1163.700 1687.380 ;
        RECT 50.240 14.320 50.500 14.580 ;
        RECT 72.320 14.320 72.580 14.580 ;
      LAYER met2 ;
        RECT 1163.430 1700.000 1163.710 1704.000 ;
        RECT 1163.500 1687.410 1163.640 1700.000 ;
        RECT 72.320 1687.090 72.580 1687.410 ;
        RECT 1163.440 1687.090 1163.700 1687.410 ;
        RECT 72.380 14.610 72.520 1687.090 ;
        RECT 50.240 14.290 50.500 14.610 ;
        RECT 72.320 14.290 72.580 14.610 ;
        RECT 50.300 2.400 50.440 14.290 ;
        RECT 50.090 -4.800 50.650 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 0.300 ;
=======
      LAYER li1 ;
        RECT 1197.525 18.445 1198.155 18.615 ;
        RECT 1186.945 17.255 1187.115 17.935 ;
        RECT 1186.945 17.085 1188.495 17.255 ;
        RECT 1196.605 16.915 1196.775 17.255 ;
        RECT 1197.525 16.915 1197.695 18.445 ;
        RECT 1196.605 16.745 1197.695 16.915 ;
      LAYER mcon ;
        RECT 1197.985 18.445 1198.155 18.615 ;
        RECT 1186.945 17.765 1187.115 17.935 ;
        RECT 1188.325 17.085 1188.495 17.255 ;
        RECT 1196.605 17.085 1196.775 17.255 ;
      LAYER met1 ;
        RECT 1214.470 1678.140 1214.790 1678.200 ;
        RECT 1216.770 1678.140 1217.090 1678.200 ;
        RECT 1214.470 1678.000 1217.090 1678.140 ;
        RECT 1214.470 1677.940 1214.790 1678.000 ;
        RECT 1216.770 1677.940 1217.090 1678.000 ;
        RECT 1197.925 18.600 1198.215 18.645 ;
        RECT 1214.470 18.600 1214.790 18.660 ;
        RECT 1197.925 18.460 1214.790 18.600 ;
        RECT 1197.925 18.415 1198.215 18.460 ;
        RECT 1214.470 18.400 1214.790 18.460 ;
        RECT 252.610 17.920 252.930 17.980 ;
        RECT 1186.885 17.920 1187.175 17.965 ;
        RECT 252.610 17.780 1187.175 17.920 ;
        RECT 252.610 17.720 252.930 17.780 ;
        RECT 1186.885 17.735 1187.175 17.780 ;
        RECT 1188.265 17.240 1188.555 17.285 ;
        RECT 1196.545 17.240 1196.835 17.285 ;
        RECT 1188.265 17.100 1196.835 17.240 ;
        RECT 1188.265 17.055 1188.555 17.100 ;
        RECT 1196.545 17.055 1196.835 17.100 ;
      LAYER via ;
        RECT 1214.500 1677.940 1214.760 1678.200 ;
        RECT 1216.800 1677.940 1217.060 1678.200 ;
        RECT 1214.500 18.400 1214.760 18.660 ;
        RECT 252.640 17.720 252.900 17.980 ;
      LAYER met2 ;
        RECT 1218.170 1700.410 1218.450 1704.000 ;
        RECT 1216.860 1700.270 1218.450 1700.410 ;
        RECT 1216.860 1678.230 1217.000 1700.270 ;
        RECT 1218.170 1700.000 1218.450 1700.270 ;
        RECT 1214.500 1677.910 1214.760 1678.230 ;
        RECT 1216.800 1677.910 1217.060 1678.230 ;
        RECT 1214.560 18.690 1214.700 1677.910 ;
        RECT 1214.500 18.370 1214.760 18.690 ;
        RECT 252.640 17.690 252.900 18.010 ;
        RECT 252.700 2.400 252.840 17.690 ;
        RECT 252.490 -4.800 253.050 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 0.300 ;
=======
      LAYER li1 ;
        RECT 1207.645 17.425 1207.815 34.595 ;
      LAYER mcon ;
        RECT 1207.645 34.425 1207.815 34.595 ;
      LAYER met1 ;
        RECT 1207.585 34.580 1207.875 34.625 ;
        RECT 1221.830 34.580 1222.150 34.640 ;
        RECT 1207.585 34.440 1222.150 34.580 ;
        RECT 1207.585 34.395 1207.875 34.440 ;
        RECT 1221.830 34.380 1222.150 34.440 ;
        RECT 270.090 18.260 270.410 18.320 ;
        RECT 1173.070 18.260 1173.390 18.320 ;
        RECT 270.090 18.120 1173.390 18.260 ;
        RECT 270.090 18.060 270.410 18.120 ;
        RECT 1173.070 18.060 1173.390 18.120 ;
        RECT 1202.970 17.580 1203.290 17.640 ;
        RECT 1207.585 17.580 1207.875 17.625 ;
        RECT 1202.970 17.440 1207.875 17.580 ;
        RECT 1202.970 17.380 1203.290 17.440 ;
        RECT 1207.585 17.395 1207.875 17.440 ;
      LAYER via ;
        RECT 1221.860 34.380 1222.120 34.640 ;
        RECT 270.120 18.060 270.380 18.320 ;
        RECT 1173.100 18.060 1173.360 18.320 ;
        RECT 1203.000 17.380 1203.260 17.640 ;
      LAYER met2 ;
        RECT 1222.770 1700.410 1223.050 1704.000 ;
        RECT 1221.920 1700.270 1223.050 1700.410 ;
        RECT 1221.920 34.670 1222.060 1700.270 ;
        RECT 1222.770 1700.000 1223.050 1700.270 ;
        RECT 1221.860 34.350 1222.120 34.670 ;
        RECT 270.120 18.030 270.380 18.350 ;
        RECT 1173.100 18.205 1173.360 18.350 ;
        RECT 270.180 2.400 270.320 18.030 ;
        RECT 1173.090 17.835 1173.370 18.205 ;
        RECT 1202.990 17.835 1203.270 18.205 ;
        RECT 1203.060 17.670 1203.200 17.835 ;
        RECT 1203.000 17.350 1203.260 17.670 ;
        RECT 269.970 -4.800 270.530 2.400 ;
      LAYER via2 ;
        RECT 1173.090 17.880 1173.370 18.160 ;
        RECT 1202.990 17.880 1203.270 18.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 1223.205 1380.210 1223.535 1380.225 ;
        RECT 1224.125 1380.210 1224.455 1380.225 ;
        RECT 1223.205 1379.910 1224.455 1380.210 ;
        RECT 1223.205 1379.895 1223.535 1379.910 ;
        RECT 1224.125 1379.895 1224.455 1379.910 ;
        RECT 1222.745 1283.650 1223.075 1283.665 ;
        RECT 1223.665 1283.650 1223.995 1283.665 ;
        RECT 1222.745 1283.350 1223.995 1283.650 ;
        RECT 1222.745 1283.335 1223.075 1283.350 ;
        RECT 1223.665 1283.335 1223.995 1283.350 ;
        RECT 1223.205 1152.410 1223.535 1152.425 ;
        RECT 1224.125 1152.410 1224.455 1152.425 ;
        RECT 1223.205 1152.110 1224.455 1152.410 ;
        RECT 1223.205 1152.095 1223.535 1152.110 ;
        RECT 1224.125 1152.095 1224.455 1152.110 ;
        RECT 1223.205 966.090 1223.535 966.105 ;
        RECT 1224.125 966.090 1224.455 966.105 ;
        RECT 1223.205 965.790 1224.455 966.090 ;
        RECT 1223.205 965.775 1223.535 965.790 ;
        RECT 1224.125 965.775 1224.455 965.790 ;
        RECT 1222.745 330.970 1223.075 330.985 ;
        RECT 1222.070 330.670 1223.075 330.970 ;
        RECT 1222.070 330.290 1222.370 330.670 ;
        RECT 1222.745 330.655 1223.075 330.670 ;
        RECT 1223.205 330.290 1223.535 330.305 ;
        RECT 1222.070 329.990 1223.535 330.290 ;
        RECT 1223.205 329.975 1223.535 329.990 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1173.065 18.170 1173.395 18.185 ;
        RECT 1202.965 18.170 1203.295 18.185 ;
        RECT 1173.065 17.870 1203.295 18.170 ;
        RECT 1173.065 17.855 1173.395 17.870 ;
        RECT 1202.965 17.855 1203.295 17.870 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 0.300 ;
=======
      LAYER met1 ;
        RECT 1223.670 1677.460 1223.990 1677.520 ;
        RECT 1226.430 1677.460 1226.750 1677.520 ;
        RECT 1223.670 1677.320 1226.750 1677.460 ;
        RECT 1223.670 1677.260 1223.990 1677.320 ;
        RECT 1226.430 1677.260 1226.750 1677.320 ;
        RECT 1223.670 18.940 1223.990 19.000 ;
        RECT 1197.540 18.800 1223.990 18.940 ;
        RECT 288.030 18.600 288.350 18.660 ;
        RECT 1197.540 18.600 1197.680 18.800 ;
        RECT 1223.670 18.740 1223.990 18.800 ;
        RECT 288.030 18.460 1197.680 18.600 ;
        RECT 288.030 18.400 288.350 18.460 ;
      LAYER via ;
        RECT 1223.700 1677.260 1223.960 1677.520 ;
        RECT 1226.460 1677.260 1226.720 1677.520 ;
        RECT 288.060 18.400 288.320 18.660 ;
        RECT 1223.700 18.740 1223.960 19.000 ;
      LAYER met2 ;
        RECT 1227.830 1700.410 1228.110 1704.000 ;
        RECT 1226.520 1700.270 1228.110 1700.410 ;
        RECT 1226.520 1677.550 1226.660 1700.270 ;
        RECT 1227.830 1700.000 1228.110 1700.270 ;
        RECT 1223.700 1677.230 1223.960 1677.550 ;
        RECT 1226.460 1677.230 1226.720 1677.550 ;
        RECT 1223.760 19.030 1223.900 1677.230 ;
        RECT 1223.700 18.710 1223.960 19.030 ;
        RECT 288.060 18.370 288.320 18.690 ;
        RECT 288.120 2.400 288.260 18.370 ;
        RECT 287.910 -4.800 288.470 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 0.300 ;
=======
      LAYER li1 ;
        RECT 1178.665 1687.505 1178.835 1689.035 ;
      LAYER mcon ;
        RECT 1178.665 1688.865 1178.835 1689.035 ;
      LAYER met1 ;
        RECT 310.110 1689.020 310.430 1689.080 ;
        RECT 1178.605 1689.020 1178.895 1689.065 ;
        RECT 310.110 1688.880 1178.895 1689.020 ;
        RECT 310.110 1688.820 310.430 1688.880 ;
        RECT 1178.605 1688.835 1178.895 1688.880 ;
        RECT 1178.605 1687.660 1178.895 1687.705 ;
        RECT 1232.410 1687.660 1232.730 1687.720 ;
        RECT 1178.605 1687.520 1232.730 1687.660 ;
        RECT 1178.605 1687.475 1178.895 1687.520 ;
        RECT 1232.410 1687.460 1232.730 1687.520 ;
        RECT 305.970 16.900 306.290 16.960 ;
        RECT 310.110 16.900 310.430 16.960 ;
        RECT 305.970 16.760 310.430 16.900 ;
        RECT 305.970 16.700 306.290 16.760 ;
        RECT 310.110 16.700 310.430 16.760 ;
      LAYER via ;
        RECT 310.140 1688.820 310.400 1689.080 ;
        RECT 1232.440 1687.460 1232.700 1687.720 ;
        RECT 306.000 16.700 306.260 16.960 ;
        RECT 310.140 16.700 310.400 16.960 ;
      LAYER met2 ;
        RECT 1232.430 1700.000 1232.710 1704.000 ;
        RECT 310.140 1688.790 310.400 1689.110 ;
        RECT 310.200 16.990 310.340 1688.790 ;
        RECT 1232.500 1687.750 1232.640 1700.000 ;
        RECT 1232.440 1687.430 1232.700 1687.750 ;
        RECT 306.000 16.670 306.260 16.990 ;
        RECT 310.140 16.670 310.400 16.990 ;
        RECT 306.060 2.400 306.200 16.670 ;
=======
      LAYER met1 ;
        RECT 1228.270 1678.140 1228.590 1678.200 ;
        RECT 1231.490 1678.140 1231.810 1678.200 ;
        RECT 1228.270 1678.000 1231.810 1678.140 ;
        RECT 1228.270 1677.940 1228.590 1678.000 ;
        RECT 1231.490 1677.940 1231.810 1678.000 ;
        RECT 1228.270 19.280 1228.590 19.340 ;
        RECT 1197.080 19.140 1228.590 19.280 ;
        RECT 305.970 18.940 306.290 19.000 ;
        RECT 1197.080 18.940 1197.220 19.140 ;
        RECT 1228.270 19.080 1228.590 19.140 ;
        RECT 305.970 18.800 1197.220 18.940 ;
        RECT 305.970 18.740 306.290 18.800 ;
      LAYER via ;
        RECT 1228.300 1677.940 1228.560 1678.200 ;
        RECT 1231.520 1677.940 1231.780 1678.200 ;
        RECT 306.000 18.740 306.260 19.000 ;
        RECT 1228.300 19.080 1228.560 19.340 ;
      LAYER met2 ;
        RECT 1232.430 1700.410 1232.710 1704.000 ;
        RECT 1231.580 1700.270 1232.710 1700.410 ;
        RECT 1231.580 1678.230 1231.720 1700.270 ;
        RECT 1232.430 1700.000 1232.710 1700.270 ;
        RECT 1228.300 1677.910 1228.560 1678.230 ;
        RECT 1231.520 1677.910 1231.780 1678.230 ;
        RECT 1228.360 19.370 1228.500 1677.910 ;
        RECT 1228.300 19.050 1228.560 19.370 ;
        RECT 306.000 18.710 306.260 19.030 ;
        RECT 306.060 2.400 306.200 18.710 ;
>>>>>>> re-updated local openlane
        RECT 305.850 -4.800 306.410 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 0.300 ;
=======
      LAYER li1 ;
        RECT 1196.605 17.765 1196.775 19.295 ;
        RECT 1215.005 17.765 1215.175 19.975 ;
      LAYER mcon ;
        RECT 1215.005 19.805 1215.175 19.975 ;
        RECT 1196.605 19.125 1196.775 19.295 ;
      LAYER met1 ;
        RECT 1235.170 1695.480 1235.490 1695.540 ;
        RECT 1237.470 1695.480 1237.790 1695.540 ;
        RECT 1235.170 1695.340 1237.790 1695.480 ;
        RECT 1235.170 1695.280 1235.490 1695.340 ;
        RECT 1237.470 1695.280 1237.790 1695.340 ;
        RECT 1214.945 19.960 1215.235 20.005 ;
        RECT 1235.170 19.960 1235.490 20.020 ;
        RECT 1214.945 19.820 1235.490 19.960 ;
        RECT 1214.945 19.775 1215.235 19.820 ;
        RECT 1235.170 19.760 1235.490 19.820 ;
        RECT 323.450 19.280 323.770 19.340 ;
        RECT 1196.545 19.280 1196.835 19.325 ;
        RECT 323.450 19.140 1196.835 19.280 ;
        RECT 323.450 19.080 323.770 19.140 ;
        RECT 1196.545 19.095 1196.835 19.140 ;
        RECT 1196.545 17.920 1196.835 17.965 ;
        RECT 1214.945 17.920 1215.235 17.965 ;
        RECT 1196.545 17.780 1215.235 17.920 ;
        RECT 1196.545 17.735 1196.835 17.780 ;
        RECT 1214.945 17.735 1215.235 17.780 ;
      LAYER via ;
        RECT 1235.200 1695.280 1235.460 1695.540 ;
        RECT 1237.500 1695.280 1237.760 1695.540 ;
        RECT 1235.200 19.760 1235.460 20.020 ;
        RECT 323.480 19.080 323.740 19.340 ;
      LAYER met2 ;
        RECT 1237.490 1700.000 1237.770 1704.000 ;
        RECT 1237.560 1695.570 1237.700 1700.000 ;
        RECT 1235.200 1695.250 1235.460 1695.570 ;
        RECT 1237.500 1695.250 1237.760 1695.570 ;
        RECT 1235.260 20.050 1235.400 1695.250 ;
        RECT 1235.200 19.730 1235.460 20.050 ;
        RECT 323.480 19.050 323.740 19.370 ;
        RECT 323.540 9.930 323.680 19.050 ;
        RECT 323.540 9.790 324.140 9.930 ;
        RECT 324.000 2.400 324.140 9.790 ;
        RECT 323.790 -4.800 324.350 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 0.300 ;
=======
      LAYER met1 ;
        RECT 341.390 19.620 341.710 19.680 ;
        RECT 1242.530 19.620 1242.850 19.680 ;
        RECT 341.390 19.480 1242.850 19.620 ;
        RECT 341.390 19.420 341.710 19.480 ;
        RECT 1242.530 19.420 1242.850 19.480 ;
      LAYER via ;
        RECT 341.420 19.420 341.680 19.680 ;
        RECT 1242.560 19.420 1242.820 19.680 ;
      LAYER met2 ;
        RECT 1242.090 1700.410 1242.370 1704.000 ;
        RECT 1242.090 1700.270 1242.760 1700.410 ;
        RECT 1242.090 1700.000 1242.370 1700.270 ;
        RECT 1242.620 19.710 1242.760 1700.270 ;
        RECT 341.420 19.390 341.680 19.710 ;
        RECT 1242.560 19.390 1242.820 19.710 ;
        RECT 341.480 2.400 341.620 19.390 ;
        RECT 341.270 -4.800 341.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 0.300 ;
=======
      LAYER met1 ;
        RECT 365.310 1689.700 365.630 1689.760 ;
        RECT 1246.670 1689.700 1246.990 1689.760 ;
        RECT 365.310 1689.560 1246.990 1689.700 ;
        RECT 365.310 1689.500 365.630 1689.560 ;
        RECT 1246.670 1689.500 1246.990 1689.560 ;
        RECT 359.330 16.900 359.650 16.960 ;
        RECT 365.310 16.900 365.630 16.960 ;
        RECT 359.330 16.760 365.630 16.900 ;
        RECT 359.330 16.700 359.650 16.760 ;
        RECT 365.310 16.700 365.630 16.760 ;
      LAYER via ;
        RECT 365.340 1689.500 365.600 1689.760 ;
        RECT 1246.700 1689.500 1246.960 1689.760 ;
        RECT 359.360 16.700 359.620 16.960 ;
        RECT 365.340 16.700 365.600 16.960 ;
      LAYER met2 ;
        RECT 1246.690 1700.000 1246.970 1704.000 ;
        RECT 1246.760 1689.790 1246.900 1700.000 ;
        RECT 365.340 1689.470 365.600 1689.790 ;
        RECT 1246.700 1689.470 1246.960 1689.790 ;
        RECT 365.400 16.990 365.540 1689.470 ;
        RECT 359.360 16.670 359.620 16.990 ;
        RECT 365.340 16.670 365.600 16.990 ;
        RECT 359.420 2.400 359.560 16.670 ;
        RECT 359.210 -4.800 359.770 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1243.985 1580.065 1244.155 1669.655 ;
        RECT 1244.445 1049.325 1244.615 1097.095 ;
        RECT 1244.445 1024.165 1244.615 1048.815 ;
        RECT 1243.985 848.725 1244.155 896.835 ;
        RECT 1243.985 807.245 1244.155 832.915 ;
        RECT 1243.985 730.745 1244.155 738.735 ;
        RECT 1243.985 379.525 1244.155 427.635 ;
      LAYER mcon ;
        RECT 1243.985 1669.485 1244.155 1669.655 ;
        RECT 1244.445 1096.925 1244.615 1097.095 ;
        RECT 1244.445 1048.645 1244.615 1048.815 ;
        RECT 1243.985 896.665 1244.155 896.835 ;
        RECT 1243.985 832.745 1244.155 832.915 ;
        RECT 1243.985 738.565 1244.155 738.735 ;
        RECT 1243.985 427.465 1244.155 427.635 ;
      LAYER met1 ;
        RECT 1243.925 1669.640 1244.215 1669.685 ;
        RECT 1244.370 1669.640 1244.690 1669.700 ;
        RECT 1243.925 1669.500 1244.690 1669.640 ;
        RECT 1243.925 1669.455 1244.215 1669.500 ;
        RECT 1244.370 1669.440 1244.690 1669.500 ;
        RECT 1243.910 1580.220 1244.230 1580.280 ;
        RECT 1243.715 1580.080 1244.230 1580.220 ;
        RECT 1243.910 1580.020 1244.230 1580.080 ;
        RECT 1243.910 1490.800 1244.230 1490.860 ;
        RECT 1244.830 1490.800 1245.150 1490.860 ;
        RECT 1243.910 1490.660 1245.150 1490.800 ;
        RECT 1243.910 1490.600 1244.230 1490.660 ;
        RECT 1244.830 1490.600 1245.150 1490.660 ;
        RECT 1245.290 1435.380 1245.610 1435.440 ;
        RECT 1246.210 1435.380 1246.530 1435.440 ;
        RECT 1245.290 1435.240 1246.530 1435.380 ;
        RECT 1245.290 1435.180 1245.610 1435.240 ;
        RECT 1246.210 1435.180 1246.530 1435.240 ;
        RECT 1243.910 1269.600 1244.230 1269.860 ;
        RECT 1244.000 1269.120 1244.140 1269.600 ;
        RECT 1244.370 1269.120 1244.690 1269.180 ;
        RECT 1244.000 1268.980 1244.690 1269.120 ;
        RECT 1244.370 1268.920 1244.690 1268.980 ;
        RECT 1244.370 1207.920 1244.690 1207.980 ;
        RECT 1244.000 1207.780 1244.690 1207.920 ;
        RECT 1244.000 1207.640 1244.140 1207.780 ;
        RECT 1244.370 1207.720 1244.690 1207.780 ;
        RECT 1243.910 1207.380 1244.230 1207.640 ;
        RECT 1243.910 1173.040 1244.230 1173.300 ;
        RECT 1244.000 1172.560 1244.140 1173.040 ;
        RECT 1244.370 1172.560 1244.690 1172.620 ;
        RECT 1244.000 1172.420 1244.690 1172.560 ;
        RECT 1244.370 1172.360 1244.690 1172.420 ;
        RECT 1244.370 1097.080 1244.690 1097.140 ;
        RECT 1244.175 1096.940 1244.690 1097.080 ;
        RECT 1244.370 1096.880 1244.690 1096.940 ;
        RECT 1244.370 1049.480 1244.690 1049.540 ;
        RECT 1244.175 1049.340 1244.690 1049.480 ;
        RECT 1244.370 1049.280 1244.690 1049.340 ;
        RECT 1244.370 1048.800 1244.690 1048.860 ;
        RECT 1244.175 1048.660 1244.690 1048.800 ;
        RECT 1244.370 1048.600 1244.690 1048.660 ;
        RECT 1244.370 1024.320 1244.690 1024.380 ;
        RECT 1244.175 1024.180 1244.690 1024.320 ;
        RECT 1244.370 1024.120 1244.690 1024.180 ;
        RECT 1244.370 1000.520 1244.690 1000.580 ;
        RECT 1245.290 1000.520 1245.610 1000.580 ;
        RECT 1244.370 1000.380 1245.610 1000.520 ;
        RECT 1244.370 1000.320 1244.690 1000.380 ;
        RECT 1245.290 1000.320 1245.610 1000.380 ;
        RECT 1243.910 934.900 1244.230 934.960 ;
        RECT 1244.830 934.900 1245.150 934.960 ;
        RECT 1243.910 934.760 1245.150 934.900 ;
        RECT 1243.910 934.700 1244.230 934.760 ;
        RECT 1244.830 934.700 1245.150 934.760 ;
        RECT 1243.910 896.820 1244.230 896.880 ;
        RECT 1243.715 896.680 1244.230 896.820 ;
        RECT 1243.910 896.620 1244.230 896.680 ;
        RECT 1243.925 848.880 1244.215 848.925 ;
        RECT 1244.370 848.880 1244.690 848.940 ;
        RECT 1243.925 848.740 1244.690 848.880 ;
        RECT 1243.925 848.695 1244.215 848.740 ;
        RECT 1244.370 848.680 1244.690 848.740 ;
        RECT 1243.925 832.900 1244.215 832.945 ;
        RECT 1244.370 832.900 1244.690 832.960 ;
        RECT 1243.925 832.760 1244.690 832.900 ;
        RECT 1243.925 832.715 1244.215 832.760 ;
        RECT 1244.370 832.700 1244.690 832.760 ;
        RECT 1243.910 807.400 1244.230 807.460 ;
        RECT 1243.715 807.260 1244.230 807.400 ;
        RECT 1243.910 807.200 1244.230 807.260 ;
        RECT 1243.925 738.720 1244.215 738.765 ;
        RECT 1244.370 738.720 1244.690 738.780 ;
        RECT 1243.925 738.580 1244.690 738.720 ;
        RECT 1243.925 738.535 1244.215 738.580 ;
        RECT 1244.370 738.520 1244.690 738.580 ;
        RECT 1243.910 730.900 1244.230 730.960 ;
        RECT 1243.715 730.760 1244.230 730.900 ;
        RECT 1243.910 730.700 1244.230 730.760 ;
        RECT 1244.370 545.600 1244.690 545.660 ;
        RECT 1244.000 545.460 1244.690 545.600 ;
        RECT 1244.000 544.980 1244.140 545.460 ;
        RECT 1244.370 545.400 1244.690 545.460 ;
        RECT 1243.910 544.720 1244.230 544.980 ;
        RECT 1243.910 496.780 1244.230 497.040 ;
        RECT 1244.000 496.640 1244.140 496.780 ;
        RECT 1244.370 496.640 1244.690 496.700 ;
        RECT 1244.000 496.500 1244.690 496.640 ;
        RECT 1244.370 496.440 1244.690 496.500 ;
        RECT 1244.370 448.500 1244.690 448.760 ;
        RECT 1244.460 448.360 1244.600 448.500 ;
        RECT 1244.830 448.360 1245.150 448.420 ;
        RECT 1244.460 448.220 1245.150 448.360 ;
        RECT 1244.830 448.160 1245.150 448.220 ;
        RECT 1243.925 427.620 1244.215 427.665 ;
        RECT 1244.830 427.620 1245.150 427.680 ;
        RECT 1243.925 427.480 1245.150 427.620 ;
        RECT 1243.925 427.435 1244.215 427.480 ;
        RECT 1244.830 427.420 1245.150 427.480 ;
        RECT 1243.910 379.680 1244.230 379.740 ;
        RECT 1243.715 379.540 1244.230 379.680 ;
        RECT 1243.910 379.480 1244.230 379.540 ;
        RECT 1244.370 283.120 1244.690 283.180 ;
        RECT 1244.830 283.120 1245.150 283.180 ;
        RECT 1244.370 282.980 1245.150 283.120 ;
        RECT 1244.370 282.920 1244.690 282.980 ;
        RECT 1244.830 282.920 1245.150 282.980 ;
        RECT 1244.370 235.180 1244.690 235.240 ;
        RECT 1244.000 235.040 1244.690 235.180 ;
        RECT 1244.000 234.900 1244.140 235.040 ;
        RECT 1244.370 234.980 1244.690 235.040 ;
        RECT 1243.910 234.640 1244.230 234.900 ;
        RECT 1243.910 137.940 1244.230 138.000 ;
        RECT 1244.370 137.940 1244.690 138.000 ;
        RECT 1243.910 137.800 1244.690 137.940 ;
        RECT 1243.910 137.740 1244.230 137.800 ;
        RECT 1244.370 137.740 1244.690 137.800 ;
        RECT 1244.370 20.300 1244.690 20.360 ;
        RECT 1214.560 20.160 1244.690 20.300 ;
        RECT 359.330 19.960 359.650 20.020 ;
        RECT 1214.560 19.960 1214.700 20.160 ;
        RECT 1244.370 20.100 1244.690 20.160 ;
        RECT 359.330 19.820 1214.700 19.960 ;
        RECT 359.330 19.760 359.650 19.820 ;
      LAYER via ;
        RECT 1244.400 1669.440 1244.660 1669.700 ;
        RECT 1243.940 1580.020 1244.200 1580.280 ;
        RECT 1243.940 1490.600 1244.200 1490.860 ;
        RECT 1244.860 1490.600 1245.120 1490.860 ;
        RECT 1245.320 1435.180 1245.580 1435.440 ;
        RECT 1246.240 1435.180 1246.500 1435.440 ;
        RECT 1243.940 1269.600 1244.200 1269.860 ;
        RECT 1244.400 1268.920 1244.660 1269.180 ;
        RECT 1244.400 1207.720 1244.660 1207.980 ;
        RECT 1243.940 1207.380 1244.200 1207.640 ;
        RECT 1243.940 1173.040 1244.200 1173.300 ;
        RECT 1244.400 1172.360 1244.660 1172.620 ;
        RECT 1244.400 1096.880 1244.660 1097.140 ;
        RECT 1244.400 1049.280 1244.660 1049.540 ;
        RECT 1244.400 1048.600 1244.660 1048.860 ;
        RECT 1244.400 1024.120 1244.660 1024.380 ;
        RECT 1244.400 1000.320 1244.660 1000.580 ;
        RECT 1245.320 1000.320 1245.580 1000.580 ;
        RECT 1243.940 934.700 1244.200 934.960 ;
        RECT 1244.860 934.700 1245.120 934.960 ;
        RECT 1243.940 896.620 1244.200 896.880 ;
        RECT 1244.400 848.680 1244.660 848.940 ;
        RECT 1244.400 832.700 1244.660 832.960 ;
        RECT 1243.940 807.200 1244.200 807.460 ;
        RECT 1244.400 738.520 1244.660 738.780 ;
        RECT 1243.940 730.700 1244.200 730.960 ;
        RECT 1244.400 545.400 1244.660 545.660 ;
        RECT 1243.940 544.720 1244.200 544.980 ;
        RECT 1243.940 496.780 1244.200 497.040 ;
        RECT 1244.400 496.440 1244.660 496.700 ;
        RECT 1244.400 448.500 1244.660 448.760 ;
        RECT 1244.860 448.160 1245.120 448.420 ;
        RECT 1244.860 427.420 1245.120 427.680 ;
        RECT 1243.940 379.480 1244.200 379.740 ;
        RECT 1244.400 282.920 1244.660 283.180 ;
        RECT 1244.860 282.920 1245.120 283.180 ;
        RECT 1244.400 234.980 1244.660 235.240 ;
        RECT 1243.940 234.640 1244.200 234.900 ;
        RECT 1243.940 137.740 1244.200 138.000 ;
        RECT 1244.400 137.740 1244.660 138.000 ;
        RECT 359.360 19.760 359.620 20.020 ;
        RECT 1244.400 20.100 1244.660 20.360 ;
      LAYER met2 ;
        RECT 1247.150 1700.410 1247.430 1704.000 ;
        RECT 1245.840 1700.270 1247.430 1700.410 ;
        RECT 1245.840 1676.725 1245.980 1700.270 ;
        RECT 1247.150 1700.000 1247.430 1700.270 ;
        RECT 1244.390 1676.355 1244.670 1676.725 ;
        RECT 1245.770 1676.355 1246.050 1676.725 ;
        RECT 1244.460 1669.730 1244.600 1676.355 ;
        RECT 1244.400 1669.410 1244.660 1669.730 ;
        RECT 1243.940 1579.990 1244.200 1580.310 ;
        RECT 1244.000 1490.890 1244.140 1579.990 ;
        RECT 1243.940 1490.570 1244.200 1490.890 ;
        RECT 1244.860 1490.570 1245.120 1490.890 ;
        RECT 1244.920 1483.605 1245.060 1490.570 ;
        RECT 1244.850 1483.235 1245.130 1483.605 ;
        RECT 1246.230 1483.235 1246.510 1483.605 ;
        RECT 1246.300 1435.470 1246.440 1483.235 ;
        RECT 1245.320 1435.150 1245.580 1435.470 ;
        RECT 1246.240 1435.150 1246.500 1435.470 ;
        RECT 1245.380 1418.210 1245.520 1435.150 ;
        RECT 1244.000 1418.070 1245.520 1418.210 ;
        RECT 1244.000 1269.890 1244.140 1418.070 ;
        RECT 1243.940 1269.570 1244.200 1269.890 ;
        RECT 1244.400 1268.890 1244.660 1269.210 ;
        RECT 1244.460 1208.010 1244.600 1268.890 ;
        RECT 1244.400 1207.690 1244.660 1208.010 ;
        RECT 1243.940 1207.350 1244.200 1207.670 ;
        RECT 1244.000 1173.330 1244.140 1207.350 ;
        RECT 1243.940 1173.010 1244.200 1173.330 ;
        RECT 1244.400 1172.330 1244.660 1172.650 ;
        RECT 1244.460 1097.170 1244.600 1172.330 ;
        RECT 1244.400 1096.850 1244.660 1097.170 ;
        RECT 1244.400 1049.250 1244.660 1049.570 ;
        RECT 1244.460 1048.890 1244.600 1049.250 ;
        RECT 1244.400 1048.570 1244.660 1048.890 ;
        RECT 1244.400 1024.090 1244.660 1024.410 ;
        RECT 1244.460 1000.610 1244.600 1024.090 ;
        RECT 1244.400 1000.290 1244.660 1000.610 ;
        RECT 1245.320 1000.290 1245.580 1000.610 ;
        RECT 1245.380 959.040 1245.520 1000.290 ;
        RECT 1244.920 958.900 1245.520 959.040 ;
        RECT 1244.920 934.990 1245.060 958.900 ;
        RECT 1243.940 934.670 1244.200 934.990 ;
        RECT 1244.860 934.670 1245.120 934.990 ;
        RECT 1244.000 896.910 1244.140 934.670 ;
        RECT 1243.940 896.590 1244.200 896.910 ;
        RECT 1244.400 848.650 1244.660 848.970 ;
        RECT 1244.460 832.990 1244.600 848.650 ;
        RECT 1244.400 832.670 1244.660 832.990 ;
        RECT 1243.940 807.170 1244.200 807.490 ;
        RECT 1244.000 783.090 1244.140 807.170 ;
        RECT 1244.000 782.950 1244.600 783.090 ;
        RECT 1244.460 738.810 1244.600 782.950 ;
        RECT 1244.400 738.490 1244.660 738.810 ;
        RECT 1243.940 730.670 1244.200 730.990 ;
        RECT 1244.000 686.530 1244.140 730.670 ;
        RECT 1244.000 686.390 1245.060 686.530 ;
        RECT 1244.920 596.090 1245.060 686.390 ;
        RECT 1244.460 595.950 1245.060 596.090 ;
        RECT 1244.460 545.690 1244.600 595.950 ;
        RECT 1244.400 545.370 1244.660 545.690 ;
        RECT 1243.940 544.690 1244.200 545.010 ;
        RECT 1244.000 497.070 1244.140 544.690 ;
        RECT 1243.940 496.750 1244.200 497.070 ;
        RECT 1244.400 496.410 1244.660 496.730 ;
        RECT 1244.460 448.790 1244.600 496.410 ;
        RECT 1244.400 448.470 1244.660 448.790 ;
        RECT 1244.860 448.130 1245.120 448.450 ;
        RECT 1244.920 427.710 1245.060 448.130 ;
        RECT 1244.860 427.390 1245.120 427.710 ;
        RECT 1243.940 379.450 1244.200 379.770 ;
        RECT 1244.000 331.005 1244.140 379.450 ;
        RECT 1243.930 330.635 1244.210 331.005 ;
        RECT 1244.850 329.955 1245.130 330.325 ;
        RECT 1244.920 283.210 1245.060 329.955 ;
        RECT 1244.400 282.890 1244.660 283.210 ;
        RECT 1244.860 282.890 1245.120 283.210 ;
        RECT 1244.460 235.270 1244.600 282.890 ;
        RECT 1244.400 234.950 1244.660 235.270 ;
        RECT 1243.940 234.610 1244.200 234.930 ;
        RECT 1244.000 186.050 1244.140 234.610 ;
        RECT 1244.000 185.910 1244.600 186.050 ;
        RECT 1244.460 139.245 1244.600 185.910 ;
        RECT 1244.390 138.875 1244.670 139.245 ;
        RECT 1243.930 138.195 1244.210 138.565 ;
        RECT 1244.000 138.030 1244.140 138.195 ;
        RECT 1243.940 137.710 1244.200 138.030 ;
        RECT 1244.400 137.710 1244.660 138.030 ;
        RECT 1244.460 20.390 1244.600 137.710 ;
        RECT 1244.400 20.070 1244.660 20.390 ;
        RECT 359.360 19.730 359.620 20.050 ;
        RECT 359.420 2.400 359.560 19.730 ;
        RECT 359.210 -4.800 359.770 2.400 ;
      LAYER via2 ;
        RECT 1244.390 1676.400 1244.670 1676.680 ;
        RECT 1245.770 1676.400 1246.050 1676.680 ;
        RECT 1244.850 1483.280 1245.130 1483.560 ;
        RECT 1246.230 1483.280 1246.510 1483.560 ;
        RECT 1243.930 330.680 1244.210 330.960 ;
        RECT 1244.850 330.000 1245.130 330.280 ;
        RECT 1244.390 138.920 1244.670 139.200 ;
        RECT 1243.930 138.240 1244.210 138.520 ;
      LAYER met3 ;
        RECT 1244.365 1676.690 1244.695 1676.705 ;
        RECT 1245.745 1676.690 1246.075 1676.705 ;
        RECT 1244.365 1676.390 1246.075 1676.690 ;
        RECT 1244.365 1676.375 1244.695 1676.390 ;
        RECT 1245.745 1676.375 1246.075 1676.390 ;
        RECT 1244.825 1483.570 1245.155 1483.585 ;
        RECT 1246.205 1483.570 1246.535 1483.585 ;
        RECT 1244.825 1483.270 1246.535 1483.570 ;
        RECT 1244.825 1483.255 1245.155 1483.270 ;
        RECT 1246.205 1483.255 1246.535 1483.270 ;
        RECT 1243.905 330.970 1244.235 330.985 ;
        RECT 1243.230 330.670 1244.235 330.970 ;
        RECT 1243.230 330.290 1243.530 330.670 ;
        RECT 1243.905 330.655 1244.235 330.670 ;
        RECT 1244.825 330.290 1245.155 330.305 ;
        RECT 1243.230 329.990 1245.155 330.290 ;
        RECT 1244.825 329.975 1245.155 329.990 ;
        RECT 1244.365 139.210 1244.695 139.225 ;
        RECT 1243.230 138.910 1244.695 139.210 ;
        RECT 1243.230 138.530 1243.530 138.910 ;
        RECT 1244.365 138.895 1244.695 138.910 ;
        RECT 1243.905 138.530 1244.235 138.545 ;
        RECT 1243.230 138.230 1244.235 138.530 ;
        RECT 1243.905 138.215 1244.235 138.230 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 0.300 ;
=======
      LAYER li1 ;
        RECT 1197.065 17.085 1197.235 20.315 ;
      LAYER mcon ;
        RECT 1197.065 20.145 1197.235 20.315 ;
      LAYER met1 ;
        RECT 1248.970 1661.480 1249.290 1661.540 ;
        RECT 1250.810 1661.480 1251.130 1661.540 ;
        RECT 1248.970 1661.340 1251.130 1661.480 ;
        RECT 1248.970 1661.280 1249.290 1661.340 ;
        RECT 1250.810 1661.280 1251.130 1661.340 ;
        RECT 377.270 20.300 377.590 20.360 ;
        RECT 1197.005 20.300 1197.295 20.345 ;
        RECT 377.270 20.160 1197.295 20.300 ;
        RECT 377.270 20.100 377.590 20.160 ;
        RECT 1197.005 20.115 1197.295 20.160 ;
        RECT 1197.005 17.240 1197.295 17.285 ;
        RECT 1248.970 17.240 1249.290 17.300 ;
        RECT 1197.005 17.100 1249.290 17.240 ;
        RECT 1197.005 17.055 1197.295 17.100 ;
        RECT 1248.970 17.040 1249.290 17.100 ;
      LAYER via ;
        RECT 1249.000 1661.280 1249.260 1661.540 ;
        RECT 1250.840 1661.280 1251.100 1661.540 ;
        RECT 377.300 20.100 377.560 20.360 ;
        RECT 1249.000 17.040 1249.260 17.300 ;
      LAYER met2 ;
        RECT 1251.750 1700.410 1252.030 1704.000 ;
        RECT 1250.900 1700.270 1252.030 1700.410 ;
        RECT 1250.900 1661.570 1251.040 1700.270 ;
        RECT 1251.750 1700.000 1252.030 1700.270 ;
        RECT 1249.000 1661.250 1249.260 1661.570 ;
        RECT 1250.840 1661.250 1251.100 1661.570 ;
        RECT 377.300 20.070 377.560 20.390 ;
        RECT 377.360 2.400 377.500 20.070 ;
        RECT 1249.060 17.330 1249.200 1661.250 ;
        RECT 1249.000 17.010 1249.260 17.330 ;
        RECT 377.150 -4.800 377.710 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 0.300 ;
=======
      LAYER met1 ;
        RECT 395.210 20.640 395.530 20.700 ;
        RECT 1255.870 20.640 1256.190 20.700 ;
        RECT 395.210 20.500 1256.190 20.640 ;
        RECT 395.210 20.440 395.530 20.500 ;
        RECT 1255.870 20.440 1256.190 20.500 ;
      LAYER via ;
        RECT 395.240 20.440 395.500 20.700 ;
        RECT 1255.900 20.440 1256.160 20.700 ;
      LAYER met2 ;
        RECT 1256.810 1700.410 1257.090 1704.000 ;
        RECT 1255.960 1700.270 1257.090 1700.410 ;
        RECT 1255.960 20.730 1256.100 1700.270 ;
        RECT 1256.810 1700.000 1257.090 1700.270 ;
        RECT 395.240 20.410 395.500 20.730 ;
        RECT 1255.900 20.410 1256.160 20.730 ;
        RECT 395.300 2.400 395.440 20.410 ;
        RECT 395.090 -4.800 395.650 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 0.300 ;
=======
      LAYER met1 ;
        RECT 1256.330 1672.360 1256.650 1672.420 ;
        RECT 1260.470 1672.360 1260.790 1672.420 ;
        RECT 1256.330 1672.220 1260.790 1672.360 ;
        RECT 1256.330 1672.160 1256.650 1672.220 ;
        RECT 1260.470 1672.160 1260.790 1672.220 ;
        RECT 1256.330 16.900 1256.650 16.960 ;
        RECT 414.160 16.760 1256.650 16.900 ;
        RECT 413.150 16.220 413.470 16.280 ;
        RECT 414.160 16.220 414.300 16.760 ;
        RECT 1256.330 16.700 1256.650 16.760 ;
        RECT 413.150 16.080 414.300 16.220 ;
        RECT 413.150 16.020 413.470 16.080 ;
      LAYER via ;
        RECT 1256.360 1672.160 1256.620 1672.420 ;
        RECT 1260.500 1672.160 1260.760 1672.420 ;
        RECT 413.180 16.020 413.440 16.280 ;
        RECT 1256.360 16.700 1256.620 16.960 ;
      LAYER met2 ;
        RECT 1261.410 1700.410 1261.690 1704.000 ;
        RECT 1260.560 1700.270 1261.690 1700.410 ;
        RECT 1260.560 1672.450 1260.700 1700.270 ;
        RECT 1261.410 1700.000 1261.690 1700.270 ;
        RECT 1256.360 1672.130 1256.620 1672.450 ;
        RECT 1260.500 1672.130 1260.760 1672.450 ;
        RECT 1256.420 16.990 1256.560 1672.130 ;
        RECT 1256.360 16.670 1256.620 16.990 ;
        RECT 413.180 15.990 413.440 16.310 ;
        RECT 413.240 2.400 413.380 15.990 ;
        RECT 413.030 -4.800 413.590 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 74.010 -4.800 74.570 0.300 ;
=======
        RECT 1169.410 1700.410 1169.690 1704.000 ;
        RECT 1169.020 1700.270 1169.690 1700.410 ;
        RECT 1169.020 18.885 1169.160 1700.270 ;
        RECT 1169.410 1700.000 1169.690 1700.270 ;
        RECT 74.150 18.515 74.430 18.885 ;
        RECT 1168.950 18.515 1169.230 18.885 ;
        RECT 74.220 2.400 74.360 18.515 ;
=======
      LAYER li1 ;
        RECT 1168.545 1635.485 1168.715 1683.595 ;
        RECT 1168.545 1538.925 1168.715 1587.035 ;
        RECT 1168.545 1442.025 1168.715 1490.475 ;
        RECT 1168.545 572.645 1168.715 620.755 ;
        RECT 1168.545 476.085 1168.715 524.195 ;
        RECT 1168.545 379.525 1168.715 427.635 ;
        RECT 1168.545 282.965 1168.715 331.075 ;
        RECT 1167.625 186.405 1167.795 234.515 ;
        RECT 1167.625 48.365 1167.795 137.955 ;
      LAYER mcon ;
        RECT 1168.545 1683.425 1168.715 1683.595 ;
        RECT 1168.545 1586.865 1168.715 1587.035 ;
        RECT 1168.545 1490.305 1168.715 1490.475 ;
        RECT 1168.545 620.585 1168.715 620.755 ;
        RECT 1168.545 524.025 1168.715 524.195 ;
        RECT 1168.545 427.465 1168.715 427.635 ;
        RECT 1168.545 330.905 1168.715 331.075 ;
        RECT 1167.625 234.345 1167.795 234.515 ;
        RECT 1167.625 137.785 1167.795 137.955 ;
      LAYER met1 ;
        RECT 1168.470 1683.580 1168.790 1683.640 ;
        RECT 1168.275 1683.440 1168.790 1683.580 ;
        RECT 1168.470 1683.380 1168.790 1683.440 ;
        RECT 1168.470 1635.640 1168.790 1635.700 ;
        RECT 1168.275 1635.500 1168.790 1635.640 ;
        RECT 1168.470 1635.440 1168.790 1635.500 ;
        RECT 1168.470 1587.020 1168.790 1587.080 ;
        RECT 1168.275 1586.880 1168.790 1587.020 ;
        RECT 1168.470 1586.820 1168.790 1586.880 ;
        RECT 1168.470 1539.080 1168.790 1539.140 ;
        RECT 1168.275 1538.940 1168.790 1539.080 ;
        RECT 1168.470 1538.880 1168.790 1538.940 ;
        RECT 1168.470 1490.460 1168.790 1490.520 ;
        RECT 1168.275 1490.320 1168.790 1490.460 ;
        RECT 1168.470 1490.260 1168.790 1490.320 ;
        RECT 1168.470 1442.180 1168.790 1442.240 ;
        RECT 1168.275 1442.040 1168.790 1442.180 ;
        RECT 1168.470 1441.980 1168.790 1442.040 ;
        RECT 1168.470 1345.620 1168.790 1345.680 ;
        RECT 1169.390 1345.620 1169.710 1345.680 ;
        RECT 1168.470 1345.480 1169.710 1345.620 ;
        RECT 1168.470 1345.420 1168.790 1345.480 ;
        RECT 1169.390 1345.420 1169.710 1345.480 ;
        RECT 1168.470 1249.060 1168.790 1249.120 ;
        RECT 1169.390 1249.060 1169.710 1249.120 ;
        RECT 1168.470 1248.920 1169.710 1249.060 ;
        RECT 1168.470 1248.860 1168.790 1248.920 ;
        RECT 1169.390 1248.860 1169.710 1248.920 ;
        RECT 1168.470 1152.500 1168.790 1152.560 ;
        RECT 1169.390 1152.500 1169.710 1152.560 ;
        RECT 1168.470 1152.360 1169.710 1152.500 ;
        RECT 1168.470 1152.300 1168.790 1152.360 ;
        RECT 1169.390 1152.300 1169.710 1152.360 ;
        RECT 1168.470 1007.320 1168.790 1007.380 ;
        RECT 1169.390 1007.320 1169.710 1007.380 ;
        RECT 1168.470 1007.180 1169.710 1007.320 ;
        RECT 1168.470 1007.120 1168.790 1007.180 ;
        RECT 1169.390 1007.120 1169.710 1007.180 ;
        RECT 1168.470 910.760 1168.790 910.820 ;
        RECT 1169.390 910.760 1169.710 910.820 ;
        RECT 1168.470 910.620 1169.710 910.760 ;
        RECT 1168.470 910.560 1168.790 910.620 ;
        RECT 1169.390 910.560 1169.710 910.620 ;
        RECT 1168.470 620.740 1168.790 620.800 ;
        RECT 1168.275 620.600 1168.790 620.740 ;
        RECT 1168.470 620.540 1168.790 620.600 ;
        RECT 1168.470 572.800 1168.790 572.860 ;
        RECT 1168.275 572.660 1168.790 572.800 ;
        RECT 1168.470 572.600 1168.790 572.660 ;
        RECT 1168.470 524.180 1168.790 524.240 ;
        RECT 1168.275 524.040 1168.790 524.180 ;
        RECT 1168.470 523.980 1168.790 524.040 ;
        RECT 1168.470 476.240 1168.790 476.300 ;
        RECT 1168.275 476.100 1168.790 476.240 ;
        RECT 1168.470 476.040 1168.790 476.100 ;
        RECT 1168.470 427.620 1168.790 427.680 ;
        RECT 1168.275 427.480 1168.790 427.620 ;
        RECT 1168.470 427.420 1168.790 427.480 ;
        RECT 1168.470 379.680 1168.790 379.740 ;
        RECT 1168.275 379.540 1168.790 379.680 ;
        RECT 1168.470 379.480 1168.790 379.540 ;
        RECT 1168.470 331.060 1168.790 331.120 ;
        RECT 1168.275 330.920 1168.790 331.060 ;
        RECT 1168.470 330.860 1168.790 330.920 ;
        RECT 1168.470 283.120 1168.790 283.180 ;
        RECT 1168.275 282.980 1168.790 283.120 ;
        RECT 1168.470 282.920 1168.790 282.980 ;
        RECT 1167.565 234.500 1167.855 234.545 ;
        RECT 1168.470 234.500 1168.790 234.560 ;
        RECT 1167.565 234.360 1168.790 234.500 ;
        RECT 1167.565 234.315 1167.855 234.360 ;
        RECT 1168.470 234.300 1168.790 234.360 ;
        RECT 1167.550 186.560 1167.870 186.620 ;
        RECT 1167.355 186.420 1167.870 186.560 ;
        RECT 1167.550 186.360 1167.870 186.420 ;
        RECT 1167.565 137.940 1167.855 137.985 ;
        RECT 1168.470 137.940 1168.790 138.000 ;
        RECT 1167.565 137.800 1168.790 137.940 ;
        RECT 1167.565 137.755 1167.855 137.800 ;
        RECT 1168.470 137.740 1168.790 137.800 ;
        RECT 1167.550 48.520 1167.870 48.580 ;
        RECT 1167.355 48.380 1167.870 48.520 ;
        RECT 1167.550 48.320 1167.870 48.380 ;
      LAYER via ;
        RECT 1168.500 1683.380 1168.760 1683.640 ;
        RECT 1168.500 1635.440 1168.760 1635.700 ;
        RECT 1168.500 1586.820 1168.760 1587.080 ;
        RECT 1168.500 1538.880 1168.760 1539.140 ;
        RECT 1168.500 1490.260 1168.760 1490.520 ;
        RECT 1168.500 1441.980 1168.760 1442.240 ;
        RECT 1168.500 1345.420 1168.760 1345.680 ;
        RECT 1169.420 1345.420 1169.680 1345.680 ;
        RECT 1168.500 1248.860 1168.760 1249.120 ;
        RECT 1169.420 1248.860 1169.680 1249.120 ;
        RECT 1168.500 1152.300 1168.760 1152.560 ;
        RECT 1169.420 1152.300 1169.680 1152.560 ;
        RECT 1168.500 1007.120 1168.760 1007.380 ;
        RECT 1169.420 1007.120 1169.680 1007.380 ;
        RECT 1168.500 910.560 1168.760 910.820 ;
        RECT 1169.420 910.560 1169.680 910.820 ;
        RECT 1168.500 620.540 1168.760 620.800 ;
        RECT 1168.500 572.600 1168.760 572.860 ;
        RECT 1168.500 523.980 1168.760 524.240 ;
        RECT 1168.500 476.040 1168.760 476.300 ;
        RECT 1168.500 427.420 1168.760 427.680 ;
        RECT 1168.500 379.480 1168.760 379.740 ;
        RECT 1168.500 330.860 1168.760 331.120 ;
        RECT 1168.500 282.920 1168.760 283.180 ;
        RECT 1168.500 234.300 1168.760 234.560 ;
        RECT 1167.580 186.360 1167.840 186.620 ;
        RECT 1168.500 137.740 1168.760 138.000 ;
        RECT 1167.580 48.320 1167.840 48.580 ;
      LAYER met2 ;
        RECT 1169.870 1700.410 1170.150 1704.000 ;
        RECT 1168.560 1700.270 1170.150 1700.410 ;
        RECT 1168.560 1683.670 1168.700 1700.270 ;
        RECT 1169.870 1700.000 1170.150 1700.270 ;
        RECT 1168.500 1683.350 1168.760 1683.670 ;
        RECT 1168.500 1635.410 1168.760 1635.730 ;
        RECT 1168.560 1587.110 1168.700 1635.410 ;
        RECT 1168.500 1586.790 1168.760 1587.110 ;
        RECT 1168.500 1538.850 1168.760 1539.170 ;
        RECT 1168.560 1490.550 1168.700 1538.850 ;
        RECT 1168.500 1490.230 1168.760 1490.550 ;
        RECT 1168.500 1441.950 1168.760 1442.270 ;
        RECT 1168.560 1393.845 1168.700 1441.950 ;
        RECT 1168.490 1393.475 1168.770 1393.845 ;
        RECT 1169.410 1393.475 1169.690 1393.845 ;
        RECT 1169.480 1345.710 1169.620 1393.475 ;
        RECT 1168.500 1345.390 1168.760 1345.710 ;
        RECT 1169.420 1345.390 1169.680 1345.710 ;
        RECT 1168.560 1297.285 1168.700 1345.390 ;
        RECT 1168.490 1296.915 1168.770 1297.285 ;
        RECT 1169.410 1296.915 1169.690 1297.285 ;
        RECT 1169.480 1249.150 1169.620 1296.915 ;
        RECT 1168.500 1248.830 1168.760 1249.150 ;
        RECT 1169.420 1248.830 1169.680 1249.150 ;
        RECT 1168.560 1208.885 1168.700 1248.830 ;
        RECT 1168.490 1208.515 1168.770 1208.885 ;
        RECT 1168.490 1207.835 1168.770 1208.205 ;
        RECT 1168.560 1200.725 1168.700 1207.835 ;
        RECT 1168.490 1200.355 1168.770 1200.725 ;
        RECT 1169.410 1200.355 1169.690 1200.725 ;
        RECT 1169.480 1152.590 1169.620 1200.355 ;
        RECT 1168.500 1152.270 1168.760 1152.590 ;
        RECT 1169.420 1152.270 1169.680 1152.590 ;
        RECT 1168.560 1104.165 1168.700 1152.270 ;
        RECT 1168.490 1103.795 1168.770 1104.165 ;
        RECT 1169.410 1103.795 1169.690 1104.165 ;
        RECT 1169.480 1055.885 1169.620 1103.795 ;
        RECT 1168.490 1055.515 1168.770 1055.885 ;
        RECT 1169.410 1055.515 1169.690 1055.885 ;
        RECT 1168.560 1007.410 1168.700 1055.515 ;
        RECT 1168.500 1007.090 1168.760 1007.410 ;
        RECT 1169.420 1007.090 1169.680 1007.410 ;
        RECT 1169.480 959.325 1169.620 1007.090 ;
        RECT 1168.490 958.955 1168.770 959.325 ;
        RECT 1169.410 958.955 1169.690 959.325 ;
        RECT 1168.560 910.850 1168.700 958.955 ;
        RECT 1168.500 910.530 1168.760 910.850 ;
        RECT 1169.420 910.530 1169.680 910.850 ;
        RECT 1169.480 862.765 1169.620 910.530 ;
        RECT 1168.490 862.395 1168.770 862.765 ;
        RECT 1169.410 862.395 1169.690 862.765 ;
        RECT 1168.560 628.845 1168.700 862.395 ;
        RECT 1168.490 628.475 1168.770 628.845 ;
        RECT 1168.490 627.795 1168.770 628.165 ;
        RECT 1168.560 620.830 1168.700 627.795 ;
        RECT 1168.500 620.510 1168.760 620.830 ;
        RECT 1168.500 572.570 1168.760 572.890 ;
        RECT 1168.560 524.270 1168.700 572.570 ;
        RECT 1168.500 523.950 1168.760 524.270 ;
        RECT 1168.500 476.010 1168.760 476.330 ;
        RECT 1168.560 427.710 1168.700 476.010 ;
        RECT 1168.500 427.390 1168.760 427.710 ;
        RECT 1168.500 379.450 1168.760 379.770 ;
        RECT 1168.560 331.150 1168.700 379.450 ;
        RECT 1168.500 330.830 1168.760 331.150 ;
        RECT 1168.500 282.890 1168.760 283.210 ;
        RECT 1168.560 234.590 1168.700 282.890 ;
        RECT 1168.500 234.270 1168.760 234.590 ;
        RECT 1167.580 186.330 1167.840 186.650 ;
        RECT 1167.640 145.365 1167.780 186.330 ;
        RECT 1167.570 144.995 1167.850 145.365 ;
        RECT 1168.490 144.995 1168.770 145.365 ;
        RECT 1168.560 138.030 1168.700 144.995 ;
        RECT 1168.500 137.710 1168.760 138.030 ;
        RECT 1167.580 48.290 1167.840 48.610 ;
        RECT 1167.640 17.525 1167.780 48.290 ;
        RECT 74.150 17.155 74.430 17.525 ;
        RECT 1167.570 17.155 1167.850 17.525 ;
        RECT 74.220 2.400 74.360 17.155 ;
>>>>>>> re-updated local openlane
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 1168.490 1393.520 1168.770 1393.800 ;
        RECT 1169.410 1393.520 1169.690 1393.800 ;
        RECT 1168.490 1296.960 1168.770 1297.240 ;
        RECT 1169.410 1296.960 1169.690 1297.240 ;
        RECT 1168.490 1208.560 1168.770 1208.840 ;
        RECT 1168.490 1207.880 1168.770 1208.160 ;
        RECT 1168.490 1200.400 1168.770 1200.680 ;
        RECT 1169.410 1200.400 1169.690 1200.680 ;
        RECT 1168.490 1103.840 1168.770 1104.120 ;
        RECT 1169.410 1103.840 1169.690 1104.120 ;
        RECT 1168.490 1055.560 1168.770 1055.840 ;
        RECT 1169.410 1055.560 1169.690 1055.840 ;
        RECT 1168.490 959.000 1168.770 959.280 ;
        RECT 1169.410 959.000 1169.690 959.280 ;
        RECT 1168.490 862.440 1168.770 862.720 ;
        RECT 1169.410 862.440 1169.690 862.720 ;
        RECT 1168.490 628.520 1168.770 628.800 ;
        RECT 1168.490 627.840 1168.770 628.120 ;
        RECT 1167.570 145.040 1167.850 145.320 ;
        RECT 1168.490 145.040 1168.770 145.320 ;
        RECT 74.150 17.200 74.430 17.480 ;
        RECT 1167.570 17.200 1167.850 17.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 74.125 18.850 74.455 18.865 ;
        RECT 1168.925 18.850 1169.255 18.865 ;
        RECT 74.125 18.550 1169.255 18.850 ;
        RECT 74.125 18.535 74.455 18.550 ;
        RECT 1168.925 18.535 1169.255 18.550 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1168.465 1393.810 1168.795 1393.825 ;
        RECT 1169.385 1393.810 1169.715 1393.825 ;
        RECT 1168.465 1393.510 1169.715 1393.810 ;
        RECT 1168.465 1393.495 1168.795 1393.510 ;
        RECT 1169.385 1393.495 1169.715 1393.510 ;
        RECT 1168.465 1297.250 1168.795 1297.265 ;
        RECT 1169.385 1297.250 1169.715 1297.265 ;
        RECT 1168.465 1296.950 1169.715 1297.250 ;
        RECT 1168.465 1296.935 1168.795 1296.950 ;
        RECT 1169.385 1296.935 1169.715 1296.950 ;
        RECT 1168.465 1208.850 1168.795 1208.865 ;
        RECT 1167.790 1208.550 1168.795 1208.850 ;
        RECT 1167.790 1208.170 1168.090 1208.550 ;
        RECT 1168.465 1208.535 1168.795 1208.550 ;
        RECT 1168.465 1208.170 1168.795 1208.185 ;
        RECT 1167.790 1207.870 1168.795 1208.170 ;
        RECT 1168.465 1207.855 1168.795 1207.870 ;
        RECT 1168.465 1200.690 1168.795 1200.705 ;
        RECT 1169.385 1200.690 1169.715 1200.705 ;
        RECT 1168.465 1200.390 1169.715 1200.690 ;
        RECT 1168.465 1200.375 1168.795 1200.390 ;
        RECT 1169.385 1200.375 1169.715 1200.390 ;
        RECT 1168.465 1104.130 1168.795 1104.145 ;
        RECT 1169.385 1104.130 1169.715 1104.145 ;
        RECT 1168.465 1103.830 1169.715 1104.130 ;
        RECT 1168.465 1103.815 1168.795 1103.830 ;
        RECT 1169.385 1103.815 1169.715 1103.830 ;
        RECT 1168.465 1055.850 1168.795 1055.865 ;
        RECT 1169.385 1055.850 1169.715 1055.865 ;
        RECT 1168.465 1055.550 1169.715 1055.850 ;
        RECT 1168.465 1055.535 1168.795 1055.550 ;
        RECT 1169.385 1055.535 1169.715 1055.550 ;
        RECT 1168.465 959.290 1168.795 959.305 ;
        RECT 1169.385 959.290 1169.715 959.305 ;
        RECT 1168.465 958.990 1169.715 959.290 ;
        RECT 1168.465 958.975 1168.795 958.990 ;
        RECT 1169.385 958.975 1169.715 958.990 ;
        RECT 1168.465 862.730 1168.795 862.745 ;
        RECT 1169.385 862.730 1169.715 862.745 ;
        RECT 1168.465 862.430 1169.715 862.730 ;
        RECT 1168.465 862.415 1168.795 862.430 ;
        RECT 1169.385 862.415 1169.715 862.430 ;
        RECT 1168.465 628.810 1168.795 628.825 ;
        RECT 1168.465 628.495 1169.010 628.810 ;
        RECT 1168.710 628.145 1169.010 628.495 ;
        RECT 1168.465 627.830 1169.010 628.145 ;
        RECT 1168.465 627.815 1168.795 627.830 ;
        RECT 1167.545 145.330 1167.875 145.345 ;
        RECT 1168.465 145.330 1168.795 145.345 ;
        RECT 1167.545 145.030 1168.795 145.330 ;
        RECT 1167.545 145.015 1167.875 145.030 ;
        RECT 1168.465 145.015 1168.795 145.030 ;
        RECT 74.125 17.490 74.455 17.505 ;
        RECT 1167.545 17.490 1167.875 17.505 ;
        RECT 74.125 17.190 1167.875 17.490 ;
        RECT 74.125 17.175 74.455 17.190 ;
        RECT 1167.545 17.175 1167.875 17.190 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 0.300 ;
=======
      LAYER met1 ;
        RECT 1264.150 16.560 1264.470 16.620 ;
        RECT 448.200 16.420 1264.470 16.560 ;
        RECT 430.630 16.220 430.950 16.280 ;
        RECT 448.200 16.220 448.340 16.420 ;
        RECT 1264.150 16.360 1264.470 16.420 ;
        RECT 430.630 16.080 448.340 16.220 ;
        RECT 430.630 16.020 430.950 16.080 ;
      LAYER via ;
        RECT 430.660 16.020 430.920 16.280 ;
        RECT 1264.180 16.360 1264.440 16.620 ;
      LAYER met2 ;
        RECT 1266.470 1700.410 1266.750 1704.000 ;
        RECT 1265.160 1700.270 1266.750 1700.410 ;
        RECT 1265.160 1677.970 1265.300 1700.270 ;
        RECT 1266.470 1700.000 1266.750 1700.270 ;
        RECT 1264.240 1677.830 1265.300 1677.970 ;
        RECT 1264.240 16.650 1264.380 1677.830 ;
        RECT 1264.180 16.330 1264.440 16.650 ;
        RECT 430.660 15.990 430.920 16.310 ;
        RECT 430.720 2.400 430.860 15.990 ;
        RECT 430.510 -4.800 431.070 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 0.300 ;
=======
      LAYER met1 ;
        RECT 448.570 16.220 448.890 16.280 ;
        RECT 1270.130 16.220 1270.450 16.280 ;
        RECT 448.570 16.080 1270.450 16.220 ;
        RECT 448.570 16.020 448.890 16.080 ;
        RECT 1270.130 16.020 1270.450 16.080 ;
      LAYER via ;
        RECT 448.600 16.020 448.860 16.280 ;
        RECT 1270.160 16.020 1270.420 16.280 ;
      LAYER met2 ;
        RECT 1271.070 1700.410 1271.350 1704.000 ;
        RECT 1270.220 1700.270 1271.350 1700.410 ;
        RECT 1270.220 16.310 1270.360 1700.270 ;
        RECT 1271.070 1700.000 1271.350 1700.270 ;
        RECT 448.600 15.990 448.860 16.310 ;
        RECT 1270.160 15.990 1270.420 16.310 ;
        RECT 448.660 2.400 448.800 15.990 ;
        RECT 448.450 -4.800 449.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 0.300 ;
=======
      LAYER met1 ;
        RECT 1271.510 1659.100 1271.830 1659.160 ;
        RECT 1274.730 1659.100 1275.050 1659.160 ;
        RECT 1271.510 1658.960 1275.050 1659.100 ;
        RECT 1271.510 1658.900 1271.830 1658.960 ;
        RECT 1274.730 1658.900 1275.050 1658.960 ;
        RECT 466.510 15.880 466.830 15.940 ;
        RECT 1271.510 15.880 1271.830 15.940 ;
        RECT 466.510 15.740 1271.830 15.880 ;
        RECT 466.510 15.680 466.830 15.740 ;
        RECT 1271.510 15.680 1271.830 15.740 ;
      LAYER via ;
        RECT 1271.540 1658.900 1271.800 1659.160 ;
        RECT 1274.760 1658.900 1275.020 1659.160 ;
        RECT 466.540 15.680 466.800 15.940 ;
        RECT 1271.540 15.680 1271.800 15.940 ;
      LAYER met2 ;
        RECT 1276.130 1700.410 1276.410 1704.000 ;
        RECT 1274.820 1700.270 1276.410 1700.410 ;
        RECT 1274.820 1659.190 1274.960 1700.270 ;
        RECT 1276.130 1700.000 1276.410 1700.270 ;
        RECT 1271.540 1658.870 1271.800 1659.190 ;
        RECT 1274.760 1658.870 1275.020 1659.190 ;
        RECT 1271.600 15.970 1271.740 1658.870 ;
        RECT 466.540 15.650 466.800 15.970 ;
        RECT 1271.540 15.650 1271.800 15.970 ;
        RECT 466.600 2.400 466.740 15.650 ;
        RECT 466.390 -4.800 466.950 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 0.300 ;
=======
      LAYER met1 ;
        RECT 489.510 1686.300 489.830 1686.360 ;
        RECT 1280.250 1686.300 1280.570 1686.360 ;
        RECT 489.510 1686.160 1280.570 1686.300 ;
        RECT 489.510 1686.100 489.830 1686.160 ;
        RECT 1280.250 1686.100 1280.570 1686.160 ;
        RECT 484.450 15.880 484.770 15.940 ;
        RECT 489.510 15.880 489.830 15.940 ;
        RECT 484.450 15.740 489.830 15.880 ;
        RECT 484.450 15.680 484.770 15.740 ;
        RECT 489.510 15.680 489.830 15.740 ;
      LAYER via ;
        RECT 489.540 1686.100 489.800 1686.360 ;
        RECT 1280.280 1686.100 1280.540 1686.360 ;
        RECT 484.480 15.680 484.740 15.940 ;
        RECT 489.540 15.680 489.800 15.940 ;
      LAYER met2 ;
        RECT 1280.270 1700.000 1280.550 1704.000 ;
        RECT 1280.340 1686.390 1280.480 1700.000 ;
        RECT 489.540 1686.070 489.800 1686.390 ;
        RECT 1280.280 1686.070 1280.540 1686.390 ;
        RECT 489.600 15.970 489.740 1686.070 ;
        RECT 484.480 15.650 484.740 15.970 ;
        RECT 489.540 15.650 489.800 15.970 ;
        RECT 484.540 2.400 484.680 15.650 ;
        RECT 484.330 -4.800 484.890 2.400 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER li1 ;
        RECT 1278.945 1558.985 1279.115 1593.835 ;
        RECT 1278.025 1261.485 1278.195 1304.155 ;
        RECT 1278.025 908.565 1278.195 959.055 ;
        RECT 1278.025 848.725 1278.195 896.835 ;
        RECT 1278.025 589.985 1278.195 627.895 ;
        RECT 1278.485 510.765 1278.655 558.875 ;
      LAYER mcon ;
        RECT 1278.945 1593.665 1279.115 1593.835 ;
        RECT 1278.025 1303.985 1278.195 1304.155 ;
        RECT 1278.025 958.885 1278.195 959.055 ;
        RECT 1278.025 896.665 1278.195 896.835 ;
        RECT 1278.025 627.725 1278.195 627.895 ;
        RECT 1278.485 558.705 1278.655 558.875 ;
      LAYER met1 ;
        RECT 1278.870 1593.820 1279.190 1593.880 ;
        RECT 1278.675 1593.680 1279.190 1593.820 ;
        RECT 1278.870 1593.620 1279.190 1593.680 ;
        RECT 1278.885 1559.140 1279.175 1559.185 ;
        RECT 1279.330 1559.140 1279.650 1559.200 ;
        RECT 1278.885 1559.000 1279.650 1559.140 ;
        RECT 1278.885 1558.955 1279.175 1559.000 ;
        RECT 1279.330 1558.940 1279.650 1559.000 ;
        RECT 1277.950 1414.440 1278.270 1414.700 ;
        RECT 1278.040 1413.960 1278.180 1414.440 ;
        RECT 1278.410 1413.960 1278.730 1414.020 ;
        RECT 1278.040 1413.820 1278.730 1413.960 ;
        RECT 1278.410 1413.760 1278.730 1413.820 ;
        RECT 1276.570 1400.700 1276.890 1400.760 ;
        RECT 1278.410 1400.700 1278.730 1400.760 ;
        RECT 1276.570 1400.560 1278.730 1400.700 ;
        RECT 1276.570 1400.500 1276.890 1400.560 ;
        RECT 1278.410 1400.500 1278.730 1400.560 ;
        RECT 1278.410 1317.880 1278.730 1318.140 ;
        RECT 1278.500 1317.460 1278.640 1317.880 ;
        RECT 1278.410 1317.200 1278.730 1317.460 ;
        RECT 1277.965 1304.140 1278.255 1304.185 ;
        RECT 1278.410 1304.140 1278.730 1304.200 ;
        RECT 1277.965 1304.000 1278.730 1304.140 ;
        RECT 1277.965 1303.955 1278.255 1304.000 ;
        RECT 1278.410 1303.940 1278.730 1304.000 ;
        RECT 1277.950 1261.640 1278.270 1261.700 ;
        RECT 1277.755 1261.500 1278.270 1261.640 ;
        RECT 1277.950 1261.440 1278.270 1261.500 ;
        RECT 1277.950 1221.320 1278.270 1221.580 ;
        RECT 1278.040 1220.840 1278.180 1221.320 ;
        RECT 1278.410 1220.840 1278.730 1220.900 ;
        RECT 1278.040 1220.700 1278.730 1220.840 ;
        RECT 1278.410 1220.640 1278.730 1220.700 ;
        RECT 1278.410 1200.440 1278.730 1200.500 ;
        RECT 1279.330 1200.440 1279.650 1200.500 ;
        RECT 1278.410 1200.300 1279.650 1200.440 ;
        RECT 1278.410 1200.240 1278.730 1200.300 ;
        RECT 1279.330 1200.240 1279.650 1200.300 ;
        RECT 1278.410 1031.460 1278.730 1031.520 ;
        RECT 1279.330 1031.460 1279.650 1031.520 ;
        RECT 1278.410 1031.320 1279.650 1031.460 ;
        RECT 1278.410 1031.260 1278.730 1031.320 ;
        RECT 1279.330 1031.260 1279.650 1031.320 ;
        RECT 1277.965 959.040 1278.255 959.085 ;
        RECT 1278.870 959.040 1279.190 959.100 ;
        RECT 1277.965 958.900 1279.190 959.040 ;
        RECT 1277.965 958.855 1278.255 958.900 ;
        RECT 1278.870 958.840 1279.190 958.900 ;
        RECT 1277.950 908.720 1278.270 908.780 ;
        RECT 1277.755 908.580 1278.270 908.720 ;
        RECT 1277.950 908.520 1278.270 908.580 ;
        RECT 1277.950 896.820 1278.270 896.880 ;
        RECT 1277.755 896.680 1278.270 896.820 ;
        RECT 1277.950 896.620 1278.270 896.680 ;
        RECT 1277.950 848.880 1278.270 848.940 ;
        RECT 1277.755 848.740 1278.270 848.880 ;
        RECT 1277.950 848.680 1278.270 848.740 ;
        RECT 1277.950 807.060 1278.270 807.120 ;
        RECT 1278.410 807.060 1278.730 807.120 ;
        RECT 1277.950 806.920 1278.730 807.060 ;
        RECT 1277.950 806.860 1278.270 806.920 ;
        RECT 1278.410 806.860 1278.730 806.920 ;
        RECT 1277.950 725.260 1278.270 725.520 ;
        RECT 1278.040 724.840 1278.180 725.260 ;
        RECT 1277.950 724.580 1278.270 724.840 ;
        RECT 1277.950 717.640 1278.270 717.700 ;
        RECT 1278.870 717.640 1279.190 717.700 ;
        RECT 1277.950 717.500 1279.190 717.640 ;
        RECT 1277.950 717.440 1278.270 717.500 ;
        RECT 1278.870 717.440 1279.190 717.500 ;
        RECT 1277.965 627.880 1278.255 627.925 ;
        RECT 1278.410 627.880 1278.730 627.940 ;
        RECT 1277.965 627.740 1278.730 627.880 ;
        RECT 1277.965 627.695 1278.255 627.740 ;
        RECT 1278.410 627.680 1278.730 627.740 ;
        RECT 1277.965 590.140 1278.255 590.185 ;
        RECT 1278.870 590.140 1279.190 590.200 ;
        RECT 1277.965 590.000 1279.190 590.140 ;
        RECT 1277.965 589.955 1278.255 590.000 ;
        RECT 1278.870 589.940 1279.190 590.000 ;
        RECT 1278.425 558.860 1278.715 558.905 ;
        RECT 1278.870 558.860 1279.190 558.920 ;
        RECT 1278.425 558.720 1279.190 558.860 ;
        RECT 1278.425 558.675 1278.715 558.720 ;
        RECT 1278.870 558.660 1279.190 558.720 ;
        RECT 1278.410 510.920 1278.730 510.980 ;
        RECT 1278.215 510.780 1278.730 510.920 ;
        RECT 1278.410 510.720 1278.730 510.780 ;
        RECT 1277.950 421.300 1278.270 421.560 ;
        RECT 1276.570 420.820 1276.890 420.880 ;
        RECT 1278.040 420.820 1278.180 421.300 ;
        RECT 1276.570 420.680 1278.180 420.820 ;
        RECT 1276.570 420.620 1276.890 420.680 ;
        RECT 1277.950 317.460 1278.270 317.520 ;
        RECT 1279.330 317.460 1279.650 317.520 ;
        RECT 1277.950 317.320 1279.650 317.460 ;
        RECT 1277.950 317.260 1278.270 317.320 ;
        RECT 1279.330 317.260 1279.650 317.320 ;
        RECT 1277.950 251.840 1278.270 251.900 ;
        RECT 1279.330 251.840 1279.650 251.900 ;
        RECT 1277.950 251.700 1279.650 251.840 ;
        RECT 1277.950 251.640 1278.270 251.700 ;
        RECT 1279.330 251.640 1279.650 251.700 ;
        RECT 1277.950 15.540 1278.270 15.600 ;
        RECT 541.580 15.400 1278.270 15.540 ;
        RECT 484.450 15.200 484.770 15.260 ;
        RECT 541.580 15.200 541.720 15.400 ;
        RECT 1277.950 15.340 1278.270 15.400 ;
        RECT 484.450 15.060 541.720 15.200 ;
        RECT 484.450 15.000 484.770 15.060 ;
      LAYER via ;
        RECT 1278.900 1593.620 1279.160 1593.880 ;
        RECT 1279.360 1558.940 1279.620 1559.200 ;
        RECT 1277.980 1414.440 1278.240 1414.700 ;
        RECT 1278.440 1413.760 1278.700 1414.020 ;
        RECT 1276.600 1400.500 1276.860 1400.760 ;
        RECT 1278.440 1400.500 1278.700 1400.760 ;
        RECT 1278.440 1317.880 1278.700 1318.140 ;
        RECT 1278.440 1317.200 1278.700 1317.460 ;
        RECT 1278.440 1303.940 1278.700 1304.200 ;
        RECT 1277.980 1261.440 1278.240 1261.700 ;
        RECT 1277.980 1221.320 1278.240 1221.580 ;
        RECT 1278.440 1220.640 1278.700 1220.900 ;
        RECT 1278.440 1200.240 1278.700 1200.500 ;
        RECT 1279.360 1200.240 1279.620 1200.500 ;
        RECT 1278.440 1031.260 1278.700 1031.520 ;
        RECT 1279.360 1031.260 1279.620 1031.520 ;
        RECT 1278.900 958.840 1279.160 959.100 ;
        RECT 1277.980 908.520 1278.240 908.780 ;
        RECT 1277.980 896.620 1278.240 896.880 ;
        RECT 1277.980 848.680 1278.240 848.940 ;
        RECT 1277.980 806.860 1278.240 807.120 ;
        RECT 1278.440 806.860 1278.700 807.120 ;
        RECT 1277.980 725.260 1278.240 725.520 ;
        RECT 1277.980 724.580 1278.240 724.840 ;
        RECT 1277.980 717.440 1278.240 717.700 ;
        RECT 1278.900 717.440 1279.160 717.700 ;
        RECT 1278.440 627.680 1278.700 627.940 ;
        RECT 1278.900 589.940 1279.160 590.200 ;
        RECT 1278.900 558.660 1279.160 558.920 ;
        RECT 1278.440 510.720 1278.700 510.980 ;
        RECT 1277.980 421.300 1278.240 421.560 ;
        RECT 1276.600 420.620 1276.860 420.880 ;
        RECT 1277.980 317.260 1278.240 317.520 ;
        RECT 1279.360 317.260 1279.620 317.520 ;
        RECT 1277.980 251.640 1278.240 251.900 ;
        RECT 1279.360 251.640 1279.620 251.900 ;
        RECT 484.480 15.000 484.740 15.260 ;
        RECT 1277.980 15.340 1278.240 15.600 ;
      LAYER met2 ;
        RECT 1280.730 1700.410 1281.010 1704.000 ;
        RECT 1280.340 1700.270 1281.010 1700.410 ;
        RECT 1280.340 1656.210 1280.480 1700.270 ;
        RECT 1280.730 1700.000 1281.010 1700.270 ;
        RECT 1279.420 1656.070 1280.480 1656.210 ;
        RECT 1279.420 1594.330 1279.560 1656.070 ;
        RECT 1278.960 1594.190 1279.560 1594.330 ;
        RECT 1278.960 1593.910 1279.100 1594.190 ;
        RECT 1278.900 1593.590 1279.160 1593.910 ;
        RECT 1279.360 1558.910 1279.620 1559.230 ;
        RECT 1279.420 1463.090 1279.560 1558.910 ;
        RECT 1278.040 1462.950 1279.560 1463.090 ;
        RECT 1278.040 1414.730 1278.180 1462.950 ;
        RECT 1277.980 1414.410 1278.240 1414.730 ;
        RECT 1278.440 1413.730 1278.700 1414.050 ;
        RECT 1278.500 1400.790 1278.640 1413.730 ;
        RECT 1276.600 1400.470 1276.860 1400.790 ;
        RECT 1278.440 1400.470 1278.700 1400.790 ;
        RECT 1276.660 1353.045 1276.800 1400.470 ;
        RECT 1276.590 1352.675 1276.870 1353.045 ;
        RECT 1278.430 1351.995 1278.710 1352.365 ;
        RECT 1278.500 1318.170 1278.640 1351.995 ;
        RECT 1278.440 1317.850 1278.700 1318.170 ;
        RECT 1278.440 1317.170 1278.700 1317.490 ;
        RECT 1278.500 1304.230 1278.640 1317.170 ;
        RECT 1278.440 1303.910 1278.700 1304.230 ;
        RECT 1277.980 1261.410 1278.240 1261.730 ;
        RECT 1278.040 1221.610 1278.180 1261.410 ;
        RECT 1277.980 1221.290 1278.240 1221.610 ;
        RECT 1278.440 1220.610 1278.700 1220.930 ;
        RECT 1278.500 1200.530 1278.640 1220.610 ;
        RECT 1278.440 1200.210 1278.700 1200.530 ;
        RECT 1279.360 1200.210 1279.620 1200.530 ;
        RECT 1279.420 1152.445 1279.560 1200.210 ;
        RECT 1278.430 1152.075 1278.710 1152.445 ;
        RECT 1279.350 1152.075 1279.630 1152.445 ;
        RECT 1278.500 1031.550 1278.640 1152.075 ;
        RECT 1278.440 1031.230 1278.700 1031.550 ;
        RECT 1279.360 1031.230 1279.620 1031.550 ;
        RECT 1279.420 1007.605 1279.560 1031.230 ;
        RECT 1278.430 1007.235 1278.710 1007.605 ;
        RECT 1279.350 1007.235 1279.630 1007.605 ;
        RECT 1278.500 983.010 1278.640 1007.235 ;
        RECT 1278.500 982.870 1279.100 983.010 ;
        RECT 1278.960 959.130 1279.100 982.870 ;
        RECT 1278.900 958.810 1279.160 959.130 ;
        RECT 1277.980 908.490 1278.240 908.810 ;
        RECT 1278.040 896.910 1278.180 908.490 ;
        RECT 1277.980 896.590 1278.240 896.910 ;
        RECT 1277.980 848.650 1278.240 848.970 ;
        RECT 1278.040 835.450 1278.180 848.650 ;
        RECT 1278.040 835.310 1278.640 835.450 ;
        RECT 1278.500 807.150 1278.640 835.310 ;
        RECT 1277.980 806.830 1278.240 807.150 ;
        RECT 1278.440 806.830 1278.700 807.150 ;
        RECT 1278.040 725.550 1278.180 806.830 ;
        RECT 1277.980 725.230 1278.240 725.550 ;
        RECT 1277.980 724.550 1278.240 724.870 ;
        RECT 1278.040 717.730 1278.180 724.550 ;
        RECT 1277.980 717.410 1278.240 717.730 ;
        RECT 1278.900 717.410 1279.160 717.730 ;
        RECT 1278.960 641.650 1279.100 717.410 ;
        RECT 1278.500 641.510 1279.100 641.650 ;
        RECT 1278.500 627.970 1278.640 641.510 ;
        RECT 1278.440 627.650 1278.700 627.970 ;
        RECT 1278.900 589.910 1279.160 590.230 ;
        RECT 1278.960 558.950 1279.100 589.910 ;
        RECT 1278.900 558.630 1279.160 558.950 ;
        RECT 1278.440 510.690 1278.700 511.010 ;
        RECT 1278.500 510.410 1278.640 510.690 ;
        RECT 1278.040 510.270 1278.640 510.410 ;
        RECT 1278.040 421.590 1278.180 510.270 ;
        RECT 1277.980 421.270 1278.240 421.590 ;
        RECT 1276.600 420.590 1276.860 420.910 ;
        RECT 1276.660 373.165 1276.800 420.590 ;
        RECT 1276.590 372.795 1276.870 373.165 ;
        RECT 1276.590 372.115 1276.870 372.485 ;
        RECT 1276.660 324.885 1276.800 372.115 ;
        RECT 1276.590 324.515 1276.870 324.885 ;
        RECT 1277.970 324.515 1278.250 324.885 ;
        RECT 1278.040 317.550 1278.180 324.515 ;
        RECT 1277.980 317.230 1278.240 317.550 ;
        RECT 1279.360 317.230 1279.620 317.550 ;
        RECT 1279.420 251.930 1279.560 317.230 ;
        RECT 1277.980 251.610 1278.240 251.930 ;
        RECT 1279.360 251.610 1279.620 251.930 ;
        RECT 1278.040 158.170 1278.180 251.610 ;
        RECT 1278.040 158.030 1278.640 158.170 ;
        RECT 1278.500 62.290 1278.640 158.030 ;
        RECT 1278.040 62.150 1278.640 62.290 ;
        RECT 1278.040 15.630 1278.180 62.150 ;
        RECT 1277.980 15.310 1278.240 15.630 ;
        RECT 484.480 14.970 484.740 15.290 ;
        RECT 484.540 2.400 484.680 14.970 ;
        RECT 484.330 -4.800 484.890 2.400 ;
      LAYER via2 ;
        RECT 1276.590 1352.720 1276.870 1353.000 ;
        RECT 1278.430 1352.040 1278.710 1352.320 ;
        RECT 1278.430 1152.120 1278.710 1152.400 ;
        RECT 1279.350 1152.120 1279.630 1152.400 ;
        RECT 1278.430 1007.280 1278.710 1007.560 ;
        RECT 1279.350 1007.280 1279.630 1007.560 ;
        RECT 1276.590 372.840 1276.870 373.120 ;
        RECT 1276.590 372.160 1276.870 372.440 ;
        RECT 1276.590 324.560 1276.870 324.840 ;
        RECT 1277.970 324.560 1278.250 324.840 ;
      LAYER met3 ;
        RECT 1276.565 1353.010 1276.895 1353.025 ;
        RECT 1276.565 1352.710 1277.570 1353.010 ;
        RECT 1276.565 1352.695 1276.895 1352.710 ;
        RECT 1277.270 1352.330 1277.570 1352.710 ;
        RECT 1278.405 1352.330 1278.735 1352.345 ;
        RECT 1277.270 1352.030 1278.735 1352.330 ;
        RECT 1278.405 1352.015 1278.735 1352.030 ;
        RECT 1278.405 1152.410 1278.735 1152.425 ;
        RECT 1279.325 1152.410 1279.655 1152.425 ;
        RECT 1278.405 1152.110 1279.655 1152.410 ;
        RECT 1278.405 1152.095 1278.735 1152.110 ;
        RECT 1279.325 1152.095 1279.655 1152.110 ;
        RECT 1278.405 1007.570 1278.735 1007.585 ;
        RECT 1279.325 1007.570 1279.655 1007.585 ;
        RECT 1278.405 1007.270 1279.655 1007.570 ;
        RECT 1278.405 1007.255 1278.735 1007.270 ;
        RECT 1279.325 1007.255 1279.655 1007.270 ;
        RECT 1276.565 373.130 1276.895 373.145 ;
        RECT 1276.565 372.830 1277.570 373.130 ;
        RECT 1276.565 372.815 1276.895 372.830 ;
        RECT 1276.565 372.450 1276.895 372.465 ;
        RECT 1277.270 372.450 1277.570 372.830 ;
        RECT 1276.565 372.150 1277.570 372.450 ;
        RECT 1276.565 372.135 1276.895 372.150 ;
        RECT 1276.565 324.850 1276.895 324.865 ;
        RECT 1277.945 324.850 1278.275 324.865 ;
        RECT 1276.565 324.550 1278.275 324.850 ;
        RECT 1276.565 324.535 1276.895 324.550 ;
        RECT 1277.945 324.535 1278.275 324.550 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 0.300 ;
=======
      LAYER met1 ;
        RECT 503.310 1689.700 503.630 1689.760 ;
        RECT 1285.770 1689.700 1286.090 1689.760 ;
        RECT 503.310 1689.560 1286.090 1689.700 ;
        RECT 503.310 1689.500 503.630 1689.560 ;
        RECT 1285.770 1689.500 1286.090 1689.560 ;
      LAYER via ;
        RECT 503.340 1689.500 503.600 1689.760 ;
        RECT 1285.800 1689.500 1286.060 1689.760 ;
      LAYER met2 ;
        RECT 1285.790 1700.000 1286.070 1704.000 ;
        RECT 1285.860 1689.790 1286.000 1700.000 ;
        RECT 503.340 1689.470 503.600 1689.790 ;
        RECT 1285.800 1689.470 1286.060 1689.790 ;
        RECT 503.400 3.130 503.540 1689.470 ;
        RECT 502.480 2.990 503.540 3.130 ;
        RECT 502.480 2.400 502.620 2.990 ;
        RECT 502.270 -4.800 502.830 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 0.300 ;
=======
      LAYER met1 ;
        RECT 1291.750 15.200 1292.070 15.260 ;
        RECT 542.040 15.060 1292.070 15.200 ;
        RECT 519.870 14.860 520.190 14.920 ;
        RECT 542.040 14.860 542.180 15.060 ;
        RECT 1291.750 15.000 1292.070 15.060 ;
        RECT 519.870 14.720 542.180 14.860 ;
        RECT 519.870 14.660 520.190 14.720 ;
      LAYER via ;
        RECT 519.900 14.660 520.160 14.920 ;
        RECT 1291.780 15.000 1292.040 15.260 ;
      LAYER met2 ;
        RECT 1290.850 1700.410 1291.130 1704.000 ;
        RECT 1290.850 1700.270 1291.980 1700.410 ;
        RECT 1290.850 1700.000 1291.130 1700.270 ;
        RECT 1291.840 15.290 1291.980 1700.270 ;
        RECT 1291.780 14.970 1292.040 15.290 ;
        RECT 519.900 14.630 520.160 14.950 ;
        RECT 519.960 2.400 520.100 14.630 ;
        RECT 519.750 -4.800 520.310 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 0.300 ;
=======
      LAYER met1 ;
        RECT 537.810 1690.040 538.130 1690.100 ;
        RECT 1295.430 1690.040 1295.750 1690.100 ;
        RECT 537.810 1689.900 1295.750 1690.040 ;
        RECT 537.810 1689.840 538.130 1689.900 ;
        RECT 1295.430 1689.840 1295.750 1689.900 ;
      LAYER via ;
        RECT 537.840 1689.840 538.100 1690.100 ;
        RECT 1295.460 1689.840 1295.720 1690.100 ;
      LAYER met2 ;
        RECT 1295.450 1700.000 1295.730 1704.000 ;
        RECT 1295.520 1690.130 1295.660 1700.000 ;
        RECT 537.840 1689.810 538.100 1690.130 ;
        RECT 1295.460 1689.810 1295.720 1690.130 ;
        RECT 537.900 2.400 538.040 1689.810 ;
        RECT 537.690 -4.800 538.250 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 0.300 ;
=======
      LAYER met1 ;
        RECT 1298.650 14.860 1298.970 14.920 ;
        RECT 607.360 14.720 1298.970 14.860 ;
        RECT 555.750 14.520 556.070 14.580 ;
        RECT 607.360 14.520 607.500 14.720 ;
        RECT 1298.650 14.660 1298.970 14.720 ;
        RECT 555.750 14.380 607.500 14.520 ;
        RECT 555.750 14.320 556.070 14.380 ;
      LAYER via ;
        RECT 555.780 14.320 556.040 14.580 ;
        RECT 1298.680 14.660 1298.940 14.920 ;
      LAYER met2 ;
        RECT 1300.510 1700.410 1300.790 1704.000 ;
        RECT 1299.200 1700.270 1300.790 1700.410 ;
        RECT 1299.200 18.770 1299.340 1700.270 ;
        RECT 1300.510 1700.000 1300.790 1700.270 ;
        RECT 1298.740 18.630 1299.340 18.770 ;
        RECT 1298.740 14.950 1298.880 18.630 ;
        RECT 1298.680 14.630 1298.940 14.950 ;
        RECT 555.780 14.290 556.040 14.610 ;
        RECT 555.840 2.400 555.980 14.290 ;
        RECT 555.630 -4.800 556.190 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 0.300 ;
=======
      LAYER met1 ;
        RECT 579.210 1686.640 579.530 1686.700 ;
        RECT 1305.090 1686.640 1305.410 1686.700 ;
        RECT 579.210 1686.500 1305.410 1686.640 ;
        RECT 579.210 1686.440 579.530 1686.500 ;
        RECT 1305.090 1686.440 1305.410 1686.500 ;
        RECT 573.690 14.860 574.010 14.920 ;
        RECT 579.210 14.860 579.530 14.920 ;
        RECT 573.690 14.720 579.530 14.860 ;
        RECT 573.690 14.660 574.010 14.720 ;
        RECT 579.210 14.660 579.530 14.720 ;
      LAYER via ;
        RECT 579.240 1686.440 579.500 1686.700 ;
        RECT 1305.120 1686.440 1305.380 1686.700 ;
        RECT 573.720 14.660 573.980 14.920 ;
        RECT 579.240 14.660 579.500 14.920 ;
      LAYER met2 ;
        RECT 1305.110 1700.000 1305.390 1704.000 ;
        RECT 1305.180 1686.730 1305.320 1700.000 ;
        RECT 579.240 1686.410 579.500 1686.730 ;
        RECT 1305.120 1686.410 1305.380 1686.730 ;
        RECT 579.300 14.950 579.440 1686.410 ;
        RECT 573.720 14.630 573.980 14.950 ;
        RECT 579.240 14.630 579.500 14.950 ;
        RECT 573.780 2.400 573.920 14.630 ;
        RECT 573.570 -4.800 574.130 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 0.300 ;
=======
      LAYER met1 ;
        RECT 1305.550 1677.460 1305.870 1677.520 ;
        RECT 1308.770 1677.460 1309.090 1677.520 ;
        RECT 1305.550 1677.320 1309.090 1677.460 ;
        RECT 1305.550 1677.260 1305.870 1677.320 ;
        RECT 1308.770 1677.260 1309.090 1677.320 ;
        RECT 1305.550 14.520 1305.870 14.580 ;
        RECT 607.820 14.380 1305.870 14.520 ;
        RECT 591.170 14.180 591.490 14.240 ;
        RECT 607.820 14.180 607.960 14.380 ;
        RECT 1305.550 14.320 1305.870 14.380 ;
        RECT 591.170 14.040 607.960 14.180 ;
        RECT 591.170 13.980 591.490 14.040 ;
      LAYER via ;
        RECT 1305.580 1677.260 1305.840 1677.520 ;
        RECT 1308.800 1677.260 1309.060 1677.520 ;
        RECT 591.200 13.980 591.460 14.240 ;
        RECT 1305.580 14.320 1305.840 14.580 ;
      LAYER met2 ;
        RECT 1310.170 1700.410 1310.450 1704.000 ;
        RECT 1308.860 1700.270 1310.450 1700.410 ;
        RECT 1308.860 1677.550 1309.000 1700.270 ;
        RECT 1310.170 1700.000 1310.450 1700.270 ;
        RECT 1305.580 1677.230 1305.840 1677.550 ;
        RECT 1308.800 1677.230 1309.060 1677.550 ;
        RECT 1305.640 14.610 1305.780 1677.230 ;
        RECT 1305.580 14.290 1305.840 14.610 ;
        RECT 591.200 13.950 591.460 14.270 ;
        RECT 591.260 2.400 591.400 13.950 ;
        RECT 591.050 -4.800 591.610 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 97.470 -4.800 98.030 0.300 ;
=======
        RECT 1175.850 1700.410 1176.130 1704.000 ;
        RECT 1175.000 1700.270 1176.130 1700.410 ;
        RECT 1175.000 1678.140 1175.140 1700.270 ;
        RECT 1175.850 1700.000 1176.130 1700.270 ;
        RECT 1173.620 1678.000 1175.140 1678.140 ;
        RECT 1173.620 20.245 1173.760 1678.000 ;
        RECT 97.610 19.875 97.890 20.245 ;
        RECT 1173.550 19.875 1173.830 20.245 ;
        RECT 97.680 2.400 97.820 19.875 ;
        RECT 97.470 -4.800 98.030 2.400 ;
      LAYER via2 ;
        RECT 97.610 19.920 97.890 20.200 ;
        RECT 1173.550 19.920 1173.830 20.200 ;
      LAYER met3 ;
        RECT 97.585 20.210 97.915 20.225 ;
        RECT 1173.525 20.210 1173.855 20.225 ;
        RECT 97.585 19.910 1173.855 20.210 ;
        RECT 97.585 19.895 97.915 19.910 ;
        RECT 1173.525 19.895 1173.855 19.910 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 141.290 1687.660 141.610 1687.720 ;
        RECT 1176.290 1687.660 1176.610 1687.720 ;
        RECT 141.290 1687.520 1176.610 1687.660 ;
        RECT 141.290 1687.460 141.610 1687.520 ;
        RECT 1176.290 1687.460 1176.610 1687.520 ;
        RECT 97.590 20.300 97.910 20.360 ;
        RECT 141.290 20.300 141.610 20.360 ;
        RECT 97.590 20.160 141.610 20.300 ;
        RECT 97.590 20.100 97.910 20.160 ;
        RECT 141.290 20.100 141.610 20.160 ;
      LAYER via ;
        RECT 141.320 1687.460 141.580 1687.720 ;
        RECT 1176.320 1687.460 1176.580 1687.720 ;
        RECT 97.620 20.100 97.880 20.360 ;
        RECT 141.320 20.100 141.580 20.360 ;
      LAYER met2 ;
        RECT 1176.310 1700.000 1176.590 1704.000 ;
        RECT 1176.380 1687.750 1176.520 1700.000 ;
        RECT 141.320 1687.430 141.580 1687.750 ;
        RECT 1176.320 1687.430 1176.580 1687.750 ;
        RECT 141.380 20.390 141.520 1687.430 ;
        RECT 97.620 20.070 97.880 20.390 ;
        RECT 141.320 20.070 141.580 20.390 ;
        RECT 97.680 2.400 97.820 20.070 ;
        RECT 97.470 -4.800 98.030 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 0.300 ;
=======
      LAYER met1 ;
        RECT 955.490 1683.920 955.810 1683.980 ;
        RECT 1314.290 1683.920 1314.610 1683.980 ;
        RECT 955.490 1683.780 1314.610 1683.920 ;
        RECT 955.490 1683.720 955.810 1683.780 ;
        RECT 1314.290 1683.720 1314.610 1683.780 ;
        RECT 609.110 27.440 609.430 27.500 ;
        RECT 955.490 27.440 955.810 27.500 ;
        RECT 609.110 27.300 955.810 27.440 ;
        RECT 609.110 27.240 609.430 27.300 ;
        RECT 955.490 27.240 955.810 27.300 ;
      LAYER via ;
        RECT 955.520 1683.720 955.780 1683.980 ;
        RECT 1314.320 1683.720 1314.580 1683.980 ;
        RECT 609.140 27.240 609.400 27.500 ;
        RECT 955.520 27.240 955.780 27.500 ;
      LAYER met2 ;
        RECT 1314.310 1700.000 1314.590 1704.000 ;
        RECT 1314.380 1684.010 1314.520 1700.000 ;
        RECT 955.520 1683.690 955.780 1684.010 ;
        RECT 1314.320 1683.690 1314.580 1684.010 ;
        RECT 955.580 27.530 955.720 1683.690 ;
        RECT 609.140 27.210 609.400 27.530 ;
        RECT 955.520 27.210 955.780 27.530 ;
        RECT 609.200 2.400 609.340 27.210 ;
=======
      LAYER li1 ;
        RECT 1312.985 572.645 1313.155 620.755 ;
        RECT 1312.985 524.365 1313.155 545.275 ;
        RECT 1312.985 386.325 1313.155 493.595 ;
      LAYER mcon ;
        RECT 1312.985 620.585 1313.155 620.755 ;
        RECT 1312.985 545.105 1313.155 545.275 ;
        RECT 1312.985 493.425 1313.155 493.595 ;
      LAYER met1 ;
        RECT 1312.910 1642.440 1313.230 1642.500 ;
        RECT 1314.290 1642.440 1314.610 1642.500 ;
        RECT 1312.910 1642.300 1314.610 1642.440 ;
        RECT 1312.910 1642.240 1313.230 1642.300 ;
        RECT 1314.290 1642.240 1314.610 1642.300 ;
        RECT 1312.910 717.640 1313.230 717.700 ;
        RECT 1313.370 717.640 1313.690 717.700 ;
        RECT 1312.910 717.500 1313.690 717.640 ;
        RECT 1312.910 717.440 1313.230 717.500 ;
        RECT 1313.370 717.440 1313.690 717.500 ;
        RECT 1312.910 620.740 1313.230 620.800 ;
        RECT 1312.715 620.600 1313.230 620.740 ;
        RECT 1312.910 620.540 1313.230 620.600 ;
        RECT 1312.910 572.800 1313.230 572.860 ;
        RECT 1312.715 572.660 1313.230 572.800 ;
        RECT 1312.910 572.600 1313.230 572.660 ;
        RECT 1312.910 545.260 1313.230 545.320 ;
        RECT 1312.715 545.120 1313.230 545.260 ;
        RECT 1312.910 545.060 1313.230 545.120 ;
        RECT 1312.910 524.520 1313.230 524.580 ;
        RECT 1312.715 524.380 1313.230 524.520 ;
        RECT 1312.910 524.320 1313.230 524.380 ;
        RECT 1312.910 493.580 1313.230 493.640 ;
        RECT 1312.715 493.440 1313.230 493.580 ;
        RECT 1312.910 493.380 1313.230 493.440 ;
        RECT 1312.910 386.480 1313.230 386.540 ;
        RECT 1312.715 386.340 1313.230 386.480 ;
        RECT 1312.910 386.280 1313.230 386.340 ;
        RECT 609.110 14.180 609.430 14.240 ;
        RECT 1312.910 14.180 1313.230 14.240 ;
        RECT 609.110 14.040 1313.230 14.180 ;
        RECT 609.110 13.980 609.430 14.040 ;
        RECT 1312.910 13.980 1313.230 14.040 ;
      LAYER via ;
        RECT 1312.940 1642.240 1313.200 1642.500 ;
        RECT 1314.320 1642.240 1314.580 1642.500 ;
        RECT 1312.940 717.440 1313.200 717.700 ;
        RECT 1313.400 717.440 1313.660 717.700 ;
        RECT 1312.940 620.540 1313.200 620.800 ;
        RECT 1312.940 572.600 1313.200 572.860 ;
        RECT 1312.940 545.060 1313.200 545.320 ;
        RECT 1312.940 524.320 1313.200 524.580 ;
        RECT 1312.940 493.380 1313.200 493.640 ;
        RECT 1312.940 386.280 1313.200 386.540 ;
        RECT 609.140 13.980 609.400 14.240 ;
        RECT 1312.940 13.980 1313.200 14.240 ;
      LAYER met2 ;
        RECT 1314.770 1700.410 1315.050 1704.000 ;
        RECT 1314.380 1700.270 1315.050 1700.410 ;
        RECT 1314.380 1642.530 1314.520 1700.270 ;
        RECT 1314.770 1700.000 1315.050 1700.270 ;
        RECT 1312.940 1642.210 1313.200 1642.530 ;
        RECT 1314.320 1642.210 1314.580 1642.530 ;
        RECT 1313.000 737.530 1313.140 1642.210 ;
        RECT 1313.000 737.390 1313.600 737.530 ;
        RECT 1313.460 717.730 1313.600 737.390 ;
        RECT 1312.940 717.410 1313.200 717.730 ;
        RECT 1313.400 717.410 1313.660 717.730 ;
        RECT 1313.000 620.830 1313.140 717.410 ;
        RECT 1312.940 620.510 1313.200 620.830 ;
        RECT 1312.940 572.570 1313.200 572.890 ;
        RECT 1313.000 545.350 1313.140 572.570 ;
        RECT 1312.940 545.030 1313.200 545.350 ;
        RECT 1312.940 524.290 1313.200 524.610 ;
        RECT 1313.000 493.670 1313.140 524.290 ;
        RECT 1312.940 493.350 1313.200 493.670 ;
        RECT 1312.940 386.250 1313.200 386.570 ;
        RECT 1313.000 14.270 1313.140 386.250 ;
        RECT 609.140 13.950 609.400 14.270 ;
        RECT 1312.940 13.950 1313.200 14.270 ;
        RECT 609.200 2.400 609.340 13.950 ;
>>>>>>> re-updated local openlane
        RECT 608.990 -4.800 609.550 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 0.300 ;
=======
      LAYER met1 ;
        RECT 1317.970 14.520 1318.290 14.580 ;
        RECT 632.200 14.380 1318.290 14.520 ;
        RECT 627.050 14.180 627.370 14.240 ;
        RECT 632.200 14.180 632.340 14.380 ;
        RECT 1317.970 14.320 1318.290 14.380 ;
        RECT 627.050 14.040 632.340 14.180 ;
        RECT 627.050 13.980 627.370 14.040 ;
      LAYER via ;
        RECT 627.080 13.980 627.340 14.240 ;
        RECT 1318.000 14.320 1318.260 14.580 ;
      LAYER met2 ;
        RECT 1318.910 1700.410 1319.190 1704.000 ;
        RECT 1318.060 1700.270 1319.190 1700.410 ;
        RECT 1318.060 14.610 1318.200 1700.270 ;
        RECT 1318.910 1700.000 1319.190 1700.270 ;
        RECT 1318.000 14.290 1318.260 14.610 ;
        RECT 627.080 13.950 627.340 14.270 ;
        RECT 627.140 2.400 627.280 13.950 ;
=======
      LAYER li1 ;
        RECT 627.585 1642.285 627.755 1685.975 ;
        RECT 628.045 1685.125 628.215 1685.975 ;
        RECT 675.885 1685.125 676.055 1685.975 ;
        RECT 724.645 1685.125 724.815 1685.975 ;
        RECT 772.485 1685.125 772.655 1685.975 ;
        RECT 821.245 1685.125 821.415 1685.975 ;
        RECT 869.085 1685.125 869.255 1685.975 ;
        RECT 917.845 1685.125 918.015 1685.975 ;
        RECT 965.685 1685.125 965.855 1685.975 ;
        RECT 1014.445 1685.125 1014.615 1685.975 ;
        RECT 1062.285 1685.125 1062.455 1685.975 ;
        RECT 1104.145 1685.125 1104.315 1685.975 ;
        RECT 1151.985 1685.125 1152.155 1685.975 ;
        RECT 1200.745 1685.125 1200.915 1686.315 ;
        RECT 1272.965 1684.785 1273.135 1686.315 ;
      LAYER mcon ;
        RECT 1200.745 1686.145 1200.915 1686.315 ;
        RECT 627.585 1685.805 627.755 1685.975 ;
        RECT 628.045 1685.805 628.215 1685.975 ;
        RECT 675.885 1685.805 676.055 1685.975 ;
        RECT 724.645 1685.805 724.815 1685.975 ;
        RECT 772.485 1685.805 772.655 1685.975 ;
        RECT 821.245 1685.805 821.415 1685.975 ;
        RECT 869.085 1685.805 869.255 1685.975 ;
        RECT 917.845 1685.805 918.015 1685.975 ;
        RECT 965.685 1685.805 965.855 1685.975 ;
        RECT 1014.445 1685.805 1014.615 1685.975 ;
        RECT 1062.285 1685.805 1062.455 1685.975 ;
        RECT 1104.145 1685.805 1104.315 1685.975 ;
        RECT 1151.985 1685.805 1152.155 1685.975 ;
        RECT 1272.965 1686.145 1273.135 1686.315 ;
      LAYER met1 ;
        RECT 1319.810 1686.640 1320.130 1686.700 ;
        RECT 1312.080 1686.500 1320.130 1686.640 ;
        RECT 676.270 1686.300 676.590 1686.360 ;
        RECT 772.870 1686.300 773.190 1686.360 ;
        RECT 869.470 1686.300 869.790 1686.360 ;
        RECT 966.070 1686.300 966.390 1686.360 ;
        RECT 1062.670 1686.300 1062.990 1686.360 ;
        RECT 1200.685 1686.300 1200.975 1686.345 ;
        RECT 627.600 1686.160 628.200 1686.300 ;
        RECT 627.600 1686.005 627.740 1686.160 ;
        RECT 628.060 1686.005 628.200 1686.160 ;
        RECT 675.900 1686.160 676.590 1686.300 ;
        RECT 675.900 1686.005 676.040 1686.160 ;
        RECT 676.270 1686.100 676.590 1686.160 ;
        RECT 724.200 1686.160 724.800 1686.300 ;
        RECT 627.525 1685.775 627.815 1686.005 ;
        RECT 627.985 1685.775 628.275 1686.005 ;
        RECT 675.825 1685.775 676.115 1686.005 ;
        RECT 676.730 1685.960 677.050 1686.020 ;
        RECT 724.200 1685.960 724.340 1686.160 ;
        RECT 724.660 1686.005 724.800 1686.160 ;
        RECT 772.500 1686.160 773.190 1686.300 ;
        RECT 772.500 1686.005 772.640 1686.160 ;
        RECT 772.870 1686.100 773.190 1686.160 ;
        RECT 820.800 1686.160 821.400 1686.300 ;
        RECT 676.730 1685.820 724.340 1685.960 ;
        RECT 676.730 1685.760 677.050 1685.820 ;
        RECT 724.585 1685.775 724.875 1686.005 ;
        RECT 772.425 1685.775 772.715 1686.005 ;
        RECT 773.330 1685.960 773.650 1686.020 ;
        RECT 820.800 1685.960 820.940 1686.160 ;
        RECT 821.260 1686.005 821.400 1686.160 ;
        RECT 869.100 1686.160 869.790 1686.300 ;
        RECT 869.100 1686.005 869.240 1686.160 ;
        RECT 869.470 1686.100 869.790 1686.160 ;
        RECT 917.400 1686.160 918.000 1686.300 ;
        RECT 773.330 1685.820 820.940 1685.960 ;
        RECT 773.330 1685.760 773.650 1685.820 ;
        RECT 821.185 1685.775 821.475 1686.005 ;
        RECT 869.025 1685.775 869.315 1686.005 ;
        RECT 869.930 1685.960 870.250 1686.020 ;
        RECT 917.400 1685.960 917.540 1686.160 ;
        RECT 917.860 1686.005 918.000 1686.160 ;
        RECT 965.700 1686.160 966.390 1686.300 ;
        RECT 965.700 1686.005 965.840 1686.160 ;
        RECT 966.070 1686.100 966.390 1686.160 ;
        RECT 1014.000 1686.160 1014.600 1686.300 ;
        RECT 869.930 1685.820 917.540 1685.960 ;
        RECT 869.930 1685.760 870.250 1685.820 ;
        RECT 917.785 1685.775 918.075 1686.005 ;
        RECT 965.625 1685.775 965.915 1686.005 ;
        RECT 966.530 1685.960 966.850 1686.020 ;
        RECT 1014.000 1685.960 1014.140 1686.160 ;
        RECT 1014.460 1686.005 1014.600 1686.160 ;
        RECT 1062.300 1686.160 1062.990 1686.300 ;
        RECT 1062.300 1686.005 1062.440 1686.160 ;
        RECT 1062.670 1686.100 1062.990 1686.160 ;
        RECT 1152.000 1686.160 1200.975 1686.300 ;
        RECT 966.530 1685.820 1014.140 1685.960 ;
        RECT 966.530 1685.760 966.850 1685.820 ;
        RECT 1014.385 1685.775 1014.675 1686.005 ;
        RECT 1062.225 1685.775 1062.515 1686.005 ;
        RECT 1063.130 1685.960 1063.450 1686.020 ;
        RECT 1152.000 1686.005 1152.140 1686.160 ;
        RECT 1200.685 1686.115 1200.975 1686.160 ;
        RECT 1272.905 1686.300 1273.195 1686.345 ;
        RECT 1312.080 1686.300 1312.220 1686.500 ;
        RECT 1319.810 1686.440 1320.130 1686.500 ;
        RECT 1272.905 1686.160 1312.220 1686.300 ;
        RECT 1272.905 1686.115 1273.195 1686.160 ;
        RECT 1104.085 1685.960 1104.375 1686.005 ;
        RECT 1063.130 1685.820 1104.375 1685.960 ;
        RECT 1063.130 1685.760 1063.450 1685.820 ;
        RECT 1104.085 1685.775 1104.375 1685.820 ;
        RECT 1151.925 1685.775 1152.215 1686.005 ;
        RECT 627.985 1685.280 628.275 1685.325 ;
        RECT 675.825 1685.280 676.115 1685.325 ;
        RECT 627.985 1685.140 676.115 1685.280 ;
        RECT 627.985 1685.095 628.275 1685.140 ;
        RECT 675.825 1685.095 676.115 1685.140 ;
        RECT 724.585 1685.280 724.875 1685.325 ;
        RECT 772.425 1685.280 772.715 1685.325 ;
        RECT 724.585 1685.140 772.715 1685.280 ;
        RECT 724.585 1685.095 724.875 1685.140 ;
        RECT 772.425 1685.095 772.715 1685.140 ;
        RECT 821.185 1685.280 821.475 1685.325 ;
        RECT 869.025 1685.280 869.315 1685.325 ;
        RECT 821.185 1685.140 869.315 1685.280 ;
        RECT 821.185 1685.095 821.475 1685.140 ;
        RECT 869.025 1685.095 869.315 1685.140 ;
        RECT 917.785 1685.280 918.075 1685.325 ;
        RECT 965.625 1685.280 965.915 1685.325 ;
        RECT 917.785 1685.140 965.915 1685.280 ;
        RECT 917.785 1685.095 918.075 1685.140 ;
        RECT 965.625 1685.095 965.915 1685.140 ;
        RECT 1014.385 1685.280 1014.675 1685.325 ;
        RECT 1062.225 1685.280 1062.515 1685.325 ;
        RECT 1014.385 1685.140 1062.515 1685.280 ;
        RECT 1014.385 1685.095 1014.675 1685.140 ;
        RECT 1062.225 1685.095 1062.515 1685.140 ;
        RECT 1104.085 1685.280 1104.375 1685.325 ;
        RECT 1151.925 1685.280 1152.215 1685.325 ;
        RECT 1104.085 1685.140 1152.215 1685.280 ;
        RECT 1104.085 1685.095 1104.375 1685.140 ;
        RECT 1151.925 1685.095 1152.215 1685.140 ;
        RECT 1200.685 1685.280 1200.975 1685.325 ;
        RECT 1200.685 1685.140 1249.200 1685.280 ;
        RECT 1200.685 1685.095 1200.975 1685.140 ;
        RECT 1249.060 1684.940 1249.200 1685.140 ;
        RECT 1272.905 1684.940 1273.195 1684.985 ;
        RECT 1249.060 1684.800 1273.195 1684.940 ;
        RECT 1272.905 1684.755 1273.195 1684.800 ;
        RECT 627.510 1642.440 627.830 1642.500 ;
        RECT 627.315 1642.300 627.830 1642.440 ;
        RECT 627.510 1642.240 627.830 1642.300 ;
      LAYER via ;
        RECT 676.300 1686.100 676.560 1686.360 ;
        RECT 676.760 1685.760 677.020 1686.020 ;
        RECT 772.900 1686.100 773.160 1686.360 ;
        RECT 773.360 1685.760 773.620 1686.020 ;
        RECT 869.500 1686.100 869.760 1686.360 ;
        RECT 869.960 1685.760 870.220 1686.020 ;
        RECT 966.100 1686.100 966.360 1686.360 ;
        RECT 966.560 1685.760 966.820 1686.020 ;
        RECT 1062.700 1686.100 1062.960 1686.360 ;
        RECT 1063.160 1685.760 1063.420 1686.020 ;
        RECT 1319.840 1686.440 1320.100 1686.700 ;
        RECT 627.540 1642.240 627.800 1642.500 ;
      LAYER met2 ;
        RECT 1319.830 1700.000 1320.110 1704.000 ;
        RECT 676.360 1686.670 676.960 1686.810 ;
        RECT 676.360 1686.390 676.500 1686.670 ;
        RECT 676.300 1686.070 676.560 1686.390 ;
        RECT 676.820 1686.050 676.960 1686.670 ;
        RECT 772.960 1686.670 773.560 1686.810 ;
        RECT 772.960 1686.390 773.100 1686.670 ;
        RECT 772.900 1686.070 773.160 1686.390 ;
        RECT 773.420 1686.050 773.560 1686.670 ;
        RECT 869.560 1686.670 870.160 1686.810 ;
        RECT 869.560 1686.390 869.700 1686.670 ;
        RECT 869.500 1686.070 869.760 1686.390 ;
        RECT 870.020 1686.050 870.160 1686.670 ;
        RECT 966.160 1686.670 966.760 1686.810 ;
        RECT 966.160 1686.390 966.300 1686.670 ;
        RECT 966.100 1686.070 966.360 1686.390 ;
        RECT 966.620 1686.050 966.760 1686.670 ;
        RECT 1062.760 1686.670 1063.360 1686.810 ;
        RECT 1319.900 1686.730 1320.040 1700.000 ;
        RECT 1062.760 1686.390 1062.900 1686.670 ;
        RECT 1062.700 1686.070 1062.960 1686.390 ;
        RECT 1063.220 1686.050 1063.360 1686.670 ;
        RECT 1319.840 1686.410 1320.100 1686.730 ;
        RECT 676.760 1685.730 677.020 1686.050 ;
        RECT 773.360 1685.730 773.620 1686.050 ;
        RECT 869.960 1685.730 870.220 1686.050 ;
        RECT 966.560 1685.730 966.820 1686.050 ;
        RECT 1063.160 1685.730 1063.420 1686.050 ;
        RECT 627.540 1642.210 627.800 1642.530 ;
        RECT 627.600 17.410 627.740 1642.210 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
>>>>>>> re-updated local openlane
        RECT 626.930 -4.800 627.490 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 0.300 ;
=======
      LAYER li1 ;
        RECT 227.845 16.405 228.015 17.935 ;
        RECT 275.685 16.405 275.855 17.935 ;
        RECT 276.605 16.065 276.775 17.935 ;
        RECT 323.525 16.065 323.695 17.935 ;
        RECT 373.205 15.045 373.375 17.935 ;
        RECT 420.125 15.045 420.295 17.935 ;
        RECT 469.805 14.705 469.975 17.935 ;
        RECT 516.725 14.705 516.895 17.935 ;
        RECT 566.405 14.365 566.575 17.935 ;
        RECT 613.325 14.025 613.495 17.935 ;
        RECT 663.005 17.765 663.175 21.675 ;
        RECT 709.465 17.935 709.635 21.675 ;
        RECT 709.465 17.765 710.095 17.935 ;
        RECT 856.205 17.765 856.375 21.335 ;
        RECT 903.125 17.765 903.295 21.335 ;
        RECT 952.805 17.765 952.975 21.335 ;
        RECT 999.725 17.765 999.895 21.335 ;
        RECT 1049.405 17.765 1049.575 21.335 ;
        RECT 1096.325 17.765 1096.495 21.335 ;
      LAYER mcon ;
        RECT 663.005 21.505 663.175 21.675 ;
        RECT 227.845 17.765 228.015 17.935 ;
        RECT 275.685 17.765 275.855 17.935 ;
        RECT 276.605 17.765 276.775 17.935 ;
        RECT 323.525 17.765 323.695 17.935 ;
        RECT 373.205 17.765 373.375 17.935 ;
        RECT 420.125 17.765 420.295 17.935 ;
        RECT 469.805 17.765 469.975 17.935 ;
        RECT 516.725 17.765 516.895 17.935 ;
        RECT 566.405 17.765 566.575 17.935 ;
        RECT 613.325 17.765 613.495 17.935 ;
        RECT 709.465 21.505 709.635 21.675 ;
        RECT 856.205 21.165 856.375 21.335 ;
        RECT 709.925 17.765 710.095 17.935 ;
        RECT 903.125 21.165 903.295 21.335 ;
        RECT 952.805 21.165 952.975 21.335 ;
        RECT 999.725 21.165 999.895 21.335 ;
        RECT 1049.405 21.165 1049.575 21.335 ;
        RECT 1096.325 21.165 1096.495 21.335 ;
      LAYER met1 ;
        RECT 662.945 21.660 663.235 21.705 ;
        RECT 709.405 21.660 709.695 21.705 ;
        RECT 662.945 21.520 709.695 21.660 ;
        RECT 662.945 21.475 663.235 21.520 ;
        RECT 709.405 21.475 709.695 21.520 ;
        RECT 856.145 21.320 856.435 21.365 ;
        RECT 903.065 21.320 903.355 21.365 ;
        RECT 856.145 21.180 903.355 21.320 ;
        RECT 856.145 21.135 856.435 21.180 ;
        RECT 903.065 21.135 903.355 21.180 ;
        RECT 952.745 21.320 953.035 21.365 ;
        RECT 999.665 21.320 999.955 21.365 ;
        RECT 952.745 21.180 999.955 21.320 ;
        RECT 952.745 21.135 953.035 21.180 ;
        RECT 999.665 21.135 999.955 21.180 ;
        RECT 1049.345 21.320 1049.635 21.365 ;
        RECT 1096.265 21.320 1096.555 21.365 ;
        RECT 1049.345 21.180 1096.555 21.320 ;
        RECT 1049.345 21.135 1049.635 21.180 ;
        RECT 1096.265 21.135 1096.555 21.180 ;
        RECT 121.510 18.600 121.830 18.660 ;
        RECT 121.510 18.460 139.220 18.600 ;
        RECT 121.510 18.400 121.830 18.460 ;
        RECT 139.080 17.920 139.220 18.460 ;
        RECT 227.785 17.920 228.075 17.965 ;
        RECT 139.080 17.780 228.075 17.920 ;
        RECT 227.785 17.735 228.075 17.780 ;
        RECT 275.625 17.920 275.915 17.965 ;
        RECT 276.545 17.920 276.835 17.965 ;
        RECT 275.625 17.780 276.835 17.920 ;
        RECT 275.625 17.735 275.915 17.780 ;
        RECT 276.545 17.735 276.835 17.780 ;
        RECT 323.465 17.920 323.755 17.965 ;
        RECT 373.145 17.920 373.435 17.965 ;
        RECT 323.465 17.780 373.435 17.920 ;
        RECT 323.465 17.735 323.755 17.780 ;
        RECT 373.145 17.735 373.435 17.780 ;
        RECT 420.065 17.920 420.355 17.965 ;
        RECT 469.745 17.920 470.035 17.965 ;
        RECT 420.065 17.780 470.035 17.920 ;
        RECT 420.065 17.735 420.355 17.780 ;
        RECT 469.745 17.735 470.035 17.780 ;
        RECT 516.665 17.920 516.955 17.965 ;
        RECT 566.345 17.920 566.635 17.965 ;
        RECT 516.665 17.780 566.635 17.920 ;
        RECT 516.665 17.735 516.955 17.780 ;
        RECT 566.345 17.735 566.635 17.780 ;
        RECT 613.265 17.920 613.555 17.965 ;
        RECT 662.945 17.920 663.235 17.965 ;
        RECT 613.265 17.780 663.235 17.920 ;
        RECT 613.265 17.735 613.555 17.780 ;
        RECT 662.945 17.735 663.235 17.780 ;
        RECT 709.865 17.920 710.155 17.965 ;
        RECT 759.530 17.920 759.850 17.980 ;
        RECT 709.865 17.780 759.850 17.920 ;
        RECT 709.865 17.735 710.155 17.780 ;
        RECT 759.530 17.720 759.850 17.780 ;
        RECT 806.450 17.920 806.770 17.980 ;
        RECT 856.145 17.920 856.435 17.965 ;
        RECT 806.450 17.780 856.435 17.920 ;
        RECT 806.450 17.720 806.770 17.780 ;
        RECT 856.145 17.735 856.435 17.780 ;
        RECT 903.065 17.920 903.355 17.965 ;
        RECT 952.745 17.920 953.035 17.965 ;
        RECT 903.065 17.780 953.035 17.920 ;
        RECT 903.065 17.735 903.355 17.780 ;
        RECT 952.745 17.735 953.035 17.780 ;
        RECT 999.665 17.920 999.955 17.965 ;
        RECT 1049.345 17.920 1049.635 17.965 ;
        RECT 999.665 17.780 1049.635 17.920 ;
        RECT 999.665 17.735 999.955 17.780 ;
        RECT 1049.345 17.735 1049.635 17.780 ;
        RECT 1096.265 17.920 1096.555 17.965 ;
        RECT 1180.430 17.920 1180.750 17.980 ;
        RECT 1096.265 17.780 1180.750 17.920 ;
        RECT 1096.265 17.735 1096.555 17.780 ;
        RECT 1180.430 17.720 1180.750 17.780 ;
        RECT 227.785 16.560 228.075 16.605 ;
        RECT 275.625 16.560 275.915 16.605 ;
        RECT 227.785 16.420 275.915 16.560 ;
        RECT 227.785 16.375 228.075 16.420 ;
        RECT 275.625 16.375 275.915 16.420 ;
        RECT 276.545 16.220 276.835 16.265 ;
        RECT 323.465 16.220 323.755 16.265 ;
        RECT 276.545 16.080 323.755 16.220 ;
        RECT 276.545 16.035 276.835 16.080 ;
        RECT 323.465 16.035 323.755 16.080 ;
        RECT 373.145 15.200 373.435 15.245 ;
        RECT 420.065 15.200 420.355 15.245 ;
        RECT 373.145 15.060 420.355 15.200 ;
        RECT 373.145 15.015 373.435 15.060 ;
        RECT 420.065 15.015 420.355 15.060 ;
        RECT 469.745 14.860 470.035 14.905 ;
        RECT 516.665 14.860 516.955 14.905 ;
        RECT 469.745 14.720 516.955 14.860 ;
        RECT 469.745 14.675 470.035 14.720 ;
        RECT 516.665 14.675 516.955 14.720 ;
        RECT 566.345 14.520 566.635 14.565 ;
        RECT 566.345 14.380 590.940 14.520 ;
        RECT 566.345 14.335 566.635 14.380 ;
        RECT 590.800 13.840 590.940 14.380 ;
        RECT 613.265 14.180 613.555 14.225 ;
        RECT 601.380 14.040 613.555 14.180 ;
        RECT 601.380 13.840 601.520 14.040 ;
        RECT 613.265 13.995 613.555 14.040 ;
        RECT 590.800 13.700 601.520 13.840 ;
      LAYER via ;
        RECT 121.540 18.400 121.800 18.660 ;
        RECT 759.560 17.720 759.820 17.980 ;
        RECT 806.480 17.720 806.740 17.980 ;
        RECT 1180.460 17.720 1180.720 17.980 ;
      LAYER met2 ;
        RECT 1182.290 1700.410 1182.570 1704.000 ;
        RECT 1181.440 1700.270 1182.570 1700.410 ;
        RECT 1181.440 1677.290 1181.580 1700.270 ;
        RECT 1182.290 1700.000 1182.570 1700.270 ;
        RECT 1180.520 1677.150 1181.580 1677.290 ;
        RECT 121.540 18.370 121.800 18.690 ;
        RECT 121.600 2.400 121.740 18.370 ;
        RECT 1180.520 18.010 1180.660 1677.150 ;
        RECT 759.560 17.690 759.820 18.010 ;
        RECT 806.480 17.690 806.740 18.010 ;
        RECT 1180.460 17.690 1180.720 18.010 ;
        RECT 759.620 16.165 759.760 17.690 ;
        RECT 806.540 16.165 806.680 17.690 ;
        RECT 759.550 15.795 759.830 16.165 ;
        RECT 806.470 15.795 806.750 16.165 ;
=======
      LAYER met1 ;
        RECT 1179.970 1679.160 1180.290 1679.220 ;
        RECT 1181.350 1679.160 1181.670 1679.220 ;
        RECT 1179.970 1679.020 1181.670 1679.160 ;
        RECT 1179.970 1678.960 1180.290 1679.020 ;
        RECT 1181.350 1678.960 1181.670 1679.020 ;
        RECT 1179.970 48.520 1180.290 48.580 ;
        RECT 1180.890 48.520 1181.210 48.580 ;
        RECT 1179.970 48.380 1181.210 48.520 ;
        RECT 1179.970 48.320 1180.290 48.380 ;
        RECT 1180.890 48.320 1181.210 48.380 ;
      LAYER via ;
        RECT 1180.000 1678.960 1180.260 1679.220 ;
        RECT 1181.380 1678.960 1181.640 1679.220 ;
        RECT 1180.000 48.320 1180.260 48.580 ;
        RECT 1180.920 48.320 1181.180 48.580 ;
      LAYER met2 ;
        RECT 1182.750 1700.410 1183.030 1704.000 ;
        RECT 1181.440 1700.270 1183.030 1700.410 ;
        RECT 1181.440 1679.250 1181.580 1700.270 ;
        RECT 1182.750 1700.000 1183.030 1700.270 ;
        RECT 1180.000 1678.930 1180.260 1679.250 ;
        RECT 1181.380 1678.930 1181.640 1679.250 ;
        RECT 1180.060 48.610 1180.200 1678.930 ;
        RECT 1180.000 48.290 1180.260 48.610 ;
        RECT 1180.920 48.290 1181.180 48.610 ;
        RECT 1180.980 18.885 1181.120 48.290 ;
        RECT 121.530 18.515 121.810 18.885 ;
        RECT 1180.910 18.515 1181.190 18.885 ;
        RECT 121.600 2.400 121.740 18.515 ;
>>>>>>> re-updated local openlane
        RECT 121.390 -4.800 121.950 2.400 ;
      LAYER via2 ;
        RECT 121.530 18.560 121.810 18.840 ;
        RECT 1180.910 18.560 1181.190 18.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 759.525 16.130 759.855 16.145 ;
        RECT 806.445 16.130 806.775 16.145 ;
        RECT 759.525 15.830 806.775 16.130 ;
        RECT 759.525 15.815 759.855 15.830 ;
        RECT 806.445 15.815 806.775 15.830 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 121.505 18.850 121.835 18.865 ;
        RECT 1180.885 18.850 1181.215 18.865 ;
        RECT 121.505 18.550 1181.215 18.850 ;
        RECT 121.505 18.535 121.835 18.550 ;
        RECT 1180.885 18.535 1181.215 18.550 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 0.300 ;
=======
      LAYER li1 ;
        RECT 276.605 18.445 276.775 20.655 ;
        RECT 323.525 18.445 323.695 20.655 ;
        RECT 373.205 18.445 373.835 18.615 ;
        RECT 373.665 16.405 373.835 18.445 ;
        RECT 419.665 18.445 420.295 18.615 ;
        RECT 469.805 18.445 470.435 18.615 ;
        RECT 419.665 16.405 419.835 18.445 ;
        RECT 470.265 14.365 470.435 18.445 ;
        RECT 516.265 18.445 516.895 18.615 ;
        RECT 566.405 18.445 566.575 20.995 ;
        RECT 613.325 18.445 613.495 20.995 ;
        RECT 759.605 18.445 759.775 21.675 ;
        RECT 806.525 18.445 806.695 21.675 ;
        RECT 1049.865 18.445 1050.035 21.675 ;
        RECT 516.265 14.365 516.435 18.445 ;
      LAYER mcon ;
        RECT 759.605 21.505 759.775 21.675 ;
        RECT 566.405 20.825 566.575 20.995 ;
        RECT 276.605 20.485 276.775 20.655 ;
        RECT 323.525 20.485 323.695 20.655 ;
        RECT 420.125 18.445 420.295 18.615 ;
        RECT 516.725 18.445 516.895 18.615 ;
        RECT 613.325 20.825 613.495 20.995 ;
        RECT 806.525 21.505 806.695 21.675 ;
        RECT 1049.865 21.505 1050.035 21.675 ;
      LAYER met1 ;
        RECT 759.545 21.660 759.835 21.705 ;
        RECT 806.465 21.660 806.755 21.705 ;
        RECT 759.545 21.520 806.755 21.660 ;
        RECT 759.545 21.475 759.835 21.520 ;
        RECT 806.465 21.475 806.755 21.520 ;
        RECT 1049.805 21.660 1050.095 21.705 ;
        RECT 1095.790 21.660 1096.110 21.720 ;
        RECT 1049.805 21.520 1096.110 21.660 ;
        RECT 1049.805 21.475 1050.095 21.520 ;
        RECT 1095.790 21.460 1096.110 21.520 ;
        RECT 566.345 20.980 566.635 21.025 ;
        RECT 613.265 20.980 613.555 21.025 ;
        RECT 566.345 20.840 613.555 20.980 ;
        RECT 566.345 20.795 566.635 20.840 ;
        RECT 613.265 20.795 613.555 20.840 ;
        RECT 276.545 20.640 276.835 20.685 ;
        RECT 323.465 20.640 323.755 20.685 ;
        RECT 276.545 20.500 323.755 20.640 ;
        RECT 276.545 20.455 276.835 20.500 ;
        RECT 323.465 20.455 323.755 20.500 ;
        RECT 145.430 18.600 145.750 18.660 ;
        RECT 276.545 18.600 276.835 18.645 ;
        RECT 145.430 18.460 276.835 18.600 ;
        RECT 145.430 18.400 145.750 18.460 ;
        RECT 276.545 18.415 276.835 18.460 ;
        RECT 323.465 18.600 323.755 18.645 ;
        RECT 373.145 18.600 373.435 18.645 ;
        RECT 323.465 18.460 373.435 18.600 ;
        RECT 323.465 18.415 323.755 18.460 ;
        RECT 373.145 18.415 373.435 18.460 ;
        RECT 420.065 18.600 420.355 18.645 ;
        RECT 469.745 18.600 470.035 18.645 ;
        RECT 420.065 18.460 470.035 18.600 ;
        RECT 420.065 18.415 420.355 18.460 ;
        RECT 469.745 18.415 470.035 18.460 ;
        RECT 516.665 18.600 516.955 18.645 ;
        RECT 566.345 18.600 566.635 18.645 ;
        RECT 516.665 18.460 566.635 18.600 ;
        RECT 516.665 18.415 516.955 18.460 ;
        RECT 566.345 18.415 566.635 18.460 ;
        RECT 613.265 18.600 613.555 18.645 ;
        RECT 663.390 18.600 663.710 18.660 ;
        RECT 613.265 18.460 663.710 18.600 ;
        RECT 613.265 18.415 613.555 18.460 ;
        RECT 663.390 18.400 663.710 18.460 ;
        RECT 709.390 18.600 709.710 18.660 ;
        RECT 759.545 18.600 759.835 18.645 ;
        RECT 709.390 18.460 759.835 18.600 ;
        RECT 709.390 18.400 709.710 18.460 ;
        RECT 759.545 18.415 759.835 18.460 ;
        RECT 806.465 18.600 806.755 18.645 ;
        RECT 856.130 18.600 856.450 18.660 ;
        RECT 806.465 18.460 856.450 18.600 ;
        RECT 806.465 18.415 806.755 18.460 ;
        RECT 856.130 18.400 856.450 18.460 ;
        RECT 903.050 18.600 903.370 18.660 ;
        RECT 952.730 18.600 953.050 18.660 ;
        RECT 903.050 18.460 953.050 18.600 ;
        RECT 903.050 18.400 903.370 18.460 ;
        RECT 952.730 18.400 953.050 18.460 ;
        RECT 999.650 18.600 999.970 18.660 ;
        RECT 1049.805 18.600 1050.095 18.645 ;
        RECT 999.650 18.460 1050.095 18.600 ;
        RECT 999.650 18.400 999.970 18.460 ;
        RECT 1049.805 18.415 1050.095 18.460 ;
        RECT 1096.250 18.600 1096.570 18.660 ;
        RECT 1188.710 18.600 1189.030 18.660 ;
        RECT 1096.250 18.460 1189.030 18.600 ;
        RECT 1096.250 18.400 1096.570 18.460 ;
        RECT 1188.710 18.400 1189.030 18.460 ;
        RECT 373.605 16.560 373.895 16.605 ;
        RECT 419.605 16.560 419.895 16.605 ;
        RECT 373.605 16.420 419.895 16.560 ;
        RECT 373.605 16.375 373.895 16.420 ;
        RECT 419.605 16.375 419.895 16.420 ;
        RECT 470.205 14.520 470.495 14.565 ;
        RECT 516.205 14.520 516.495 14.565 ;
        RECT 470.205 14.380 516.495 14.520 ;
        RECT 470.205 14.335 470.495 14.380 ;
        RECT 516.205 14.335 516.495 14.380 ;
      LAYER via ;
        RECT 1095.820 21.460 1096.080 21.720 ;
        RECT 145.460 18.400 145.720 18.660 ;
        RECT 663.420 18.400 663.680 18.660 ;
        RECT 709.420 18.400 709.680 18.660 ;
        RECT 856.160 18.400 856.420 18.660 ;
        RECT 903.080 18.400 903.340 18.660 ;
        RECT 952.760 18.400 953.020 18.660 ;
        RECT 999.680 18.400 999.940 18.660 ;
        RECT 1096.280 18.400 1096.540 18.660 ;
        RECT 1188.740 18.400 1189.000 18.660 ;
      LAYER met2 ;
        RECT 1188.730 1700.000 1189.010 1704.000 ;
        RECT 1095.820 21.490 1096.080 21.750 ;
        RECT 1095.820 21.430 1096.480 21.490 ;
        RECT 1095.880 21.350 1096.480 21.430 ;
        RECT 663.410 20.555 663.690 20.925 ;
        RECT 709.410 20.555 709.690 20.925 ;
        RECT 856.150 20.555 856.430 20.925 ;
        RECT 903.070 20.555 903.350 20.925 ;
        RECT 952.750 20.555 953.030 20.925 ;
        RECT 999.670 20.555 999.950 20.925 ;
        RECT 663.480 18.690 663.620 20.555 ;
        RECT 709.480 18.690 709.620 20.555 ;
        RECT 856.220 18.690 856.360 20.555 ;
        RECT 903.140 18.690 903.280 20.555 ;
        RECT 952.820 18.690 952.960 20.555 ;
        RECT 999.740 18.690 999.880 20.555 ;
        RECT 1096.340 18.690 1096.480 21.350 ;
        RECT 1188.800 18.690 1188.940 1700.000 ;
        RECT 145.460 18.370 145.720 18.690 ;
        RECT 663.420 18.370 663.680 18.690 ;
        RECT 709.420 18.370 709.680 18.690 ;
        RECT 856.160 18.370 856.420 18.690 ;
        RECT 903.080 18.370 903.340 18.690 ;
        RECT 952.760 18.370 953.020 18.690 ;
        RECT 999.680 18.370 999.940 18.690 ;
        RECT 1096.280 18.370 1096.540 18.690 ;
        RECT 1188.740 18.370 1189.000 18.690 ;
        RECT 145.520 2.400 145.660 18.370 ;
        RECT 145.310 -4.800 145.870 2.400 ;
      LAYER via2 ;
        RECT 663.410 20.600 663.690 20.880 ;
        RECT 709.410 20.600 709.690 20.880 ;
        RECT 856.150 20.600 856.430 20.880 ;
        RECT 903.070 20.600 903.350 20.880 ;
        RECT 952.750 20.600 953.030 20.880 ;
        RECT 999.670 20.600 999.950 20.880 ;
      LAYER met3 ;
        RECT 663.385 20.890 663.715 20.905 ;
        RECT 709.385 20.890 709.715 20.905 ;
        RECT 663.385 20.590 709.715 20.890 ;
        RECT 663.385 20.575 663.715 20.590 ;
        RECT 709.385 20.575 709.715 20.590 ;
        RECT 856.125 20.890 856.455 20.905 ;
        RECT 903.045 20.890 903.375 20.905 ;
        RECT 856.125 20.590 903.375 20.890 ;
        RECT 856.125 20.575 856.455 20.590 ;
        RECT 903.045 20.575 903.375 20.590 ;
        RECT 952.725 20.890 953.055 20.905 ;
        RECT 999.645 20.890 999.975 20.905 ;
        RECT 952.725 20.590 999.975 20.890 ;
        RECT 952.725 20.575 953.055 20.590 ;
        RECT 999.645 20.575 999.975 20.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
      LAYER met1 ;
        RECT 175.790 1688.340 176.110 1688.400 ;
        RECT 175.790 1688.200 1165.480 1688.340 ;
        RECT 175.790 1688.140 176.110 1688.200 ;
        RECT 1165.340 1688.000 1165.480 1688.200 ;
        RECT 1189.170 1688.000 1189.490 1688.060 ;
        RECT 1165.340 1687.860 1189.490 1688.000 ;
        RECT 1189.170 1687.800 1189.490 1687.860 ;
        RECT 145.430 17.920 145.750 17.980 ;
        RECT 175.790 17.920 176.110 17.980 ;
        RECT 145.430 17.780 176.110 17.920 ;
        RECT 145.430 17.720 145.750 17.780 ;
        RECT 175.790 17.720 176.110 17.780 ;
      LAYER via ;
        RECT 175.820 1688.140 176.080 1688.400 ;
        RECT 1189.200 1687.800 1189.460 1688.060 ;
        RECT 145.460 17.720 145.720 17.980 ;
        RECT 175.820 17.720 176.080 17.980 ;
      LAYER met2 ;
        RECT 1189.190 1700.000 1189.470 1704.000 ;
        RECT 175.820 1688.110 176.080 1688.430 ;
        RECT 175.880 18.010 176.020 1688.110 ;
        RECT 1189.260 1688.090 1189.400 1700.000 ;
        RECT 1189.200 1687.770 1189.460 1688.090 ;
        RECT 145.460 17.690 145.720 18.010 ;
        RECT 175.820 17.690 176.080 18.010 ;
        RECT 145.520 2.400 145.660 17.690 ;
        RECT 145.310 -4.800 145.870 2.400 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 0.300 ;
=======
      LAYER met1 ;
        RECT 163.370 14.180 163.690 14.240 ;
        RECT 165.210 14.180 165.530 14.240 ;
        RECT 163.370 14.040 165.530 14.180 ;
        RECT 163.370 13.980 163.690 14.040 ;
        RECT 165.210 13.980 165.530 14.040 ;
      LAYER via ;
        RECT 163.400 13.980 163.660 14.240 ;
        RECT 165.240 13.980 165.500 14.240 ;
=======
>>>>>>> re-updated local openlane
      LAYER met2 ;
        RECT 1193.790 1700.000 1194.070 1704.000 ;
        RECT 1193.860 20.245 1194.000 1700.000 ;
        RECT 163.390 19.875 163.670 20.245 ;
        RECT 1193.790 19.875 1194.070 20.245 ;
        RECT 163.460 2.400 163.600 19.875 ;
        RECT 163.250 -4.800 163.810 2.400 ;
      LAYER via2 ;
        RECT 163.390 19.920 163.670 20.200 ;
        RECT 1193.790 19.920 1194.070 20.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 165.205 1689.610 165.535 1689.625 ;
        RECT 1193.765 1689.610 1194.095 1689.625 ;
        RECT 165.205 1689.310 1194.095 1689.610 ;
        RECT 165.205 1689.295 165.535 1689.310 ;
        RECT 1193.765 1689.295 1194.095 1689.310 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 163.365 20.210 163.695 20.225 ;
        RECT 1193.765 20.210 1194.095 20.225 ;
        RECT 163.365 19.910 1194.095 20.210 ;
        RECT 163.365 19.895 163.695 19.910 ;
        RECT 1193.765 19.895 1194.095 19.910 ;
>>>>>>> re-updated local openlane
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 0.300 ;
=======
      LAYER li1 ;
        RECT 1149.225 17.425 1149.395 19.295 ;
      LAYER mcon ;
        RECT 1149.225 19.125 1149.395 19.295 ;
      LAYER met1 ;
        RECT 180.850 19.280 181.170 19.340 ;
        RECT 1149.165 19.280 1149.455 19.325 ;
        RECT 180.850 19.140 1149.455 19.280 ;
        RECT 180.850 19.080 181.170 19.140 ;
        RECT 1149.165 19.095 1149.455 19.140 ;
        RECT 1149.165 17.580 1149.455 17.625 ;
        RECT 1195.610 17.580 1195.930 17.640 ;
        RECT 1149.165 17.440 1195.930 17.580 ;
        RECT 1149.165 17.395 1149.455 17.440 ;
        RECT 1195.610 17.380 1195.930 17.440 ;
      LAYER via ;
        RECT 180.880 19.080 181.140 19.340 ;
        RECT 1195.640 17.380 1195.900 17.640 ;
      LAYER met2 ;
        RECT 1198.390 1700.410 1198.670 1704.000 ;
        RECT 1197.540 1700.270 1198.670 1700.410 ;
        RECT 1197.540 1678.140 1197.680 1700.270 ;
        RECT 1198.390 1700.000 1198.670 1700.270 ;
        RECT 1195.700 1678.000 1197.680 1678.140 ;
        RECT 180.880 19.050 181.140 19.370 ;
        RECT 180.940 2.400 181.080 19.050 ;
        RECT 1195.700 17.670 1195.840 1678.000 ;
        RECT 1195.640 17.350 1195.900 17.670 ;
=======
      LAYER met1 ;
        RECT 196.490 1688.680 196.810 1688.740 ;
        RECT 1198.830 1688.680 1199.150 1688.740 ;
        RECT 196.490 1688.540 1199.150 1688.680 ;
        RECT 196.490 1688.480 196.810 1688.540 ;
        RECT 1198.830 1688.480 1199.150 1688.540 ;
        RECT 180.850 16.220 181.170 16.280 ;
        RECT 196.490 16.220 196.810 16.280 ;
        RECT 180.850 16.080 196.810 16.220 ;
        RECT 180.850 16.020 181.170 16.080 ;
        RECT 196.490 16.020 196.810 16.080 ;
      LAYER via ;
        RECT 196.520 1688.480 196.780 1688.740 ;
        RECT 1198.860 1688.480 1199.120 1688.740 ;
        RECT 180.880 16.020 181.140 16.280 ;
        RECT 196.520 16.020 196.780 16.280 ;
      LAYER met2 ;
        RECT 1198.850 1700.000 1199.130 1704.000 ;
        RECT 1198.920 1688.770 1199.060 1700.000 ;
        RECT 196.520 1688.450 196.780 1688.770 ;
        RECT 1198.860 1688.450 1199.120 1688.770 ;
        RECT 196.580 16.310 196.720 1688.450 ;
        RECT 180.880 15.990 181.140 16.310 ;
        RECT 196.520 15.990 196.780 16.310 ;
        RECT 180.940 2.400 181.080 15.990 ;
>>>>>>> re-updated local openlane
        RECT 180.730 -4.800 181.290 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 0.300 ;
=======
      LAYER met1 ;
        RECT 1202.510 17.580 1202.830 17.640 ;
        RECT 1187.880 17.440 1202.830 17.580 ;
        RECT 198.790 17.240 199.110 17.300 ;
        RECT 1187.880 17.240 1188.020 17.440 ;
        RECT 1202.510 17.380 1202.830 17.440 ;
        RECT 198.790 17.100 1188.020 17.240 ;
        RECT 198.790 17.040 199.110 17.100 ;
      LAYER via ;
        RECT 198.820 17.040 199.080 17.300 ;
        RECT 1202.540 17.380 1202.800 17.640 ;
      LAYER met2 ;
        RECT 1203.450 1700.410 1203.730 1704.000 ;
        RECT 1202.600 1700.270 1203.730 1700.410 ;
        RECT 1202.600 17.670 1202.740 1700.270 ;
        RECT 1203.450 1700.000 1203.730 1700.270 ;
        RECT 1202.540 17.350 1202.800 17.670 ;
        RECT 198.820 17.010 199.080 17.330 ;
        RECT 198.880 2.400 199.020 17.010 ;
        RECT 198.670 -4.800 199.230 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 0.300 ;
=======
      LAYER met1 ;
        RECT 306.890 1689.360 307.210 1689.420 ;
        RECT 1208.490 1689.360 1208.810 1689.420 ;
        RECT 306.890 1689.220 1208.810 1689.360 ;
        RECT 306.890 1689.160 307.210 1689.220 ;
        RECT 1208.490 1689.160 1208.810 1689.220 ;
        RECT 216.730 19.280 217.050 19.340 ;
        RECT 306.890 19.280 307.210 19.340 ;
        RECT 216.730 19.140 307.210 19.280 ;
        RECT 216.730 19.080 217.050 19.140 ;
        RECT 306.890 19.080 307.210 19.140 ;
      LAYER via ;
        RECT 306.920 1689.160 307.180 1689.420 ;
        RECT 1208.520 1689.160 1208.780 1689.420 ;
        RECT 216.760 19.080 217.020 19.340 ;
        RECT 306.920 19.080 307.180 19.340 ;
      LAYER met2 ;
        RECT 1208.510 1700.000 1208.790 1704.000 ;
        RECT 1208.580 1689.450 1208.720 1700.000 ;
        RECT 306.920 1689.130 307.180 1689.450 ;
        RECT 1208.520 1689.130 1208.780 1689.450 ;
        RECT 306.980 19.370 307.120 1689.130 ;
        RECT 216.760 19.050 217.020 19.370 ;
        RECT 306.920 19.050 307.180 19.370 ;
        RECT 216.820 2.400 216.960 19.050 ;
        RECT 216.610 -4.800 217.170 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 0.300 ;
=======
      LAYER met1 ;
        RECT 1213.090 1688.340 1213.410 1688.400 ;
        RECT 1177.760 1688.200 1213.410 1688.340 ;
        RECT 241.110 1688.000 241.430 1688.060 ;
        RECT 1177.760 1688.000 1177.900 1688.200 ;
        RECT 1213.090 1688.140 1213.410 1688.200 ;
        RECT 241.110 1687.860 1177.900 1688.000 ;
        RECT 241.110 1687.800 241.430 1687.860 ;
        RECT 234.670 16.900 234.990 16.960 ;
        RECT 241.110 16.900 241.430 16.960 ;
        RECT 234.670 16.760 241.430 16.900 ;
        RECT 234.670 16.700 234.990 16.760 ;
        RECT 241.110 16.700 241.430 16.760 ;
      LAYER via ;
        RECT 241.140 1687.800 241.400 1688.060 ;
        RECT 1213.120 1688.140 1213.380 1688.400 ;
        RECT 234.700 16.700 234.960 16.960 ;
        RECT 241.140 16.700 241.400 16.960 ;
      LAYER met2 ;
        RECT 1213.110 1700.000 1213.390 1704.000 ;
        RECT 1213.180 1688.430 1213.320 1700.000 ;
        RECT 1213.120 1688.110 1213.380 1688.430 ;
        RECT 241.140 1687.770 241.400 1688.090 ;
        RECT 241.200 16.990 241.340 1687.770 ;
        RECT 234.700 16.670 234.960 16.990 ;
        RECT 241.140 16.670 241.400 16.990 ;
        RECT 234.760 2.400 234.900 16.670 ;
=======
      LAYER li1 ;
        RECT 1196.145 20.485 1197.695 20.655 ;
        RECT 1196.145 17.765 1196.315 20.485 ;
        RECT 1197.525 20.145 1197.695 20.485 ;
        RECT 269.245 16.405 269.415 17.595 ;
      LAYER mcon ;
        RECT 269.245 17.425 269.415 17.595 ;
      LAYER met1 ;
        RECT 1197.465 20.300 1197.755 20.345 ;
        RECT 1208.950 20.300 1209.270 20.360 ;
        RECT 1197.465 20.160 1209.270 20.300 ;
        RECT 1197.465 20.115 1197.755 20.160 ;
        RECT 1208.950 20.100 1209.270 20.160 ;
        RECT 1196.085 17.920 1196.375 17.965 ;
        RECT 1187.420 17.780 1196.375 17.920 ;
        RECT 269.185 17.580 269.475 17.625 ;
        RECT 1187.420 17.580 1187.560 17.780 ;
        RECT 1196.085 17.735 1196.375 17.780 ;
        RECT 269.185 17.440 1187.560 17.580 ;
        RECT 269.185 17.395 269.475 17.440 ;
        RECT 234.670 16.560 234.990 16.620 ;
        RECT 269.185 16.560 269.475 16.605 ;
        RECT 234.670 16.420 269.475 16.560 ;
        RECT 234.670 16.360 234.990 16.420 ;
        RECT 269.185 16.375 269.475 16.420 ;
      LAYER via ;
        RECT 1208.980 20.100 1209.240 20.360 ;
        RECT 234.700 16.360 234.960 16.620 ;
      LAYER met2 ;
        RECT 1213.110 1700.410 1213.390 1704.000 ;
        RECT 1212.720 1700.270 1213.390 1700.410 ;
        RECT 1212.720 1677.290 1212.860 1700.270 ;
        RECT 1213.110 1700.000 1213.390 1700.270 ;
        RECT 1209.040 1677.150 1212.860 1677.290 ;
        RECT 1209.040 20.390 1209.180 1677.150 ;
        RECT 1208.980 20.070 1209.240 20.390 ;
        RECT 234.700 16.330 234.960 16.650 ;
        RECT 234.760 2.400 234.900 16.330 ;
>>>>>>> re-updated local openlane
        RECT 234.550 -4.800 235.110 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 0.300 ;
=======
      LAYER met1 ;
        RECT 79.190 1688.000 79.510 1688.060 ;
        RECT 1164.790 1688.000 1165.110 1688.060 ;
        RECT 79.190 1687.860 1165.110 1688.000 ;
        RECT 79.190 1687.800 79.510 1687.860 ;
        RECT 1164.790 1687.800 1165.110 1687.860 ;
        RECT 56.190 17.580 56.510 17.640 ;
        RECT 79.190 17.580 79.510 17.640 ;
        RECT 56.190 17.440 79.510 17.580 ;
        RECT 56.190 17.380 56.510 17.440 ;
        RECT 79.190 17.380 79.510 17.440 ;
      LAYER via ;
        RECT 79.220 1687.800 79.480 1688.060 ;
        RECT 1164.820 1687.800 1165.080 1688.060 ;
        RECT 56.220 17.380 56.480 17.640 ;
        RECT 79.220 17.380 79.480 17.640 ;
      LAYER met2 ;
        RECT 1164.810 1700.000 1165.090 1704.000 ;
        RECT 1164.880 1688.090 1165.020 1700.000 ;
        RECT 79.220 1687.770 79.480 1688.090 ;
        RECT 1164.820 1687.770 1165.080 1688.090 ;
        RECT 79.280 17.670 79.420 1687.770 ;
        RECT 56.220 17.350 56.480 17.670 ;
        RECT 79.220 17.350 79.480 17.670 ;
        RECT 56.280 2.400 56.420 17.350 ;
        RECT 56.070 -4.800 56.630 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 56.210 17.880 56.490 18.160 ;
        RECT 1159.290 17.880 1159.570 18.160 ;
      LAYER met3 ;
        RECT 56.185 18.170 56.515 18.185 ;
        RECT 1159.265 18.170 1159.595 18.185 ;
        RECT 56.185 17.870 1159.595 18.170 ;
        RECT 56.185 17.855 56.515 17.870 ;
        RECT 1159.265 17.855 1159.595 17.870 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 0.300 ;
=======
      LAYER met1 ;
        RECT 1166.170 1678.140 1166.490 1678.200 ;
        RECT 1170.310 1678.140 1170.630 1678.200 ;
        RECT 1166.170 1678.000 1170.630 1678.140 ;
        RECT 1166.170 1677.940 1166.490 1678.000 ;
        RECT 1170.310 1677.940 1170.630 1678.000 ;
      LAYER via ;
        RECT 1166.200 1677.940 1166.460 1678.200 ;
        RECT 1170.340 1677.940 1170.600 1678.200 ;
      LAYER met2 ;
        RECT 1171.250 1700.410 1171.530 1704.000 ;
        RECT 1170.400 1700.270 1171.530 1700.410 ;
        RECT 1170.400 1678.230 1170.540 1700.270 ;
        RECT 1171.250 1700.000 1171.530 1700.270 ;
        RECT 1166.200 1677.910 1166.460 1678.230 ;
        RECT 1170.340 1677.910 1170.600 1678.230 ;
        RECT 1166.260 18.205 1166.400 1677.910 ;
        RECT 80.130 17.835 80.410 18.205 ;
        RECT 1166.190 17.835 1166.470 18.205 ;
        RECT 80.200 2.400 80.340 17.835 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 80.130 17.880 80.410 18.160 ;
        RECT 1166.190 17.880 1166.470 18.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 82.405 1687.570 82.735 1687.585 ;
        RECT 1171.225 1687.570 1171.555 1687.585 ;
        RECT 82.405 1687.270 1171.555 1687.570 ;
        RECT 82.405 1687.255 82.735 1687.270 ;
        RECT 1171.225 1687.255 1171.555 1687.270 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 80.105 18.170 80.435 18.185 ;
        RECT 1166.165 18.170 1166.495 18.185 ;
        RECT 80.105 17.870 1166.495 18.170 ;
        RECT 80.105 17.855 80.435 17.870 ;
        RECT 1166.165 17.855 1166.495 17.870 ;
>>>>>>> re-updated local openlane
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
<<<<<<< HEAD
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 0.300 ;
=======
      LAYER li1 ;
        RECT 1149.685 17.255 1149.855 19.295 ;
        RECT 1148.305 17.085 1149.855 17.255 ;
      LAYER mcon ;
        RECT 1149.685 19.125 1149.855 19.295 ;
      LAYER met1 ;
        RECT 1149.625 19.280 1149.915 19.325 ;
        RECT 1173.990 19.280 1174.310 19.340 ;
        RECT 1149.625 19.140 1174.310 19.280 ;
        RECT 1149.625 19.095 1149.915 19.140 ;
        RECT 1173.990 19.080 1174.310 19.140 ;
        RECT 103.570 17.240 103.890 17.300 ;
        RECT 1148.245 17.240 1148.535 17.285 ;
        RECT 103.570 17.100 1148.535 17.240 ;
        RECT 103.570 17.040 103.890 17.100 ;
        RECT 1148.245 17.055 1148.535 17.100 ;
      LAYER via ;
        RECT 1174.020 19.080 1174.280 19.340 ;
        RECT 103.600 17.040 103.860 17.300 ;
      LAYER met2 ;
        RECT 1177.690 1700.410 1177.970 1704.000 ;
        RECT 1176.380 1700.270 1177.970 1700.410 ;
        RECT 1176.380 1677.290 1176.520 1700.270 ;
        RECT 1177.690 1700.000 1177.970 1700.270 ;
        RECT 1174.080 1677.150 1176.520 1677.290 ;
        RECT 1174.080 19.370 1174.220 1677.150 ;
        RECT 1174.020 19.050 1174.280 19.370 ;
        RECT 103.600 17.010 103.860 17.330 ;
        RECT 103.660 2.400 103.800 17.010 ;
=======
      LAYER met1 ;
        RECT 210.290 1689.020 210.610 1689.080 ;
        RECT 1177.670 1689.020 1177.990 1689.080 ;
        RECT 210.290 1688.880 1177.990 1689.020 ;
        RECT 210.290 1688.820 210.610 1688.880 ;
        RECT 1177.670 1688.820 1177.990 1688.880 ;
        RECT 210.290 17.580 210.610 17.640 ;
        RECT 121.140 17.440 210.610 17.580 ;
        RECT 103.570 16.900 103.890 16.960 ;
        RECT 121.140 16.900 121.280 17.440 ;
        RECT 210.290 17.380 210.610 17.440 ;
        RECT 103.570 16.760 121.280 16.900 ;
        RECT 103.570 16.700 103.890 16.760 ;
      LAYER via ;
        RECT 210.320 1688.820 210.580 1689.080 ;
        RECT 1177.700 1688.820 1177.960 1689.080 ;
        RECT 103.600 16.700 103.860 16.960 ;
        RECT 210.320 17.380 210.580 17.640 ;
      LAYER met2 ;
        RECT 1177.690 1700.000 1177.970 1704.000 ;
        RECT 1177.760 1689.110 1177.900 1700.000 ;
        RECT 210.320 1688.790 210.580 1689.110 ;
        RECT 1177.700 1688.790 1177.960 1689.110 ;
        RECT 210.380 17.670 210.520 1688.790 ;
        RECT 210.320 17.350 210.580 17.670 ;
        RECT 103.600 16.670 103.860 16.990 ;
        RECT 103.660 2.400 103.800 16.670 ;
>>>>>>> re-updated local openlane
        RECT 103.450 -4.800 104.010 2.400 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 0.300 ;
=======
      LAYER met1 ;
        RECT 1180.430 1677.460 1180.750 1677.520 ;
        RECT 1183.190 1677.460 1183.510 1677.520 ;
        RECT 1180.430 1677.320 1183.510 1677.460 ;
        RECT 1180.430 1677.260 1180.750 1677.320 ;
        RECT 1183.190 1677.260 1183.510 1677.320 ;
      LAYER via ;
        RECT 1180.460 1677.260 1180.720 1677.520 ;
        RECT 1183.220 1677.260 1183.480 1677.520 ;
      LAYER met2 ;
        RECT 1184.130 1700.410 1184.410 1704.000 ;
        RECT 1183.280 1700.270 1184.410 1700.410 ;
        RECT 1183.280 1677.550 1183.420 1700.270 ;
        RECT 1184.130 1700.000 1184.410 1700.270 ;
        RECT 1180.460 1677.230 1180.720 1677.550 ;
        RECT 1183.220 1677.230 1183.480 1677.550 ;
        RECT 1180.520 19.565 1180.660 1677.230 ;
        RECT 127.510 19.195 127.790 19.565 ;
        RECT 1180.450 19.195 1180.730 19.565 ;
        RECT 127.580 2.400 127.720 19.195 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 127.510 19.240 127.790 19.520 ;
        RECT 1180.450 19.240 1180.730 19.520 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 130.705 1688.250 131.035 1688.265 ;
        RECT 1184.105 1688.250 1184.435 1688.265 ;
        RECT 130.705 1687.950 1184.435 1688.250 ;
        RECT 130.705 1687.935 131.035 1687.950 ;
        RECT 1184.105 1687.935 1184.435 1687.950 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 127.485 19.530 127.815 19.545 ;
        RECT 1180.425 19.530 1180.755 19.545 ;
        RECT 127.485 19.230 1180.755 19.530 ;
        RECT 127.485 19.215 127.815 19.230 ;
        RECT 1180.425 19.215 1180.755 19.230 ;
>>>>>>> re-updated local openlane
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 0.300 ;
=======
      LAYER met1 ;
        RECT 51.590 1686.980 51.910 1687.040 ;
        RECT 1156.970 1686.980 1157.290 1687.040 ;
        RECT 51.590 1686.840 1157.290 1686.980 ;
        RECT 51.590 1686.780 51.910 1686.840 ;
        RECT 1156.970 1686.780 1157.290 1686.840 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 51.590 17.240 51.910 17.300 ;
        RECT 26.290 17.100 51.910 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 51.590 17.040 51.910 17.100 ;
      LAYER via ;
        RECT 51.620 1686.780 51.880 1687.040 ;
        RECT 1157.000 1686.780 1157.260 1687.040 ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 51.620 17.040 51.880 17.300 ;
      LAYER met2 ;
        RECT 1156.990 1700.000 1157.270 1704.000 ;
        RECT 1157.060 1687.070 1157.200 1700.000 ;
        RECT 51.620 1686.750 51.880 1687.070 ;
        RECT 1157.000 1686.750 1157.260 1687.070 ;
        RECT 51.680 17.330 51.820 1686.750 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 51.620 17.010 51.880 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
<<<<<<< HEAD
      LAYER via2 ;
        RECT 26.310 16.520 26.590 16.800 ;
        RECT 1153.770 16.520 1154.050 16.800 ;
      LAYER met3 ;
        RECT 26.285 16.810 26.615 16.825 ;
        RECT 1153.745 16.810 1154.075 16.825 ;
        RECT 26.285 16.510 1154.075 16.810 ;
        RECT 26.285 16.495 26.615 16.510 ;
        RECT 1153.745 16.495 1154.075 16.510 ;
>>>>>>> Latest run - not LVS matched yet
=======
>>>>>>> re-updated local openlane
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
<<<<<<< HEAD
        RECT 32.150 -4.800 32.710 0.300 ;
=======
        RECT 1158.370 1700.000 1158.650 1704.000 ;
        RECT 1158.440 1686.925 1158.580 1700.000 ;
        RECT 34.130 1686.555 34.410 1686.925 ;
        RECT 1158.370 1686.555 1158.650 1686.925 ;
        RECT 34.200 3.130 34.340 1686.555 ;
        RECT 32.360 2.990 34.340 3.130 ;
        RECT 32.360 2.400 32.500 2.990 ;
=======
      LAYER li1 ;
        RECT 1154.285 1594.005 1154.455 1658.095 ;
        RECT 1154.285 786.505 1154.455 821.015 ;
        RECT 1154.285 689.605 1154.455 724.455 ;
        RECT 1154.285 593.045 1154.455 627.895 ;
        RECT 1154.285 496.485 1154.455 531.335 ;
        RECT 1154.285 386.325 1154.455 434.775 ;
        RECT 1154.285 351.645 1154.455 385.815 ;
        RECT 1154.285 255.085 1154.455 289.595 ;
        RECT 1154.285 158.525 1154.455 193.035 ;
      LAYER mcon ;
        RECT 1154.285 1657.925 1154.455 1658.095 ;
        RECT 1154.285 820.845 1154.455 821.015 ;
        RECT 1154.285 724.285 1154.455 724.455 ;
        RECT 1154.285 627.725 1154.455 627.895 ;
        RECT 1154.285 531.165 1154.455 531.335 ;
        RECT 1154.285 434.605 1154.455 434.775 ;
        RECT 1154.285 385.645 1154.455 385.815 ;
        RECT 1154.285 289.425 1154.455 289.595 ;
        RECT 1154.285 192.865 1154.455 193.035 ;
      LAYER met1 ;
        RECT 1154.225 1658.080 1154.515 1658.125 ;
        RECT 1157.430 1658.080 1157.750 1658.140 ;
        RECT 1154.225 1657.940 1157.750 1658.080 ;
        RECT 1154.225 1657.895 1154.515 1657.940 ;
        RECT 1157.430 1657.880 1157.750 1657.940 ;
        RECT 1154.210 1594.160 1154.530 1594.220 ;
        RECT 1154.015 1594.020 1154.530 1594.160 ;
        RECT 1154.210 1593.960 1154.530 1594.020 ;
        RECT 1153.750 1414.640 1154.070 1414.700 ;
        RECT 1154.670 1414.640 1154.990 1414.700 ;
        RECT 1153.750 1414.500 1154.990 1414.640 ;
        RECT 1153.750 1414.440 1154.070 1414.500 ;
        RECT 1154.670 1414.440 1154.990 1414.500 ;
        RECT 1153.750 1318.080 1154.070 1318.140 ;
        RECT 1154.670 1318.080 1154.990 1318.140 ;
        RECT 1153.750 1317.940 1154.990 1318.080 ;
        RECT 1153.750 1317.880 1154.070 1317.940 ;
        RECT 1154.670 1317.880 1154.990 1317.940 ;
        RECT 1153.750 1221.520 1154.070 1221.580 ;
        RECT 1154.670 1221.520 1154.990 1221.580 ;
        RECT 1153.750 1221.380 1154.990 1221.520 ;
        RECT 1153.750 1221.320 1154.070 1221.380 ;
        RECT 1154.670 1221.320 1154.990 1221.380 ;
        RECT 1153.750 1124.960 1154.070 1125.020 ;
        RECT 1154.670 1124.960 1154.990 1125.020 ;
        RECT 1153.750 1124.820 1154.990 1124.960 ;
        RECT 1153.750 1124.760 1154.070 1124.820 ;
        RECT 1154.670 1124.760 1154.990 1124.820 ;
        RECT 1153.750 1028.400 1154.070 1028.460 ;
        RECT 1154.670 1028.400 1154.990 1028.460 ;
        RECT 1153.750 1028.260 1154.990 1028.400 ;
        RECT 1153.750 1028.200 1154.070 1028.260 ;
        RECT 1154.670 1028.200 1154.990 1028.260 ;
        RECT 1153.750 931.840 1154.070 931.900 ;
        RECT 1154.670 931.840 1154.990 931.900 ;
        RECT 1153.750 931.700 1154.990 931.840 ;
        RECT 1153.750 931.640 1154.070 931.700 ;
        RECT 1154.670 931.640 1154.990 931.700 ;
        RECT 1154.670 869.620 1154.990 869.680 ;
        RECT 1155.590 869.620 1155.910 869.680 ;
        RECT 1154.670 869.480 1155.910 869.620 ;
        RECT 1154.670 869.420 1154.990 869.480 ;
        RECT 1155.590 869.420 1155.910 869.480 ;
        RECT 1153.750 835.280 1154.070 835.340 ;
        RECT 1154.670 835.280 1154.990 835.340 ;
        RECT 1153.750 835.140 1154.990 835.280 ;
        RECT 1153.750 835.080 1154.070 835.140 ;
        RECT 1154.670 835.080 1154.990 835.140 ;
        RECT 1154.210 821.000 1154.530 821.060 ;
        RECT 1154.015 820.860 1154.530 821.000 ;
        RECT 1154.210 820.800 1154.530 820.860 ;
        RECT 1154.210 786.660 1154.530 786.720 ;
        RECT 1154.015 786.520 1154.530 786.660 ;
        RECT 1154.210 786.460 1154.530 786.520 ;
        RECT 1153.750 738.380 1154.070 738.440 ;
        RECT 1154.670 738.380 1154.990 738.440 ;
        RECT 1153.750 738.240 1154.990 738.380 ;
        RECT 1153.750 738.180 1154.070 738.240 ;
        RECT 1154.670 738.180 1154.990 738.240 ;
        RECT 1154.210 724.440 1154.530 724.500 ;
        RECT 1154.015 724.300 1154.530 724.440 ;
        RECT 1154.210 724.240 1154.530 724.300 ;
        RECT 1154.210 689.760 1154.530 689.820 ;
        RECT 1154.015 689.620 1154.530 689.760 ;
        RECT 1154.210 689.560 1154.530 689.620 ;
        RECT 1153.750 641.820 1154.070 641.880 ;
        RECT 1154.670 641.820 1154.990 641.880 ;
        RECT 1153.750 641.680 1154.990 641.820 ;
        RECT 1153.750 641.620 1154.070 641.680 ;
        RECT 1154.670 641.620 1154.990 641.680 ;
        RECT 1154.210 627.880 1154.530 627.940 ;
        RECT 1154.015 627.740 1154.530 627.880 ;
        RECT 1154.210 627.680 1154.530 627.740 ;
        RECT 1154.210 593.200 1154.530 593.260 ;
        RECT 1154.015 593.060 1154.530 593.200 ;
        RECT 1154.210 593.000 1154.530 593.060 ;
        RECT 1153.750 545.260 1154.070 545.320 ;
        RECT 1154.670 545.260 1154.990 545.320 ;
        RECT 1153.750 545.120 1154.990 545.260 ;
        RECT 1153.750 545.060 1154.070 545.120 ;
        RECT 1154.670 545.060 1154.990 545.120 ;
        RECT 1154.210 531.320 1154.530 531.380 ;
        RECT 1154.015 531.180 1154.530 531.320 ;
        RECT 1154.210 531.120 1154.530 531.180 ;
        RECT 1154.210 496.640 1154.530 496.700 ;
        RECT 1154.015 496.500 1154.530 496.640 ;
        RECT 1154.210 496.440 1154.530 496.500 ;
        RECT 1153.750 448.700 1154.070 448.760 ;
        RECT 1154.670 448.700 1154.990 448.760 ;
        RECT 1153.750 448.560 1154.990 448.700 ;
        RECT 1153.750 448.500 1154.070 448.560 ;
        RECT 1154.670 448.500 1154.990 448.560 ;
        RECT 1154.210 434.760 1154.530 434.820 ;
        RECT 1154.015 434.620 1154.530 434.760 ;
        RECT 1154.210 434.560 1154.530 434.620 ;
        RECT 1154.225 386.480 1154.515 386.525 ;
        RECT 1154.670 386.480 1154.990 386.540 ;
        RECT 1154.225 386.340 1154.990 386.480 ;
        RECT 1154.225 386.295 1154.515 386.340 ;
        RECT 1154.670 386.280 1154.990 386.340 ;
        RECT 1154.225 385.800 1154.515 385.845 ;
        RECT 1154.670 385.800 1154.990 385.860 ;
        RECT 1154.225 385.660 1154.990 385.800 ;
        RECT 1154.225 385.615 1154.515 385.660 ;
        RECT 1154.670 385.600 1154.990 385.660 ;
        RECT 1154.210 351.800 1154.530 351.860 ;
        RECT 1154.015 351.660 1154.530 351.800 ;
        RECT 1154.210 351.600 1154.530 351.660 ;
        RECT 1154.225 289.580 1154.515 289.625 ;
        RECT 1154.670 289.580 1154.990 289.640 ;
        RECT 1154.225 289.440 1154.990 289.580 ;
        RECT 1154.225 289.395 1154.515 289.440 ;
        RECT 1154.670 289.380 1154.990 289.440 ;
        RECT 1154.210 255.240 1154.530 255.300 ;
        RECT 1154.015 255.100 1154.530 255.240 ;
        RECT 1154.210 255.040 1154.530 255.100 ;
        RECT 1154.225 193.020 1154.515 193.065 ;
        RECT 1154.670 193.020 1154.990 193.080 ;
        RECT 1154.225 192.880 1154.990 193.020 ;
        RECT 1154.225 192.835 1154.515 192.880 ;
        RECT 1154.670 192.820 1154.990 192.880 ;
        RECT 1154.210 158.680 1154.530 158.740 ;
        RECT 1154.015 158.540 1154.530 158.680 ;
        RECT 1154.210 158.480 1154.530 158.540 ;
      LAYER via ;
        RECT 1157.460 1657.880 1157.720 1658.140 ;
        RECT 1154.240 1593.960 1154.500 1594.220 ;
        RECT 1153.780 1414.440 1154.040 1414.700 ;
        RECT 1154.700 1414.440 1154.960 1414.700 ;
        RECT 1153.780 1317.880 1154.040 1318.140 ;
        RECT 1154.700 1317.880 1154.960 1318.140 ;
        RECT 1153.780 1221.320 1154.040 1221.580 ;
        RECT 1154.700 1221.320 1154.960 1221.580 ;
        RECT 1153.780 1124.760 1154.040 1125.020 ;
        RECT 1154.700 1124.760 1154.960 1125.020 ;
        RECT 1153.780 1028.200 1154.040 1028.460 ;
        RECT 1154.700 1028.200 1154.960 1028.460 ;
        RECT 1153.780 931.640 1154.040 931.900 ;
        RECT 1154.700 931.640 1154.960 931.900 ;
        RECT 1154.700 869.420 1154.960 869.680 ;
        RECT 1155.620 869.420 1155.880 869.680 ;
        RECT 1153.780 835.080 1154.040 835.340 ;
        RECT 1154.700 835.080 1154.960 835.340 ;
        RECT 1154.240 820.800 1154.500 821.060 ;
        RECT 1154.240 786.460 1154.500 786.720 ;
        RECT 1153.780 738.180 1154.040 738.440 ;
        RECT 1154.700 738.180 1154.960 738.440 ;
        RECT 1154.240 724.240 1154.500 724.500 ;
        RECT 1154.240 689.560 1154.500 689.820 ;
        RECT 1153.780 641.620 1154.040 641.880 ;
        RECT 1154.700 641.620 1154.960 641.880 ;
        RECT 1154.240 627.680 1154.500 627.940 ;
        RECT 1154.240 593.000 1154.500 593.260 ;
        RECT 1153.780 545.060 1154.040 545.320 ;
        RECT 1154.700 545.060 1154.960 545.320 ;
        RECT 1154.240 531.120 1154.500 531.380 ;
        RECT 1154.240 496.440 1154.500 496.700 ;
        RECT 1153.780 448.500 1154.040 448.760 ;
        RECT 1154.700 448.500 1154.960 448.760 ;
        RECT 1154.240 434.560 1154.500 434.820 ;
        RECT 1154.700 386.280 1154.960 386.540 ;
        RECT 1154.700 385.600 1154.960 385.860 ;
        RECT 1154.240 351.600 1154.500 351.860 ;
        RECT 1154.700 289.380 1154.960 289.640 ;
        RECT 1154.240 255.040 1154.500 255.300 ;
        RECT 1154.700 192.820 1154.960 193.080 ;
        RECT 1154.240 158.480 1154.500 158.740 ;
      LAYER met2 ;
        RECT 1158.370 1700.410 1158.650 1704.000 ;
        RECT 1157.520 1700.270 1158.650 1700.410 ;
        RECT 1157.520 1658.170 1157.660 1700.270 ;
        RECT 1158.370 1700.000 1158.650 1700.270 ;
        RECT 1157.460 1657.850 1157.720 1658.170 ;
        RECT 1154.240 1593.930 1154.500 1594.250 ;
        RECT 1154.300 1569.170 1154.440 1593.930 ;
        RECT 1154.300 1569.030 1154.900 1569.170 ;
        RECT 1154.760 1414.730 1154.900 1569.030 ;
        RECT 1153.780 1414.410 1154.040 1414.730 ;
        RECT 1154.700 1414.410 1154.960 1414.730 ;
        RECT 1153.840 1414.130 1153.980 1414.410 ;
        RECT 1153.840 1413.990 1154.440 1414.130 ;
        RECT 1154.300 1366.530 1154.440 1413.990 ;
        RECT 1154.300 1366.390 1154.900 1366.530 ;
        RECT 1154.760 1318.170 1154.900 1366.390 ;
        RECT 1153.780 1317.850 1154.040 1318.170 ;
        RECT 1154.700 1317.850 1154.960 1318.170 ;
        RECT 1153.840 1317.570 1153.980 1317.850 ;
        RECT 1153.840 1317.430 1154.440 1317.570 ;
        RECT 1154.300 1269.970 1154.440 1317.430 ;
        RECT 1154.300 1269.830 1154.900 1269.970 ;
        RECT 1154.760 1221.610 1154.900 1269.830 ;
        RECT 1153.780 1221.290 1154.040 1221.610 ;
        RECT 1154.700 1221.290 1154.960 1221.610 ;
        RECT 1153.840 1221.010 1153.980 1221.290 ;
        RECT 1153.840 1220.870 1154.440 1221.010 ;
        RECT 1154.300 1173.410 1154.440 1220.870 ;
        RECT 1154.300 1173.270 1154.900 1173.410 ;
        RECT 1154.760 1125.050 1154.900 1173.270 ;
        RECT 1153.780 1124.730 1154.040 1125.050 ;
        RECT 1154.700 1124.730 1154.960 1125.050 ;
        RECT 1153.840 1124.450 1153.980 1124.730 ;
        RECT 1153.840 1124.310 1154.440 1124.450 ;
        RECT 1154.300 1076.850 1154.440 1124.310 ;
        RECT 1154.300 1076.710 1154.900 1076.850 ;
        RECT 1154.760 1028.490 1154.900 1076.710 ;
        RECT 1153.780 1028.170 1154.040 1028.490 ;
        RECT 1154.700 1028.170 1154.960 1028.490 ;
        RECT 1153.840 1027.890 1153.980 1028.170 ;
        RECT 1153.840 1027.750 1154.440 1027.890 ;
        RECT 1154.300 980.290 1154.440 1027.750 ;
        RECT 1154.300 980.150 1154.900 980.290 ;
        RECT 1154.760 931.930 1154.900 980.150 ;
        RECT 1153.780 931.610 1154.040 931.930 ;
        RECT 1154.700 931.610 1154.960 931.930 ;
        RECT 1153.840 931.330 1153.980 931.610 ;
        RECT 1153.840 931.190 1154.440 931.330 ;
        RECT 1154.300 917.845 1154.440 931.190 ;
        RECT 1154.230 917.475 1154.510 917.845 ;
        RECT 1155.610 917.475 1155.890 917.845 ;
        RECT 1155.680 869.710 1155.820 917.475 ;
        RECT 1154.700 869.390 1154.960 869.710 ;
        RECT 1155.620 869.390 1155.880 869.710 ;
        RECT 1154.760 835.370 1154.900 869.390 ;
        RECT 1153.780 835.050 1154.040 835.370 ;
        RECT 1154.700 835.050 1154.960 835.370 ;
        RECT 1153.840 834.770 1153.980 835.050 ;
        RECT 1153.840 834.630 1154.440 834.770 ;
        RECT 1154.300 821.090 1154.440 834.630 ;
        RECT 1154.240 820.770 1154.500 821.090 ;
        RECT 1154.240 786.430 1154.500 786.750 ;
        RECT 1154.300 772.890 1154.440 786.430 ;
        RECT 1154.300 772.750 1154.900 772.890 ;
        RECT 1154.760 738.470 1154.900 772.750 ;
        RECT 1153.780 738.210 1154.040 738.470 ;
        RECT 1153.780 738.150 1154.440 738.210 ;
        RECT 1154.700 738.150 1154.960 738.470 ;
        RECT 1153.840 738.070 1154.440 738.150 ;
        RECT 1154.300 724.530 1154.440 738.070 ;
        RECT 1154.240 724.210 1154.500 724.530 ;
        RECT 1154.240 689.530 1154.500 689.850 ;
        RECT 1154.300 676.330 1154.440 689.530 ;
        RECT 1154.300 676.190 1154.900 676.330 ;
        RECT 1154.760 641.910 1154.900 676.190 ;
        RECT 1153.780 641.650 1154.040 641.910 ;
        RECT 1153.780 641.590 1154.440 641.650 ;
        RECT 1154.700 641.590 1154.960 641.910 ;
        RECT 1153.840 641.510 1154.440 641.590 ;
        RECT 1154.300 627.970 1154.440 641.510 ;
        RECT 1154.240 627.650 1154.500 627.970 ;
        RECT 1154.240 592.970 1154.500 593.290 ;
        RECT 1154.300 579.770 1154.440 592.970 ;
        RECT 1154.300 579.630 1154.900 579.770 ;
        RECT 1154.760 545.350 1154.900 579.630 ;
        RECT 1153.780 545.090 1154.040 545.350 ;
        RECT 1153.780 545.030 1154.440 545.090 ;
        RECT 1154.700 545.030 1154.960 545.350 ;
        RECT 1153.840 544.950 1154.440 545.030 ;
        RECT 1154.300 531.410 1154.440 544.950 ;
        RECT 1154.240 531.090 1154.500 531.410 ;
        RECT 1154.240 496.410 1154.500 496.730 ;
        RECT 1154.300 483.210 1154.440 496.410 ;
        RECT 1154.300 483.070 1154.900 483.210 ;
        RECT 1154.760 448.790 1154.900 483.070 ;
        RECT 1153.780 448.530 1154.040 448.790 ;
        RECT 1153.780 448.470 1154.440 448.530 ;
        RECT 1154.700 448.470 1154.960 448.790 ;
        RECT 1153.840 448.390 1154.440 448.470 ;
        RECT 1154.300 434.850 1154.440 448.390 ;
        RECT 1154.240 434.530 1154.500 434.850 ;
        RECT 1154.700 386.250 1154.960 386.570 ;
        RECT 1154.760 385.890 1154.900 386.250 ;
        RECT 1154.700 385.570 1154.960 385.890 ;
        RECT 1154.240 351.570 1154.500 351.890 ;
        RECT 1154.300 303.690 1154.440 351.570 ;
        RECT 1154.300 303.550 1154.900 303.690 ;
        RECT 1154.760 289.670 1154.900 303.550 ;
        RECT 1154.700 289.350 1154.960 289.670 ;
        RECT 1154.240 255.010 1154.500 255.330 ;
        RECT 1154.300 207.130 1154.440 255.010 ;
        RECT 1154.300 206.990 1154.900 207.130 ;
        RECT 1154.760 193.110 1154.900 206.990 ;
        RECT 1154.700 192.790 1154.960 193.110 ;
        RECT 1154.240 158.450 1154.500 158.770 ;
        RECT 1154.300 110.570 1154.440 158.450 ;
        RECT 1154.300 110.430 1154.900 110.570 ;
        RECT 1154.760 62.290 1154.900 110.430 ;
        RECT 1153.840 62.150 1154.900 62.290 ;
        RECT 1153.840 16.845 1153.980 62.150 ;
        RECT 32.290 16.475 32.570 16.845 ;
        RECT 1153.770 16.475 1154.050 16.845 ;
        RECT 32.360 2.400 32.500 16.475 ;
>>>>>>> re-updated local openlane
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 1154.230 917.520 1154.510 917.800 ;
        RECT 1155.610 917.520 1155.890 917.800 ;
        RECT 32.290 16.520 32.570 16.800 ;
        RECT 1153.770 16.520 1154.050 16.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 34.105 1686.890 34.435 1686.905 ;
        RECT 1158.345 1686.890 1158.675 1686.905 ;
        RECT 34.105 1686.590 1158.675 1686.890 ;
        RECT 34.105 1686.575 34.435 1686.590 ;
        RECT 1158.345 1686.575 1158.675 1686.590 ;
>>>>>>> Latest run - not LVS matched yet
=======
        RECT 1154.205 917.810 1154.535 917.825 ;
        RECT 1155.585 917.810 1155.915 917.825 ;
        RECT 1154.205 917.510 1155.915 917.810 ;
        RECT 1154.205 917.495 1154.535 917.510 ;
        RECT 1155.585 917.495 1155.915 917.510 ;
        RECT 32.265 16.810 32.595 16.825 ;
        RECT 1153.745 16.810 1154.075 16.825 ;
        RECT 32.265 16.510 1154.075 16.810 ;
        RECT 32.265 16.495 32.595 16.510 ;
        RECT 1153.745 16.495 1154.075 16.510 ;
>>>>>>> re-updated local openlane
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
<<<<<<< HEAD
        RECT 4.020 3519.700 7.020 3529.000 ;
        RECT 184.020 3519.700 187.020 3529.000 ;
        RECT 364.020 3519.700 367.020 3529.000 ;
        RECT 544.020 3519.700 547.020 3529.000 ;
        RECT 724.020 3519.700 727.020 3529.000 ;
        RECT 904.020 3519.700 907.020 3529.000 ;
        RECT 1084.020 3519.700 1087.020 3529.000 ;
        RECT 1264.020 3519.700 1267.020 3529.000 ;
        RECT 1444.020 3519.700 1447.020 3529.000 ;
        RECT 1624.020 3519.700 1627.020 3529.000 ;
        RECT 1804.020 3519.700 1807.020 3529.000 ;
        RECT 1984.020 3519.700 1987.020 3529.000 ;
        RECT 2164.020 3519.700 2167.020 3529.000 ;
        RECT 2344.020 3519.700 2347.020 3529.000 ;
        RECT 2524.020 3519.700 2527.020 3529.000 ;
        RECT 2704.020 3519.700 2707.020 3529.000 ;
        RECT 2884.020 3519.700 2887.020 3529.000 ;
        RECT 4.020 -9.320 7.020 0.300 ;
        RECT 184.020 -9.320 187.020 0.300 ;
        RECT 364.020 -9.320 367.020 0.300 ;
        RECT 544.020 -9.320 547.020 0.300 ;
        RECT 724.020 -9.320 727.020 0.300 ;
        RECT 904.020 -9.320 907.020 0.300 ;
        RECT 1084.020 -9.320 1087.020 0.300 ;
        RECT 1264.020 -9.320 1267.020 0.300 ;
        RECT 1444.020 -9.320 1447.020 0.300 ;
        RECT 1624.020 -9.320 1627.020 0.300 ;
        RECT 1804.020 -9.320 1807.020 0.300 ;
        RECT 1984.020 -9.320 1987.020 0.300 ;
        RECT 2164.020 -9.320 2167.020 0.300 ;
        RECT 2344.020 -9.320 2347.020 0.300 ;
        RECT 2524.020 -9.320 2527.020 0.300 ;
        RECT 2704.020 -9.320 2707.020 0.300 ;
        RECT 2884.020 -9.320 2887.020 0.300 ;
=======
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 -9.220 547.020 3528.900 ;
        RECT 724.020 -9.220 727.020 3528.900 ;
        RECT 904.020 -9.220 907.020 3528.900 ;
        RECT 1084.020 -9.220 1087.020 3528.900 ;
        RECT 1264.020 -9.220 1267.020 3528.900 ;
        RECT 1444.020 -9.220 1447.020 3528.900 ;
        RECT 1624.020 -9.220 1627.020 3528.900 ;
        RECT 1804.020 -9.220 1807.020 3528.900 ;
        RECT 1984.020 -9.220 1987.020 3528.900 ;
        RECT 2164.020 -9.220 2167.020 3528.900 ;
        RECT 2344.020 -9.220 2347.020 3528.900 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
>>>>>>> Latest run - not LVS matched yet
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
<<<<<<< HEAD
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT -9.070 3430.850 -7.890 3432.030 ;
        RECT -9.070 3429.250 -7.890 3430.430 ;
        RECT -9.070 3250.850 -7.890 3252.030 ;
        RECT -9.070 3249.250 -7.890 3250.430 ;
        RECT -9.070 3070.850 -7.890 3072.030 ;
        RECT -9.070 3069.250 -7.890 3070.430 ;
        RECT -9.070 2890.850 -7.890 2892.030 ;
        RECT -9.070 2889.250 -7.890 2890.430 ;
        RECT -9.070 2710.850 -7.890 2712.030 ;
        RECT -9.070 2709.250 -7.890 2710.430 ;
        RECT -9.070 2530.850 -7.890 2532.030 ;
        RECT -9.070 2529.250 -7.890 2530.430 ;
        RECT -9.070 2350.850 -7.890 2352.030 ;
        RECT -9.070 2349.250 -7.890 2350.430 ;
        RECT -9.070 2170.850 -7.890 2172.030 ;
        RECT -9.070 2169.250 -7.890 2170.430 ;
        RECT -9.070 1990.850 -7.890 1992.030 ;
        RECT -9.070 1989.250 -7.890 1990.430 ;
        RECT -9.070 1810.850 -7.890 1812.030 ;
        RECT -9.070 1809.250 -7.890 1810.430 ;
        RECT -9.070 1630.850 -7.890 1632.030 ;
        RECT -9.070 1629.250 -7.890 1630.430 ;
        RECT -9.070 1450.850 -7.890 1452.030 ;
        RECT -9.070 1449.250 -7.890 1450.430 ;
        RECT -9.070 1270.850 -7.890 1272.030 ;
        RECT -9.070 1269.250 -7.890 1270.430 ;
        RECT -9.070 1090.850 -7.890 1092.030 ;
        RECT -9.070 1089.250 -7.890 1090.430 ;
        RECT -9.070 910.850 -7.890 912.030 ;
        RECT -9.070 909.250 -7.890 910.430 ;
        RECT -9.070 730.850 -7.890 732.030 ;
        RECT -9.070 729.250 -7.890 730.430 ;
        RECT -9.070 550.850 -7.890 552.030 ;
        RECT -9.070 549.250 -7.890 550.430 ;
        RECT -9.070 370.850 -7.890 372.030 ;
        RECT -9.070 369.250 -7.890 370.430 ;
        RECT -9.070 190.850 -7.890 192.030 ;
        RECT -9.070 189.250 -7.890 190.430 ;
        RECT -9.070 10.850 -7.890 12.030 ;
        RECT -9.070 9.250 -7.890 10.430 ;
        RECT 2927.510 3430.850 2928.690 3432.030 ;
        RECT 2927.510 3429.250 2928.690 3430.430 ;
        RECT 2927.510 3250.850 2928.690 3252.030 ;
        RECT 2927.510 3249.250 2928.690 3250.430 ;
        RECT 2927.510 3070.850 2928.690 3072.030 ;
        RECT 2927.510 3069.250 2928.690 3070.430 ;
        RECT 2927.510 2890.850 2928.690 2892.030 ;
        RECT 2927.510 2889.250 2928.690 2890.430 ;
        RECT 2927.510 2710.850 2928.690 2712.030 ;
        RECT 2927.510 2709.250 2928.690 2710.430 ;
        RECT 2927.510 2530.850 2928.690 2532.030 ;
        RECT 2927.510 2529.250 2928.690 2530.430 ;
        RECT 2927.510 2350.850 2928.690 2352.030 ;
        RECT 2927.510 2349.250 2928.690 2350.430 ;
        RECT 2927.510 2170.850 2928.690 2172.030 ;
        RECT 2927.510 2169.250 2928.690 2170.430 ;
        RECT 2927.510 1990.850 2928.690 1992.030 ;
        RECT 2927.510 1989.250 2928.690 1990.430 ;
        RECT 2927.510 1810.850 2928.690 1812.030 ;
        RECT 2927.510 1809.250 2928.690 1810.430 ;
        RECT 2927.510 1630.850 2928.690 1632.030 ;
        RECT 2927.510 1629.250 2928.690 1630.430 ;
        RECT 2927.510 1450.850 2928.690 1452.030 ;
        RECT 2927.510 1449.250 2928.690 1450.430 ;
        RECT 2927.510 1270.850 2928.690 1272.030 ;
        RECT 2927.510 1269.250 2928.690 1270.430 ;
        RECT 2927.510 1090.850 2928.690 1092.030 ;
        RECT 2927.510 1089.250 2928.690 1090.430 ;
        RECT 2927.510 910.850 2928.690 912.030 ;
        RECT 2927.510 909.250 2928.690 910.430 ;
        RECT 2927.510 730.850 2928.690 732.030 ;
        RECT 2927.510 729.250 2928.690 730.430 ;
        RECT 2927.510 550.850 2928.690 552.030 ;
        RECT 2927.510 549.250 2928.690 550.430 ;
        RECT 2927.510 370.850 2928.690 372.030 ;
        RECT 2927.510 369.250 2928.690 370.430 ;
        RECT 2927.510 190.850 2928.690 192.030 ;
        RECT 2927.510 189.250 2928.690 190.430 ;
        RECT 2927.510 10.850 2928.690 12.030 ;
        RECT 2927.510 9.250 2928.690 10.430 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
=======
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
>>>>>>> Latest run - not LVS matched yet
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
<<<<<<< HEAD
        RECT -9.980 3432.140 -6.980 3432.150 ;
        RECT 2926.600 3432.140 2929.600 3432.150 ;
        RECT -14.680 3429.140 0.300 3432.140 ;
        RECT 2919.700 3429.140 2934.300 3432.140 ;
        RECT -9.980 3429.130 -6.980 3429.140 ;
        RECT 2926.600 3429.130 2929.600 3429.140 ;
        RECT -9.980 3252.140 -6.980 3252.150 ;
        RECT 2926.600 3252.140 2929.600 3252.150 ;
        RECT -14.680 3249.140 0.300 3252.140 ;
        RECT 2919.700 3249.140 2934.300 3252.140 ;
        RECT -9.980 3249.130 -6.980 3249.140 ;
        RECT 2926.600 3249.130 2929.600 3249.140 ;
        RECT -9.980 3072.140 -6.980 3072.150 ;
        RECT 2926.600 3072.140 2929.600 3072.150 ;
        RECT -14.680 3069.140 0.300 3072.140 ;
        RECT 2919.700 3069.140 2934.300 3072.140 ;
        RECT -9.980 3069.130 -6.980 3069.140 ;
        RECT 2926.600 3069.130 2929.600 3069.140 ;
        RECT -9.980 2892.140 -6.980 2892.150 ;
        RECT 2926.600 2892.140 2929.600 2892.150 ;
        RECT -14.680 2889.140 0.300 2892.140 ;
        RECT 2919.700 2889.140 2934.300 2892.140 ;
        RECT -9.980 2889.130 -6.980 2889.140 ;
        RECT 2926.600 2889.130 2929.600 2889.140 ;
        RECT -9.980 2712.140 -6.980 2712.150 ;
        RECT 2926.600 2712.140 2929.600 2712.150 ;
        RECT -14.680 2709.140 0.300 2712.140 ;
        RECT 2919.700 2709.140 2934.300 2712.140 ;
        RECT -9.980 2709.130 -6.980 2709.140 ;
        RECT 2926.600 2709.130 2929.600 2709.140 ;
        RECT -9.980 2532.140 -6.980 2532.150 ;
        RECT 2926.600 2532.140 2929.600 2532.150 ;
        RECT -14.680 2529.140 0.300 2532.140 ;
        RECT 2919.700 2529.140 2934.300 2532.140 ;
        RECT -9.980 2529.130 -6.980 2529.140 ;
        RECT 2926.600 2529.130 2929.600 2529.140 ;
        RECT -9.980 2352.140 -6.980 2352.150 ;
        RECT 2926.600 2352.140 2929.600 2352.150 ;
        RECT -14.680 2349.140 0.300 2352.140 ;
        RECT 2919.700 2349.140 2934.300 2352.140 ;
        RECT -9.980 2349.130 -6.980 2349.140 ;
        RECT 2926.600 2349.130 2929.600 2349.140 ;
        RECT -9.980 2172.140 -6.980 2172.150 ;
        RECT 2926.600 2172.140 2929.600 2172.150 ;
        RECT -14.680 2169.140 0.300 2172.140 ;
        RECT 2919.700 2169.140 2934.300 2172.140 ;
        RECT -9.980 2169.130 -6.980 2169.140 ;
        RECT 2926.600 2169.130 2929.600 2169.140 ;
        RECT -9.980 1992.140 -6.980 1992.150 ;
        RECT 2926.600 1992.140 2929.600 1992.150 ;
        RECT -14.680 1989.140 0.300 1992.140 ;
        RECT 2919.700 1989.140 2934.300 1992.140 ;
        RECT -9.980 1989.130 -6.980 1989.140 ;
        RECT 2926.600 1989.130 2929.600 1989.140 ;
        RECT -9.980 1812.140 -6.980 1812.150 ;
        RECT 2926.600 1812.140 2929.600 1812.150 ;
        RECT -14.680 1809.140 0.300 1812.140 ;
        RECT 2919.700 1809.140 2934.300 1812.140 ;
        RECT -9.980 1809.130 -6.980 1809.140 ;
        RECT 2926.600 1809.130 2929.600 1809.140 ;
        RECT -9.980 1632.140 -6.980 1632.150 ;
        RECT 2926.600 1632.140 2929.600 1632.150 ;
        RECT -14.680 1629.140 0.300 1632.140 ;
        RECT 2919.700 1629.140 2934.300 1632.140 ;
        RECT -9.980 1629.130 -6.980 1629.140 ;
        RECT 2926.600 1629.130 2929.600 1629.140 ;
        RECT -9.980 1452.140 -6.980 1452.150 ;
        RECT 2926.600 1452.140 2929.600 1452.150 ;
        RECT -14.680 1449.140 0.300 1452.140 ;
        RECT 2919.700 1449.140 2934.300 1452.140 ;
        RECT -9.980 1449.130 -6.980 1449.140 ;
        RECT 2926.600 1449.130 2929.600 1449.140 ;
        RECT -9.980 1272.140 -6.980 1272.150 ;
        RECT 2926.600 1272.140 2929.600 1272.150 ;
        RECT -14.680 1269.140 0.300 1272.140 ;
        RECT 2919.700 1269.140 2934.300 1272.140 ;
        RECT -9.980 1269.130 -6.980 1269.140 ;
        RECT 2926.600 1269.130 2929.600 1269.140 ;
        RECT -9.980 1092.140 -6.980 1092.150 ;
        RECT 2926.600 1092.140 2929.600 1092.150 ;
        RECT -14.680 1089.140 0.300 1092.140 ;
        RECT 2919.700 1089.140 2934.300 1092.140 ;
        RECT -9.980 1089.130 -6.980 1089.140 ;
        RECT 2926.600 1089.130 2929.600 1089.140 ;
        RECT -9.980 912.140 -6.980 912.150 ;
        RECT 2926.600 912.140 2929.600 912.150 ;
        RECT -14.680 909.140 0.300 912.140 ;
        RECT 2919.700 909.140 2934.300 912.140 ;
        RECT -9.980 909.130 -6.980 909.140 ;
        RECT 2926.600 909.130 2929.600 909.140 ;
        RECT -9.980 732.140 -6.980 732.150 ;
        RECT 2926.600 732.140 2929.600 732.150 ;
        RECT -14.680 729.140 0.300 732.140 ;
        RECT 2919.700 729.140 2934.300 732.140 ;
        RECT -9.980 729.130 -6.980 729.140 ;
        RECT 2926.600 729.130 2929.600 729.140 ;
        RECT -9.980 552.140 -6.980 552.150 ;
        RECT 2926.600 552.140 2929.600 552.150 ;
        RECT -14.680 549.140 0.300 552.140 ;
        RECT 2919.700 549.140 2934.300 552.140 ;
        RECT -9.980 549.130 -6.980 549.140 ;
        RECT 2926.600 549.130 2929.600 549.140 ;
        RECT -9.980 372.140 -6.980 372.150 ;
        RECT 2926.600 372.140 2929.600 372.150 ;
        RECT -14.680 369.140 0.300 372.140 ;
        RECT 2919.700 369.140 2934.300 372.140 ;
        RECT -9.980 369.130 -6.980 369.140 ;
        RECT 2926.600 369.130 2929.600 369.140 ;
        RECT -9.980 192.140 -6.980 192.150 ;
        RECT 2926.600 192.140 2929.600 192.150 ;
        RECT -14.680 189.140 0.300 192.140 ;
        RECT 2919.700 189.140 2934.300 192.140 ;
        RECT -9.980 189.130 -6.980 189.140 ;
        RECT 2926.600 189.130 2929.600 189.140 ;
        RECT -9.980 12.140 -6.980 12.150 ;
        RECT 2926.600 12.140 2929.600 12.150 ;
        RECT -14.680 9.140 0.300 12.140 ;
        RECT 2919.700 9.140 2934.300 12.140 ;
        RECT -9.980 9.130 -6.980 9.140 ;
        RECT 2926.600 9.130 2929.600 9.140 ;
=======
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
>>>>>>> Latest run - not LVS matched yet
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 3519.700 97.020 3529.000 ;
        RECT 274.020 3519.700 277.020 3529.000 ;
        RECT 454.020 3519.700 457.020 3529.000 ;
        RECT 634.020 3519.700 637.020 3529.000 ;
        RECT 814.020 3519.700 817.020 3529.000 ;
        RECT 994.020 3519.700 997.020 3529.000 ;
        RECT 1174.020 3519.700 1177.020 3529.000 ;
        RECT 1354.020 3519.700 1357.020 3529.000 ;
        RECT 1534.020 3519.700 1537.020 3529.000 ;
        RECT 1714.020 3519.700 1717.020 3529.000 ;
        RECT 1894.020 3519.700 1897.020 3529.000 ;
        RECT 2074.020 3519.700 2077.020 3529.000 ;
        RECT 2254.020 3519.700 2257.020 3529.000 ;
        RECT 2434.020 3519.700 2437.020 3529.000 ;
        RECT 2614.020 3519.700 2617.020 3529.000 ;
        RECT 2794.020 3519.700 2797.020 3529.000 ;
        RECT 94.020 -9.320 97.020 0.300 ;
        RECT 274.020 -9.320 277.020 0.300 ;
        RECT 454.020 -9.320 457.020 0.300 ;
        RECT 634.020 -9.320 637.020 0.300 ;
        RECT 814.020 -9.320 817.020 0.300 ;
        RECT 994.020 -9.320 997.020 0.300 ;
        RECT 1174.020 -9.320 1177.020 0.300 ;
        RECT 1354.020 -9.320 1357.020 0.300 ;
        RECT 1534.020 -9.320 1537.020 0.300 ;
        RECT 1714.020 -9.320 1717.020 0.300 ;
        RECT 1894.020 -9.320 1897.020 0.300 ;
        RECT 2074.020 -9.320 2077.020 0.300 ;
        RECT 2254.020 -9.320 2257.020 0.300 ;
        RECT 2434.020 -9.320 2437.020 0.300 ;
        RECT 2614.020 -9.320 2617.020 0.300 ;
        RECT 2794.020 -9.320 2797.020 0.300 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT -13.770 3340.850 -12.590 3342.030 ;
        RECT -13.770 3339.250 -12.590 3340.430 ;
        RECT -13.770 3160.850 -12.590 3162.030 ;
        RECT -13.770 3159.250 -12.590 3160.430 ;
        RECT -13.770 2980.850 -12.590 2982.030 ;
        RECT -13.770 2979.250 -12.590 2980.430 ;
        RECT -13.770 2800.850 -12.590 2802.030 ;
        RECT -13.770 2799.250 -12.590 2800.430 ;
        RECT -13.770 2620.850 -12.590 2622.030 ;
        RECT -13.770 2619.250 -12.590 2620.430 ;
        RECT -13.770 2440.850 -12.590 2442.030 ;
        RECT -13.770 2439.250 -12.590 2440.430 ;
        RECT -13.770 2260.850 -12.590 2262.030 ;
        RECT -13.770 2259.250 -12.590 2260.430 ;
        RECT -13.770 2080.850 -12.590 2082.030 ;
        RECT -13.770 2079.250 -12.590 2080.430 ;
        RECT -13.770 1900.850 -12.590 1902.030 ;
        RECT -13.770 1899.250 -12.590 1900.430 ;
        RECT -13.770 1720.850 -12.590 1722.030 ;
        RECT -13.770 1719.250 -12.590 1720.430 ;
        RECT -13.770 1540.850 -12.590 1542.030 ;
        RECT -13.770 1539.250 -12.590 1540.430 ;
        RECT -13.770 1360.850 -12.590 1362.030 ;
        RECT -13.770 1359.250 -12.590 1360.430 ;
        RECT -13.770 1180.850 -12.590 1182.030 ;
        RECT -13.770 1179.250 -12.590 1180.430 ;
        RECT -13.770 1000.850 -12.590 1002.030 ;
        RECT -13.770 999.250 -12.590 1000.430 ;
        RECT -13.770 820.850 -12.590 822.030 ;
        RECT -13.770 819.250 -12.590 820.430 ;
        RECT -13.770 640.850 -12.590 642.030 ;
        RECT -13.770 639.250 -12.590 640.430 ;
        RECT -13.770 460.850 -12.590 462.030 ;
        RECT -13.770 459.250 -12.590 460.430 ;
        RECT -13.770 280.850 -12.590 282.030 ;
        RECT -13.770 279.250 -12.590 280.430 ;
        RECT -13.770 100.850 -12.590 102.030 ;
        RECT -13.770 99.250 -12.590 100.430 ;
        RECT 2932.210 3340.850 2933.390 3342.030 ;
        RECT 2932.210 3339.250 2933.390 3340.430 ;
        RECT 2932.210 3160.850 2933.390 3162.030 ;
        RECT 2932.210 3159.250 2933.390 3160.430 ;
        RECT 2932.210 2980.850 2933.390 2982.030 ;
        RECT 2932.210 2979.250 2933.390 2980.430 ;
        RECT 2932.210 2800.850 2933.390 2802.030 ;
        RECT 2932.210 2799.250 2933.390 2800.430 ;
        RECT 2932.210 2620.850 2933.390 2622.030 ;
        RECT 2932.210 2619.250 2933.390 2620.430 ;
        RECT 2932.210 2440.850 2933.390 2442.030 ;
        RECT 2932.210 2439.250 2933.390 2440.430 ;
        RECT 2932.210 2260.850 2933.390 2262.030 ;
        RECT 2932.210 2259.250 2933.390 2260.430 ;
        RECT 2932.210 2080.850 2933.390 2082.030 ;
        RECT 2932.210 2079.250 2933.390 2080.430 ;
        RECT 2932.210 1900.850 2933.390 1902.030 ;
        RECT 2932.210 1899.250 2933.390 1900.430 ;
        RECT 2932.210 1720.850 2933.390 1722.030 ;
        RECT 2932.210 1719.250 2933.390 1720.430 ;
        RECT 2932.210 1540.850 2933.390 1542.030 ;
        RECT 2932.210 1539.250 2933.390 1540.430 ;
        RECT 2932.210 1360.850 2933.390 1362.030 ;
        RECT 2932.210 1359.250 2933.390 1360.430 ;
        RECT 2932.210 1180.850 2933.390 1182.030 ;
        RECT 2932.210 1179.250 2933.390 1180.430 ;
        RECT 2932.210 1000.850 2933.390 1002.030 ;
        RECT 2932.210 999.250 2933.390 1000.430 ;
        RECT 2932.210 820.850 2933.390 822.030 ;
        RECT 2932.210 819.250 2933.390 820.430 ;
        RECT 2932.210 640.850 2933.390 642.030 ;
        RECT 2932.210 639.250 2933.390 640.430 ;
        RECT 2932.210 460.850 2933.390 462.030 ;
        RECT 2932.210 459.250 2933.390 460.430 ;
        RECT 2932.210 280.850 2933.390 282.030 ;
        RECT 2932.210 279.250 2933.390 280.430 ;
        RECT 2932.210 100.850 2933.390 102.030 ;
        RECT 2932.210 99.250 2933.390 100.430 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.140 -11.680 3342.150 ;
        RECT 2931.300 3342.140 2934.300 3342.150 ;
        RECT -14.680 3339.140 0.300 3342.140 ;
        RECT 2919.700 3339.140 2934.300 3342.140 ;
        RECT -14.680 3339.130 -11.680 3339.140 ;
        RECT 2931.300 3339.130 2934.300 3339.140 ;
        RECT -14.680 3162.140 -11.680 3162.150 ;
        RECT 2931.300 3162.140 2934.300 3162.150 ;
        RECT -14.680 3159.140 0.300 3162.140 ;
        RECT 2919.700 3159.140 2934.300 3162.140 ;
        RECT -14.680 3159.130 -11.680 3159.140 ;
        RECT 2931.300 3159.130 2934.300 3159.140 ;
        RECT -14.680 2982.140 -11.680 2982.150 ;
        RECT 2931.300 2982.140 2934.300 2982.150 ;
        RECT -14.680 2979.140 0.300 2982.140 ;
        RECT 2919.700 2979.140 2934.300 2982.140 ;
        RECT -14.680 2979.130 -11.680 2979.140 ;
        RECT 2931.300 2979.130 2934.300 2979.140 ;
        RECT -14.680 2802.140 -11.680 2802.150 ;
        RECT 2931.300 2802.140 2934.300 2802.150 ;
        RECT -14.680 2799.140 0.300 2802.140 ;
        RECT 2919.700 2799.140 2934.300 2802.140 ;
        RECT -14.680 2799.130 -11.680 2799.140 ;
        RECT 2931.300 2799.130 2934.300 2799.140 ;
        RECT -14.680 2622.140 -11.680 2622.150 ;
        RECT 2931.300 2622.140 2934.300 2622.150 ;
        RECT -14.680 2619.140 0.300 2622.140 ;
        RECT 2919.700 2619.140 2934.300 2622.140 ;
        RECT -14.680 2619.130 -11.680 2619.140 ;
        RECT 2931.300 2619.130 2934.300 2619.140 ;
        RECT -14.680 2442.140 -11.680 2442.150 ;
        RECT 2931.300 2442.140 2934.300 2442.150 ;
        RECT -14.680 2439.140 0.300 2442.140 ;
        RECT 2919.700 2439.140 2934.300 2442.140 ;
        RECT -14.680 2439.130 -11.680 2439.140 ;
        RECT 2931.300 2439.130 2934.300 2439.140 ;
        RECT -14.680 2262.140 -11.680 2262.150 ;
        RECT 2931.300 2262.140 2934.300 2262.150 ;
        RECT -14.680 2259.140 0.300 2262.140 ;
        RECT 2919.700 2259.140 2934.300 2262.140 ;
        RECT -14.680 2259.130 -11.680 2259.140 ;
        RECT 2931.300 2259.130 2934.300 2259.140 ;
        RECT -14.680 2082.140 -11.680 2082.150 ;
        RECT 2931.300 2082.140 2934.300 2082.150 ;
        RECT -14.680 2079.140 0.300 2082.140 ;
        RECT 2919.700 2079.140 2934.300 2082.140 ;
        RECT -14.680 2079.130 -11.680 2079.140 ;
        RECT 2931.300 2079.130 2934.300 2079.140 ;
        RECT -14.680 1902.140 -11.680 1902.150 ;
        RECT 2931.300 1902.140 2934.300 1902.150 ;
        RECT -14.680 1899.140 0.300 1902.140 ;
        RECT 2919.700 1899.140 2934.300 1902.140 ;
        RECT -14.680 1899.130 -11.680 1899.140 ;
        RECT 2931.300 1899.130 2934.300 1899.140 ;
        RECT -14.680 1722.140 -11.680 1722.150 ;
        RECT 2931.300 1722.140 2934.300 1722.150 ;
        RECT -14.680 1719.140 0.300 1722.140 ;
        RECT 2919.700 1719.140 2934.300 1722.140 ;
        RECT -14.680 1719.130 -11.680 1719.140 ;
        RECT 2931.300 1719.130 2934.300 1719.140 ;
        RECT -14.680 1542.140 -11.680 1542.150 ;
        RECT 2931.300 1542.140 2934.300 1542.150 ;
        RECT -14.680 1539.140 0.300 1542.140 ;
        RECT 2919.700 1539.140 2934.300 1542.140 ;
        RECT -14.680 1539.130 -11.680 1539.140 ;
        RECT 2931.300 1539.130 2934.300 1539.140 ;
        RECT -14.680 1362.140 -11.680 1362.150 ;
        RECT 2931.300 1362.140 2934.300 1362.150 ;
        RECT -14.680 1359.140 0.300 1362.140 ;
        RECT 2919.700 1359.140 2934.300 1362.140 ;
        RECT -14.680 1359.130 -11.680 1359.140 ;
        RECT 2931.300 1359.130 2934.300 1359.140 ;
        RECT -14.680 1182.140 -11.680 1182.150 ;
        RECT 2931.300 1182.140 2934.300 1182.150 ;
        RECT -14.680 1179.140 0.300 1182.140 ;
        RECT 2919.700 1179.140 2934.300 1182.140 ;
        RECT -14.680 1179.130 -11.680 1179.140 ;
        RECT 2931.300 1179.130 2934.300 1179.140 ;
        RECT -14.680 1002.140 -11.680 1002.150 ;
        RECT 2931.300 1002.140 2934.300 1002.150 ;
        RECT -14.680 999.140 0.300 1002.140 ;
        RECT 2919.700 999.140 2934.300 1002.140 ;
        RECT -14.680 999.130 -11.680 999.140 ;
        RECT 2931.300 999.130 2934.300 999.140 ;
        RECT -14.680 822.140 -11.680 822.150 ;
        RECT 2931.300 822.140 2934.300 822.150 ;
        RECT -14.680 819.140 0.300 822.140 ;
        RECT 2919.700 819.140 2934.300 822.140 ;
        RECT -14.680 819.130 -11.680 819.140 ;
        RECT 2931.300 819.130 2934.300 819.140 ;
        RECT -14.680 642.140 -11.680 642.150 ;
        RECT 2931.300 642.140 2934.300 642.150 ;
        RECT -14.680 639.140 0.300 642.140 ;
        RECT 2919.700 639.140 2934.300 642.140 ;
        RECT -14.680 639.130 -11.680 639.140 ;
        RECT 2931.300 639.130 2934.300 639.140 ;
        RECT -14.680 462.140 -11.680 462.150 ;
        RECT 2931.300 462.140 2934.300 462.150 ;
        RECT -14.680 459.140 0.300 462.140 ;
        RECT 2919.700 459.140 2934.300 462.140 ;
        RECT -14.680 459.130 -11.680 459.140 ;
        RECT 2931.300 459.130 2934.300 459.140 ;
        RECT -14.680 282.140 -11.680 282.150 ;
        RECT 2931.300 282.140 2934.300 282.150 ;
        RECT -14.680 279.140 0.300 282.140 ;
        RECT 2919.700 279.140 2934.300 282.140 ;
        RECT -14.680 279.130 -11.680 279.140 ;
        RECT 2931.300 279.130 2934.300 279.140 ;
        RECT -14.680 102.140 -11.680 102.150 ;
        RECT 2931.300 102.140 2934.300 102.150 ;
        RECT -14.680 99.140 0.300 102.140 ;
        RECT 2919.700 99.140 2934.300 102.140 ;
        RECT -14.680 99.130 -11.680 99.140 ;
        RECT 2931.300 99.130 2934.300 99.140 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
=======
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 -9.220 457.020 3528.900 ;
        RECT 634.020 -9.220 637.020 3528.900 ;
        RECT 814.020 -9.220 817.020 3528.900 ;
        RECT 994.020 -9.220 997.020 3528.900 ;
        RECT 1174.020 -9.220 1177.020 3528.900 ;
        RECT 1354.020 -9.220 1357.020 3528.900 ;
        RECT 1534.020 -9.220 1537.020 3528.900 ;
        RECT 1714.020 -9.220 1717.020 3528.900 ;
        RECT 1894.020 -9.220 1897.020 3528.900 ;
        RECT 2074.020 -9.220 2077.020 3528.900 ;
        RECT 2254.020 -9.220 2257.020 3528.900 ;
        RECT 2434.020 -9.220 2437.020 3528.900 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 3519.700 25.020 3538.400 ;
        RECT 202.020 3519.700 205.020 3538.400 ;
        RECT 382.020 3519.700 385.020 3538.400 ;
        RECT 562.020 3519.700 565.020 3538.400 ;
        RECT 742.020 3519.700 745.020 3538.400 ;
        RECT 922.020 3519.700 925.020 3538.400 ;
        RECT 1102.020 3519.700 1105.020 3538.400 ;
        RECT 1282.020 3519.700 1285.020 3538.400 ;
        RECT 1462.020 3519.700 1465.020 3538.400 ;
        RECT 1642.020 3519.700 1645.020 3538.400 ;
        RECT 1822.020 3519.700 1825.020 3538.400 ;
        RECT 2002.020 3519.700 2005.020 3538.400 ;
        RECT 2182.020 3519.700 2185.020 3538.400 ;
        RECT 2362.020 3519.700 2365.020 3538.400 ;
        RECT 2542.020 3519.700 2545.020 3538.400 ;
        RECT 2722.020 3519.700 2725.020 3538.400 ;
        RECT 2902.020 3519.700 2905.020 3538.400 ;
        RECT 22.020 -18.720 25.020 0.300 ;
        RECT 202.020 -18.720 205.020 0.300 ;
        RECT 382.020 -18.720 385.020 0.300 ;
        RECT 562.020 -18.720 565.020 0.300 ;
        RECT 742.020 -18.720 745.020 0.300 ;
        RECT 922.020 -18.720 925.020 0.300 ;
        RECT 1102.020 -18.720 1105.020 0.300 ;
        RECT 1282.020 -18.720 1285.020 0.300 ;
        RECT 1462.020 -18.720 1465.020 0.300 ;
        RECT 1642.020 -18.720 1645.020 0.300 ;
        RECT 1822.020 -18.720 1825.020 0.300 ;
        RECT 2002.020 -18.720 2005.020 0.300 ;
        RECT 2182.020 -18.720 2185.020 0.300 ;
        RECT 2362.020 -18.720 2365.020 0.300 ;
        RECT 2542.020 -18.720 2545.020 0.300 ;
        RECT 2722.020 -18.720 2725.020 0.300 ;
        RECT 2902.020 -18.720 2905.020 0.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 0.300 3450.380 ;
        RECT 2919.700 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 0.300 3270.380 ;
        RECT 2919.700 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 0.300 3090.380 ;
        RECT 2919.700 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 0.300 2910.380 ;
        RECT 2919.700 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 0.300 2730.380 ;
        RECT 2919.700 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 0.300 2550.380 ;
        RECT 2919.700 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 0.300 2370.380 ;
        RECT 2919.700 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 0.300 2190.380 ;
        RECT 2919.700 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 0.300 2010.380 ;
        RECT 2919.700 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 0.300 1830.380 ;
        RECT 2919.700 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 0.300 1650.380 ;
        RECT 2919.700 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 0.300 1470.380 ;
        RECT 2919.700 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 0.300 1290.380 ;
        RECT 2919.700 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 0.300 1110.380 ;
        RECT 2919.700 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 0.300 930.380 ;
        RECT 2919.700 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 0.300 750.380 ;
        RECT 2919.700 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 0.300 570.380 ;
        RECT 2919.700 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 0.300 390.380 ;
        RECT 2919.700 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 0.300 210.380 ;
        RECT 2919.700 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 0.300 30.380 ;
        RECT 2919.700 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
=======
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 -18.420 565.020 3538.100 ;
        RECT 742.020 -18.420 745.020 3538.100 ;
        RECT 922.020 -18.420 925.020 3538.100 ;
        RECT 1102.020 -18.420 1105.020 3538.100 ;
        RECT 1282.020 -18.420 1285.020 3538.100 ;
        RECT 1462.020 -18.420 1465.020 3538.100 ;
        RECT 1642.020 -18.420 1645.020 3538.100 ;
        RECT 1822.020 -18.420 1825.020 3538.100 ;
        RECT 2002.020 -18.420 2005.020 3538.100 ;
        RECT 2182.020 -18.420 2185.020 3538.100 ;
        RECT 2362.020 -18.420 2365.020 3538.100 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 3519.700 115.020 3538.400 ;
        RECT 292.020 3519.700 295.020 3538.400 ;
        RECT 472.020 3519.700 475.020 3538.400 ;
        RECT 652.020 3519.700 655.020 3538.400 ;
        RECT 832.020 3519.700 835.020 3538.400 ;
        RECT 1012.020 3519.700 1015.020 3538.400 ;
        RECT 1192.020 3519.700 1195.020 3538.400 ;
        RECT 1372.020 3519.700 1375.020 3538.400 ;
        RECT 1552.020 3519.700 1555.020 3538.400 ;
        RECT 1732.020 3519.700 1735.020 3538.400 ;
        RECT 1912.020 3519.700 1915.020 3538.400 ;
        RECT 2092.020 3519.700 2095.020 3538.400 ;
        RECT 2272.020 3519.700 2275.020 3538.400 ;
        RECT 2452.020 3519.700 2455.020 3538.400 ;
        RECT 2632.020 3519.700 2635.020 3538.400 ;
        RECT 2812.020 3519.700 2815.020 3538.400 ;
        RECT 112.020 -18.720 115.020 0.300 ;
        RECT 292.020 -18.720 295.020 0.300 ;
        RECT 472.020 -18.720 475.020 0.300 ;
        RECT 652.020 -18.720 655.020 0.300 ;
        RECT 832.020 -18.720 835.020 0.300 ;
        RECT 1012.020 -18.720 1015.020 0.300 ;
        RECT 1192.020 -18.720 1195.020 0.300 ;
        RECT 1372.020 -18.720 1375.020 0.300 ;
        RECT 1552.020 -18.720 1555.020 0.300 ;
        RECT 1732.020 -18.720 1735.020 0.300 ;
        RECT 1912.020 -18.720 1915.020 0.300 ;
        RECT 2092.020 -18.720 2095.020 0.300 ;
        RECT 2272.020 -18.720 2275.020 0.300 ;
        RECT 2452.020 -18.720 2455.020 0.300 ;
        RECT 2632.020 -18.720 2635.020 0.300 ;
        RECT 2812.020 -18.720 2815.020 0.300 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 0.300 3360.380 ;
        RECT 2919.700 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 0.300 3180.380 ;
        RECT 2919.700 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 0.300 3000.380 ;
        RECT 2919.700 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 0.300 2820.380 ;
        RECT 2919.700 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 0.300 2640.380 ;
        RECT 2919.700 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 0.300 2460.380 ;
        RECT 2919.700 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 0.300 2280.380 ;
        RECT 2919.700 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 0.300 2100.380 ;
        RECT 2919.700 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 0.300 1920.380 ;
        RECT 2919.700 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 0.300 1740.380 ;
        RECT 2919.700 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 0.300 1560.380 ;
        RECT 2919.700 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 0.300 1380.380 ;
        RECT 2919.700 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 0.300 1200.380 ;
        RECT 2919.700 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 0.300 1020.380 ;
        RECT 2919.700 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 0.300 840.380 ;
        RECT 2919.700 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 0.300 660.380 ;
        RECT 2919.700 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 0.300 480.380 ;
        RECT 2919.700 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 0.300 300.380 ;
        RECT 2919.700 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 0.300 120.380 ;
        RECT 2919.700 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
=======
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 -18.420 475.020 3538.100 ;
        RECT 652.020 -18.420 655.020 3538.100 ;
        RECT 832.020 -18.420 835.020 3538.100 ;
        RECT 1012.020 -18.420 1015.020 3538.100 ;
        RECT 1192.020 -18.420 1195.020 3538.100 ;
        RECT 1372.020 -18.420 1375.020 3538.100 ;
        RECT 1552.020 -18.420 1555.020 3538.100 ;
        RECT 1732.020 -18.420 1735.020 3538.100 ;
        RECT 1912.020 -18.420 1915.020 3538.100 ;
        RECT 2092.020 -18.420 2095.020 3538.100 ;
        RECT 2272.020 -18.420 2275.020 3538.100 ;
        RECT 2452.020 -18.420 2455.020 3538.100 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 3519.700 43.020 3547.800 ;
        RECT 220.020 3519.700 223.020 3547.800 ;
        RECT 400.020 3519.700 403.020 3547.800 ;
        RECT 580.020 3519.700 583.020 3547.800 ;
        RECT 760.020 3519.700 763.020 3547.800 ;
        RECT 940.020 3519.700 943.020 3547.800 ;
        RECT 1120.020 3519.700 1123.020 3547.800 ;
        RECT 1300.020 3519.700 1303.020 3547.800 ;
        RECT 1480.020 3519.700 1483.020 3547.800 ;
        RECT 1660.020 3519.700 1663.020 3547.800 ;
        RECT 1840.020 3519.700 1843.020 3547.800 ;
        RECT 2020.020 3519.700 2023.020 3547.800 ;
        RECT 2200.020 3519.700 2203.020 3547.800 ;
        RECT 2380.020 3519.700 2383.020 3547.800 ;
        RECT 2560.020 3519.700 2563.020 3547.800 ;
        RECT 2740.020 3519.700 2743.020 3547.800 ;
        RECT 40.020 -28.120 43.020 0.300 ;
        RECT 220.020 -28.120 223.020 0.300 ;
        RECT 400.020 -28.120 403.020 0.300 ;
        RECT 580.020 -28.120 583.020 0.300 ;
        RECT 760.020 -28.120 763.020 0.300 ;
        RECT 940.020 -28.120 943.020 0.300 ;
        RECT 1120.020 -28.120 1123.020 0.300 ;
        RECT 1300.020 -28.120 1303.020 0.300 ;
        RECT 1480.020 -28.120 1483.020 0.300 ;
        RECT 1660.020 -28.120 1663.020 0.300 ;
        RECT 1840.020 -28.120 1843.020 0.300 ;
        RECT 2020.020 -28.120 2023.020 0.300 ;
        RECT 2200.020 -28.120 2203.020 0.300 ;
        RECT 2380.020 -28.120 2383.020 0.300 ;
        RECT 2560.020 -28.120 2563.020 0.300 ;
        RECT 2740.020 -28.120 2743.020 0.300 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 0.300 3468.380 ;
        RECT 2919.700 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 0.300 3288.380 ;
        RECT 2919.700 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 0.300 3108.380 ;
        RECT 2919.700 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 0.300 2928.380 ;
        RECT 2919.700 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 0.300 2748.380 ;
        RECT 2919.700 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 0.300 2568.380 ;
        RECT 2919.700 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 0.300 2388.380 ;
        RECT 2919.700 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 0.300 2208.380 ;
        RECT 2919.700 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 0.300 2028.380 ;
        RECT 2919.700 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 0.300 1848.380 ;
        RECT 2919.700 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 0.300 1668.380 ;
        RECT 2919.700 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 0.300 1488.380 ;
        RECT 2919.700 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 0.300 1308.380 ;
        RECT 2919.700 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 0.300 1128.380 ;
        RECT 2919.700 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 0.300 948.380 ;
        RECT 2919.700 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 0.300 768.380 ;
        RECT 2919.700 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 0.300 588.380 ;
        RECT 2919.700 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 0.300 408.380 ;
        RECT 2919.700 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 0.300 228.380 ;
        RECT 2919.700 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 0.300 48.380 ;
        RECT 2919.700 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
=======
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 -27.620 583.020 3547.300 ;
        RECT 760.020 -27.620 763.020 3547.300 ;
        RECT 940.020 -27.620 943.020 3547.300 ;
        RECT 1120.020 -27.620 1123.020 3547.300 ;
        RECT 1300.020 -27.620 1303.020 3547.300 ;
        RECT 1480.020 -27.620 1483.020 3547.300 ;
        RECT 1660.020 -27.620 1663.020 3547.300 ;
        RECT 1840.020 -27.620 1843.020 3547.300 ;
        RECT 2020.020 -27.620 2023.020 3547.300 ;
        RECT 2200.020 -27.620 2203.020 3547.300 ;
        RECT 2380.020 -27.620 2383.020 3547.300 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 3519.700 133.020 3547.800 ;
        RECT 310.020 3519.700 313.020 3547.800 ;
        RECT 490.020 3519.700 493.020 3547.800 ;
        RECT 670.020 3519.700 673.020 3547.800 ;
        RECT 850.020 3519.700 853.020 3547.800 ;
        RECT 1030.020 3519.700 1033.020 3547.800 ;
        RECT 1210.020 3519.700 1213.020 3547.800 ;
        RECT 1390.020 3519.700 1393.020 3547.800 ;
        RECT 1570.020 3519.700 1573.020 3547.800 ;
        RECT 1750.020 3519.700 1753.020 3547.800 ;
        RECT 1930.020 3519.700 1933.020 3547.800 ;
        RECT 2110.020 3519.700 2113.020 3547.800 ;
        RECT 2290.020 3519.700 2293.020 3547.800 ;
        RECT 2470.020 3519.700 2473.020 3547.800 ;
        RECT 2650.020 3519.700 2653.020 3547.800 ;
        RECT 2830.020 3519.700 2833.020 3547.800 ;
        RECT 130.020 -28.120 133.020 0.300 ;
        RECT 310.020 -28.120 313.020 0.300 ;
        RECT 490.020 -28.120 493.020 0.300 ;
        RECT 670.020 -28.120 673.020 0.300 ;
        RECT 850.020 -28.120 853.020 0.300 ;
        RECT 1030.020 -28.120 1033.020 0.300 ;
        RECT 1210.020 -28.120 1213.020 0.300 ;
        RECT 1390.020 -28.120 1393.020 0.300 ;
        RECT 1570.020 -28.120 1573.020 0.300 ;
        RECT 1750.020 -28.120 1753.020 0.300 ;
        RECT 1930.020 -28.120 1933.020 0.300 ;
        RECT 2110.020 -28.120 2113.020 0.300 ;
        RECT 2290.020 -28.120 2293.020 0.300 ;
        RECT 2470.020 -28.120 2473.020 0.300 ;
        RECT 2650.020 -28.120 2653.020 0.300 ;
        RECT 2830.020 -28.120 2833.020 0.300 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 0.300 3378.380 ;
        RECT 2919.700 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 0.300 3198.380 ;
        RECT 2919.700 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 0.300 3018.380 ;
        RECT 2919.700 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 0.300 2838.380 ;
        RECT 2919.700 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 0.300 2658.380 ;
        RECT 2919.700 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 0.300 2478.380 ;
        RECT 2919.700 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 0.300 2298.380 ;
        RECT 2919.700 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 0.300 2118.380 ;
        RECT 2919.700 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 0.300 1938.380 ;
        RECT 2919.700 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 0.300 1758.380 ;
        RECT 2919.700 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 0.300 1578.380 ;
        RECT 2919.700 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 0.300 1398.380 ;
        RECT 2919.700 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 0.300 1218.380 ;
        RECT 2919.700 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 0.300 1038.380 ;
        RECT 2919.700 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 0.300 858.380 ;
        RECT 2919.700 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 0.300 678.380 ;
        RECT 2919.700 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 0.300 498.380 ;
        RECT 2919.700 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 0.300 318.380 ;
        RECT 2919.700 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 0.300 138.380 ;
        RECT 2919.700 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 3519.700 61.020 3557.200 ;
        RECT 238.020 3519.700 241.020 3557.200 ;
        RECT 418.020 3519.700 421.020 3557.200 ;
        RECT 598.020 3519.700 601.020 3557.200 ;
        RECT 778.020 3519.700 781.020 3557.200 ;
        RECT 958.020 3519.700 961.020 3557.200 ;
        RECT 1138.020 3519.700 1141.020 3557.200 ;
        RECT 1318.020 3519.700 1321.020 3557.200 ;
        RECT 1498.020 3519.700 1501.020 3557.200 ;
        RECT 1678.020 3519.700 1681.020 3557.200 ;
        RECT 1858.020 3519.700 1861.020 3557.200 ;
        RECT 2038.020 3519.700 2041.020 3557.200 ;
        RECT 2218.020 3519.700 2221.020 3557.200 ;
        RECT 2398.020 3519.700 2401.020 3557.200 ;
        RECT 2578.020 3519.700 2581.020 3557.200 ;
        RECT 2758.020 3519.700 2761.020 3557.200 ;
        RECT 58.020 -37.520 61.020 0.300 ;
        RECT 238.020 -37.520 241.020 0.300 ;
        RECT 418.020 -37.520 421.020 0.300 ;
        RECT 598.020 -37.520 601.020 0.300 ;
        RECT 778.020 -37.520 781.020 0.300 ;
        RECT 958.020 -37.520 961.020 0.300 ;
        RECT 1138.020 -37.520 1141.020 0.300 ;
        RECT 1318.020 -37.520 1321.020 0.300 ;
        RECT 1498.020 -37.520 1501.020 0.300 ;
        RECT 1678.020 -37.520 1681.020 0.300 ;
        RECT 1858.020 -37.520 1861.020 0.300 ;
        RECT 2038.020 -37.520 2041.020 0.300 ;
        RECT 2218.020 -37.520 2221.020 0.300 ;
        RECT 2398.020 -37.520 2401.020 0.300 ;
        RECT 2578.020 -37.520 2581.020 0.300 ;
        RECT 2758.020 -37.520 2761.020 0.300 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 0.300 3486.380 ;
        RECT 2919.700 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 0.300 3306.380 ;
        RECT 2919.700 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 0.300 3126.380 ;
        RECT 2919.700 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 0.300 2946.380 ;
        RECT 2919.700 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 0.300 2766.380 ;
        RECT 2919.700 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 0.300 2586.380 ;
        RECT 2919.700 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 0.300 2406.380 ;
        RECT 2919.700 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 0.300 2226.380 ;
        RECT 2919.700 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 0.300 2046.380 ;
        RECT 2919.700 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 0.300 1866.380 ;
        RECT 2919.700 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 0.300 1686.380 ;
        RECT 2919.700 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 0.300 1506.380 ;
        RECT 2919.700 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 0.300 1326.380 ;
        RECT 2919.700 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 0.300 1146.380 ;
        RECT 2919.700 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 0.300 966.380 ;
        RECT 2919.700 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 0.300 786.380 ;
        RECT 2919.700 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 0.300 606.380 ;
        RECT 2919.700 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 0.300 426.380 ;
        RECT 2919.700 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 0.300 246.380 ;
        RECT 2919.700 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 0.300 66.380 ;
        RECT 2919.700 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
=======
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 -27.620 493.020 3547.300 ;
        RECT 670.020 -27.620 673.020 3547.300 ;
        RECT 850.020 -27.620 853.020 3547.300 ;
        RECT 1030.020 -27.620 1033.020 3547.300 ;
        RECT 1210.020 -27.620 1213.020 3547.300 ;
        RECT 1390.020 -27.620 1393.020 3547.300 ;
        RECT 1570.020 -27.620 1573.020 3547.300 ;
        RECT 1750.020 -27.620 1753.020 3547.300 ;
        RECT 1930.020 -27.620 1933.020 3547.300 ;
        RECT 2110.020 -27.620 2113.020 3547.300 ;
        RECT 2290.020 -27.620 2293.020 3547.300 ;
        RECT 2470.020 -27.620 2473.020 3547.300 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 -36.820 421.020 3556.500 ;
        RECT 598.020 -36.820 601.020 3556.500 ;
        RECT 778.020 -36.820 781.020 3556.500 ;
        RECT 958.020 -36.820 961.020 3556.500 ;
        RECT 1138.020 -36.820 1141.020 3556.500 ;
        RECT 1318.020 -36.820 1321.020 3556.500 ;
        RECT 1498.020 -36.820 1501.020 3556.500 ;
        RECT 1678.020 -36.820 1681.020 3556.500 ;
        RECT 1858.020 -36.820 1861.020 3556.500 ;
        RECT 2038.020 -36.820 2041.020 3556.500 ;
        RECT 2218.020 -36.820 2221.020 3556.500 ;
        RECT 2398.020 -36.820 2401.020 3556.500 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 3519.700 151.020 3557.200 ;
        RECT 328.020 3519.700 331.020 3557.200 ;
        RECT 508.020 3519.700 511.020 3557.200 ;
        RECT 688.020 3519.700 691.020 3557.200 ;
        RECT 868.020 3519.700 871.020 3557.200 ;
        RECT 1048.020 3519.700 1051.020 3557.200 ;
        RECT 1228.020 3519.700 1231.020 3557.200 ;
        RECT 1408.020 3519.700 1411.020 3557.200 ;
        RECT 1588.020 3519.700 1591.020 3557.200 ;
        RECT 1768.020 3519.700 1771.020 3557.200 ;
        RECT 1948.020 3519.700 1951.020 3557.200 ;
        RECT 2128.020 3519.700 2131.020 3557.200 ;
        RECT 2308.020 3519.700 2311.020 3557.200 ;
        RECT 2488.020 3519.700 2491.020 3557.200 ;
        RECT 2668.020 3519.700 2671.020 3557.200 ;
        RECT 2848.020 3519.700 2851.020 3557.200 ;
        RECT 148.020 -37.520 151.020 0.300 ;
        RECT 328.020 -37.520 331.020 0.300 ;
        RECT 508.020 -37.520 511.020 0.300 ;
        RECT 688.020 -37.520 691.020 0.300 ;
        RECT 868.020 -37.520 871.020 0.300 ;
        RECT 1048.020 -37.520 1051.020 0.300 ;
        RECT 1228.020 -37.520 1231.020 0.300 ;
        RECT 1408.020 -37.520 1411.020 0.300 ;
        RECT 1588.020 -37.520 1591.020 0.300 ;
        RECT 1768.020 -37.520 1771.020 0.300 ;
        RECT 1948.020 -37.520 1951.020 0.300 ;
        RECT 2128.020 -37.520 2131.020 0.300 ;
        RECT 2308.020 -37.520 2311.020 0.300 ;
        RECT 2488.020 -37.520 2491.020 0.300 ;
        RECT 2668.020 -37.520 2671.020 0.300 ;
        RECT 2848.020 -37.520 2851.020 0.300 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 0.300 3396.380 ;
        RECT 2919.700 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 0.300 3216.380 ;
        RECT 2919.700 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 0.300 3036.380 ;
        RECT 2919.700 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 0.300 2856.380 ;
        RECT 2919.700 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 0.300 2676.380 ;
        RECT 2919.700 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 0.300 2496.380 ;
        RECT 2919.700 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 0.300 2316.380 ;
        RECT 2919.700 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 0.300 2136.380 ;
        RECT 2919.700 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 0.300 1956.380 ;
        RECT 2919.700 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 0.300 1776.380 ;
        RECT 2919.700 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 0.300 1596.380 ;
        RECT 2919.700 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 0.300 1416.380 ;
        RECT 2919.700 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 0.300 1236.380 ;
        RECT 2919.700 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 0.300 1056.380 ;
        RECT 2919.700 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 0.300 876.380 ;
        RECT 2919.700 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 0.300 696.380 ;
        RECT 2919.700 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 0.300 516.380 ;
        RECT 2919.700 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 0.300 336.380 ;
        RECT 2919.700 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 0.300 156.380 ;
        RECT 2919.700 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
=======
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 -36.820 511.020 3556.500 ;
        RECT 688.020 -36.820 691.020 3556.500 ;
        RECT 868.020 -36.820 871.020 3556.500 ;
        RECT 1048.020 -36.820 1051.020 3556.500 ;
        RECT 1228.020 -36.820 1231.020 3556.500 ;
        RECT 1408.020 -36.820 1411.020 3556.500 ;
        RECT 1588.020 -36.820 1591.020 3556.500 ;
        RECT 1768.020 -36.820 1771.020 3556.500 ;
        RECT 1948.020 -36.820 1951.020 3556.500 ;
        RECT 2128.020 -36.820 2131.020 3556.500 ;
        RECT 2308.020 -36.820 2311.020 3556.500 ;
        RECT 2488.020 -36.820 2491.020 3556.500 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
>>>>>>> Latest run - not LVS matched yet
    END
  END vssa2
  OBS
      LAYER li1 ;
<<<<<<< HEAD
        RECT 276.145 2.805 2799.415 3477.435 ;
      LAYER met1 ;
        RECT 2.830 2.760 2914.100 3512.160 ;
      LAYER met2 ;
        RECT 2.710 0.300 2917.370 3519.700 ;
      LAYER met3 ;
        RECT 0.300 10.715 2919.700 3508.965 ;
      LAYER met4 ;
        RECT 4.020 0.300 2905.020 3519.700 ;
      LAYER met5 ;
        RECT 0.300 9.130 2919.700 3486.390 ;
=======
        RECT 1155.520 1710.795 1944.420 2488.885 ;
      LAYER met1 ;
        RECT 1153.750 1708.200 1944.420 2489.040 ;
      LAYER met2 ;
        RECT 1150.550 2495.720 1153.030 2496.010 ;
        RECT 1153.870 2495.720 1159.470 2496.010 ;
        RECT 1160.310 2495.720 1165.910 2496.010 ;
        RECT 1166.750 2495.720 1172.350 2496.010 ;
        RECT 1173.190 2495.720 1178.790 2496.010 ;
        RECT 1179.630 2495.720 1185.230 2496.010 ;
        RECT 1186.070 2495.720 1191.670 2496.010 ;
        RECT 1192.510 2495.720 1198.110 2496.010 ;
        RECT 1198.950 2495.720 1204.550 2496.010 ;
        RECT 1205.390 2495.720 1210.990 2496.010 ;
        RECT 1211.830 2495.720 1217.430 2496.010 ;
        RECT 1218.270 2495.720 1223.870 2496.010 ;
        RECT 1224.710 2495.720 1230.310 2496.010 ;
        RECT 1231.150 2495.720 1236.750 2496.010 ;
        RECT 1237.590 2495.720 1243.190 2496.010 ;
        RECT 1244.030 2495.720 1249.630 2496.010 ;
        RECT 1250.470 2495.720 1256.070 2496.010 ;
        RECT 1256.910 2495.720 1262.510 2496.010 ;
        RECT 1263.350 2495.720 1268.950 2496.010 ;
        RECT 1269.790 2495.720 1275.390 2496.010 ;
        RECT 1276.230 2495.720 1281.830 2496.010 ;
        RECT 1282.670 2495.720 1288.270 2496.010 ;
        RECT 1289.110 2495.720 1294.710 2496.010 ;
        RECT 1295.550 2495.720 1301.150 2496.010 ;
        RECT 1301.990 2495.720 1307.590 2496.010 ;
        RECT 1308.430 2495.720 1314.030 2496.010 ;
        RECT 1314.870 2495.720 1320.470 2496.010 ;
        RECT 1321.310 2495.720 1326.910 2496.010 ;
        RECT 1327.750 2495.720 1333.350 2496.010 ;
        RECT 1334.190 2495.720 1339.790 2496.010 ;
        RECT 1340.630 2495.720 1346.230 2496.010 ;
        RECT 1347.070 2495.720 1352.670 2496.010 ;
        RECT 1353.510 2495.720 1359.110 2496.010 ;
        RECT 1359.950 2495.720 1365.550 2496.010 ;
        RECT 1366.390 2495.720 1371.990 2496.010 ;
        RECT 1372.830 2495.720 1378.430 2496.010 ;
        RECT 1379.270 2495.720 1384.870 2496.010 ;
        RECT 1385.710 2495.720 1391.310 2496.010 ;
        RECT 1392.150 2495.720 1397.750 2496.010 ;
        RECT 1398.590 2495.720 1404.190 2496.010 ;
        RECT 1405.030 2495.720 1410.630 2496.010 ;
        RECT 1411.470 2495.720 1417.070 2496.010 ;
        RECT 1417.910 2495.720 1423.970 2496.010 ;
        RECT 1424.810 2495.720 1430.410 2496.010 ;
        RECT 1431.250 2495.720 1436.850 2496.010 ;
        RECT 1437.690 2495.720 1443.290 2496.010 ;
        RECT 1444.130 2495.720 1449.730 2496.010 ;
        RECT 1450.570 2495.720 1456.170 2496.010 ;
        RECT 1457.010 2495.720 1462.610 2496.010 ;
        RECT 1463.450 2495.720 1469.050 2496.010 ;
        RECT 1469.890 2495.720 1475.490 2496.010 ;
        RECT 1476.330 2495.720 1481.930 2496.010 ;
        RECT 1482.770 2495.720 1488.370 2496.010 ;
        RECT 1489.210 2495.720 1494.810 2496.010 ;
        RECT 1495.650 2495.720 1501.250 2496.010 ;
        RECT 1502.090 2495.720 1507.690 2496.010 ;
        RECT 1508.530 2495.720 1514.130 2496.010 ;
        RECT 1514.970 2495.720 1520.570 2496.010 ;
        RECT 1521.410 2495.720 1527.010 2496.010 ;
        RECT 1527.850 2495.720 1533.450 2496.010 ;
        RECT 1534.290 2495.720 1539.890 2496.010 ;
        RECT 1540.730 2495.720 1546.330 2496.010 ;
        RECT 1547.170 2495.720 1552.770 2496.010 ;
        RECT 1553.610 2495.720 1559.210 2496.010 ;
        RECT 1560.050 2495.720 1565.650 2496.010 ;
        RECT 1566.490 2495.720 1572.090 2496.010 ;
        RECT 1572.930 2495.720 1578.530 2496.010 ;
        RECT 1579.370 2495.720 1584.970 2496.010 ;
        RECT 1585.810 2495.720 1591.410 2496.010 ;
        RECT 1592.250 2495.720 1597.850 2496.010 ;
        RECT 1598.690 2495.720 1604.290 2496.010 ;
        RECT 1605.130 2495.720 1610.730 2496.010 ;
        RECT 1611.570 2495.720 1617.170 2496.010 ;
        RECT 1618.010 2495.720 1623.610 2496.010 ;
        RECT 1624.450 2495.720 1630.050 2496.010 ;
        RECT 1630.890 2495.720 1636.490 2496.010 ;
        RECT 1637.330 2495.720 1642.930 2496.010 ;
        RECT 1643.770 2495.720 1649.370 2496.010 ;
        RECT 1650.210 2495.720 1655.810 2496.010 ;
        RECT 1656.650 2495.720 1662.250 2496.010 ;
        RECT 1663.090 2495.720 1668.690 2496.010 ;
        RECT 1669.530 2495.720 1675.130 2496.010 ;
        RECT 1675.970 2495.720 1681.570 2496.010 ;
        RECT 1682.410 2495.720 1688.470 2496.010 ;
        RECT 1689.310 2495.720 1694.910 2496.010 ;
        RECT 1695.750 2495.720 1701.350 2496.010 ;
        RECT 1702.190 2495.720 1707.790 2496.010 ;
        RECT 1708.630 2495.720 1714.230 2496.010 ;
        RECT 1715.070 2495.720 1720.670 2496.010 ;
        RECT 1721.510 2495.720 1727.110 2496.010 ;
        RECT 1727.950 2495.720 1733.550 2496.010 ;
        RECT 1734.390 2495.720 1739.990 2496.010 ;
        RECT 1740.830 2495.720 1746.430 2496.010 ;
        RECT 1747.270 2495.720 1752.870 2496.010 ;
        RECT 1753.710 2495.720 1759.310 2496.010 ;
        RECT 1760.150 2495.720 1765.750 2496.010 ;
        RECT 1766.590 2495.720 1772.190 2496.010 ;
        RECT 1773.030 2495.720 1778.630 2496.010 ;
        RECT 1779.470 2495.720 1785.070 2496.010 ;
        RECT 1785.910 2495.720 1791.510 2496.010 ;
        RECT 1792.350 2495.720 1797.950 2496.010 ;
        RECT 1798.790 2495.720 1804.390 2496.010 ;
        RECT 1805.230 2495.720 1810.830 2496.010 ;
        RECT 1811.670 2495.720 1817.270 2496.010 ;
        RECT 1818.110 2495.720 1823.710 2496.010 ;
        RECT 1824.550 2495.720 1830.150 2496.010 ;
        RECT 1830.990 2495.720 1836.590 2496.010 ;
        RECT 1837.430 2495.720 1843.030 2496.010 ;
        RECT 1843.870 2495.720 1849.470 2496.010 ;
        RECT 1850.310 2495.720 1855.910 2496.010 ;
        RECT 1856.750 2495.720 1862.350 2496.010 ;
        RECT 1863.190 2495.720 1868.790 2496.010 ;
        RECT 1869.630 2495.720 1875.230 2496.010 ;
        RECT 1876.070 2495.720 1881.670 2496.010 ;
        RECT 1882.510 2495.720 1888.110 2496.010 ;
        RECT 1888.950 2495.720 1894.550 2496.010 ;
        RECT 1895.390 2495.720 1900.990 2496.010 ;
        RECT 1901.830 2495.720 1907.430 2496.010 ;
        RECT 1908.270 2495.720 1913.870 2496.010 ;
        RECT 1914.710 2495.720 1920.310 2496.010 ;
        RECT 1921.150 2495.720 1926.750 2496.010 ;
        RECT 1927.590 2495.720 1933.190 2496.010 ;
        RECT 1934.030 2495.720 1939.630 2496.010 ;
        RECT 1940.470 2495.720 1940.580 2496.010 ;
        RECT 1150.550 1704.280 1940.580 2495.720 ;
        RECT 1151.110 1704.000 1151.650 1704.280 ;
        RECT 1152.490 1704.000 1153.490 1704.280 ;
        RECT 1154.330 1704.000 1154.870 1704.280 ;
        RECT 1155.710 1704.000 1156.710 1704.280 ;
        RECT 1157.550 1704.000 1158.090 1704.280 ;
        RECT 1158.930 1704.000 1159.930 1704.280 ;
        RECT 1160.770 1704.000 1161.310 1704.280 ;
        RECT 1162.150 1704.000 1163.150 1704.280 ;
        RECT 1163.990 1704.000 1164.530 1704.280 ;
        RECT 1165.370 1704.000 1166.370 1704.280 ;
        RECT 1167.210 1704.000 1167.750 1704.280 ;
        RECT 1168.590 1704.000 1169.590 1704.280 ;
        RECT 1170.430 1704.000 1170.970 1704.280 ;
        RECT 1171.810 1704.000 1172.810 1704.280 ;
        RECT 1173.650 1704.000 1174.190 1704.280 ;
        RECT 1175.030 1704.000 1176.030 1704.280 ;
        RECT 1176.870 1704.000 1177.410 1704.280 ;
        RECT 1178.250 1704.000 1179.250 1704.280 ;
        RECT 1180.090 1704.000 1180.630 1704.280 ;
        RECT 1181.470 1704.000 1182.470 1704.280 ;
        RECT 1183.310 1704.000 1183.850 1704.280 ;
        RECT 1184.690 1704.000 1185.690 1704.280 ;
        RECT 1186.530 1704.000 1187.070 1704.280 ;
        RECT 1187.910 1704.000 1188.910 1704.280 ;
        RECT 1189.750 1704.000 1190.290 1704.280 ;
        RECT 1191.130 1704.000 1192.130 1704.280 ;
        RECT 1192.970 1704.000 1193.510 1704.280 ;
        RECT 1194.350 1704.000 1195.350 1704.280 ;
        RECT 1196.190 1704.000 1196.730 1704.280 ;
        RECT 1197.570 1704.000 1198.570 1704.280 ;
        RECT 1199.410 1704.000 1199.950 1704.280 ;
        RECT 1200.790 1704.000 1201.790 1704.280 ;
        RECT 1202.630 1704.000 1203.170 1704.280 ;
        RECT 1204.010 1704.000 1205.010 1704.280 ;
        RECT 1205.850 1704.000 1206.390 1704.280 ;
        RECT 1207.230 1704.000 1208.230 1704.280 ;
        RECT 1209.070 1704.000 1209.610 1704.280 ;
        RECT 1210.450 1704.000 1211.450 1704.280 ;
        RECT 1212.290 1704.000 1212.830 1704.280 ;
        RECT 1213.670 1704.000 1214.670 1704.280 ;
        RECT 1215.510 1704.000 1216.050 1704.280 ;
        RECT 1216.890 1704.000 1217.890 1704.280 ;
        RECT 1218.730 1704.000 1219.270 1704.280 ;
        RECT 1220.110 1704.000 1221.110 1704.280 ;
        RECT 1221.950 1704.000 1222.490 1704.280 ;
        RECT 1223.330 1704.000 1224.330 1704.280 ;
        RECT 1225.170 1704.000 1225.710 1704.280 ;
        RECT 1226.550 1704.000 1227.550 1704.280 ;
        RECT 1228.390 1704.000 1228.930 1704.280 ;
        RECT 1229.770 1704.000 1230.770 1704.280 ;
        RECT 1231.610 1704.000 1232.150 1704.280 ;
        RECT 1232.990 1704.000 1233.990 1704.280 ;
        RECT 1234.830 1704.000 1235.370 1704.280 ;
        RECT 1236.210 1704.000 1237.210 1704.280 ;
        RECT 1238.050 1704.000 1238.590 1704.280 ;
        RECT 1239.430 1704.000 1240.430 1704.280 ;
        RECT 1241.270 1704.000 1241.810 1704.280 ;
        RECT 1242.650 1704.000 1243.650 1704.280 ;
        RECT 1244.490 1704.000 1245.030 1704.280 ;
        RECT 1245.870 1704.000 1246.870 1704.280 ;
        RECT 1247.710 1704.000 1248.250 1704.280 ;
        RECT 1249.090 1704.000 1250.090 1704.280 ;
        RECT 1250.930 1704.000 1251.470 1704.280 ;
        RECT 1252.310 1704.000 1253.310 1704.280 ;
        RECT 1254.150 1704.000 1254.690 1704.280 ;
        RECT 1255.530 1704.000 1256.530 1704.280 ;
        RECT 1257.370 1704.000 1257.910 1704.280 ;
        RECT 1258.750 1704.000 1259.750 1704.280 ;
        RECT 1260.590 1704.000 1261.130 1704.280 ;
        RECT 1261.970 1704.000 1262.970 1704.280 ;
        RECT 1263.810 1704.000 1264.350 1704.280 ;
        RECT 1265.190 1704.000 1266.190 1704.280 ;
        RECT 1267.030 1704.000 1267.570 1704.280 ;
        RECT 1268.410 1704.000 1269.410 1704.280 ;
        RECT 1270.250 1704.000 1270.790 1704.280 ;
        RECT 1271.630 1704.000 1272.630 1704.280 ;
        RECT 1273.470 1704.000 1274.010 1704.280 ;
        RECT 1274.850 1704.000 1275.850 1704.280 ;
        RECT 1276.690 1704.000 1277.230 1704.280 ;
        RECT 1278.070 1704.000 1279.070 1704.280 ;
        RECT 1279.910 1704.000 1280.450 1704.280 ;
        RECT 1281.290 1704.000 1282.290 1704.280 ;
        RECT 1283.130 1704.000 1284.130 1704.280 ;
        RECT 1284.970 1704.000 1285.510 1704.280 ;
        RECT 1286.350 1704.000 1287.350 1704.280 ;
        RECT 1288.190 1704.000 1288.730 1704.280 ;
        RECT 1289.570 1704.000 1290.570 1704.280 ;
        RECT 1291.410 1704.000 1291.950 1704.280 ;
        RECT 1292.790 1704.000 1293.790 1704.280 ;
        RECT 1294.630 1704.000 1295.170 1704.280 ;
        RECT 1296.010 1704.000 1297.010 1704.280 ;
        RECT 1297.850 1704.000 1298.390 1704.280 ;
        RECT 1299.230 1704.000 1300.230 1704.280 ;
        RECT 1301.070 1704.000 1301.610 1704.280 ;
        RECT 1302.450 1704.000 1303.450 1704.280 ;
        RECT 1304.290 1704.000 1304.830 1704.280 ;
        RECT 1305.670 1704.000 1306.670 1704.280 ;
        RECT 1307.510 1704.000 1308.050 1704.280 ;
        RECT 1308.890 1704.000 1309.890 1704.280 ;
        RECT 1310.730 1704.000 1311.270 1704.280 ;
        RECT 1312.110 1704.000 1313.110 1704.280 ;
        RECT 1313.950 1704.000 1314.490 1704.280 ;
        RECT 1315.330 1704.000 1316.330 1704.280 ;
        RECT 1317.170 1704.000 1317.710 1704.280 ;
        RECT 1318.550 1704.000 1319.550 1704.280 ;
        RECT 1320.390 1704.000 1320.930 1704.280 ;
        RECT 1321.770 1704.000 1322.770 1704.280 ;
        RECT 1323.610 1704.000 1324.150 1704.280 ;
        RECT 1324.990 1704.000 1325.990 1704.280 ;
        RECT 1326.830 1704.000 1327.370 1704.280 ;
        RECT 1328.210 1704.000 1329.210 1704.280 ;
        RECT 1330.050 1704.000 1330.590 1704.280 ;
        RECT 1331.430 1704.000 1332.430 1704.280 ;
        RECT 1333.270 1704.000 1333.810 1704.280 ;
        RECT 1334.650 1704.000 1335.650 1704.280 ;
        RECT 1336.490 1704.000 1337.030 1704.280 ;
        RECT 1337.870 1704.000 1338.870 1704.280 ;
        RECT 1339.710 1704.000 1340.250 1704.280 ;
        RECT 1341.090 1704.000 1342.090 1704.280 ;
        RECT 1342.930 1704.000 1343.470 1704.280 ;
        RECT 1344.310 1704.000 1345.310 1704.280 ;
        RECT 1346.150 1704.000 1346.690 1704.280 ;
        RECT 1347.530 1704.000 1348.530 1704.280 ;
        RECT 1349.370 1704.000 1349.910 1704.280 ;
        RECT 1350.750 1704.000 1351.750 1704.280 ;
        RECT 1352.590 1704.000 1353.130 1704.280 ;
        RECT 1353.970 1704.000 1354.970 1704.280 ;
        RECT 1355.810 1704.000 1356.350 1704.280 ;
        RECT 1357.190 1704.000 1358.190 1704.280 ;
        RECT 1359.030 1704.000 1359.570 1704.280 ;
        RECT 1360.410 1704.000 1361.410 1704.280 ;
        RECT 1362.250 1704.000 1362.790 1704.280 ;
        RECT 1363.630 1704.000 1364.630 1704.280 ;
        RECT 1365.470 1704.000 1366.010 1704.280 ;
        RECT 1366.850 1704.000 1367.850 1704.280 ;
        RECT 1368.690 1704.000 1369.230 1704.280 ;
        RECT 1370.070 1704.000 1371.070 1704.280 ;
        RECT 1371.910 1704.000 1372.450 1704.280 ;
        RECT 1373.290 1704.000 1374.290 1704.280 ;
        RECT 1375.130 1704.000 1375.670 1704.280 ;
        RECT 1376.510 1704.000 1377.510 1704.280 ;
        RECT 1378.350 1704.000 1378.890 1704.280 ;
        RECT 1379.730 1704.000 1380.730 1704.280 ;
        RECT 1381.570 1704.000 1382.110 1704.280 ;
        RECT 1382.950 1704.000 1383.950 1704.280 ;
        RECT 1384.790 1704.000 1385.330 1704.280 ;
        RECT 1386.170 1704.000 1387.170 1704.280 ;
        RECT 1388.010 1704.000 1388.550 1704.280 ;
        RECT 1389.390 1704.000 1390.390 1704.280 ;
        RECT 1391.230 1704.000 1391.770 1704.280 ;
        RECT 1392.610 1704.000 1393.610 1704.280 ;
        RECT 1394.450 1704.000 1394.990 1704.280 ;
        RECT 1395.830 1704.000 1396.830 1704.280 ;
        RECT 1397.670 1704.000 1398.210 1704.280 ;
        RECT 1399.050 1704.000 1400.050 1704.280 ;
        RECT 1400.890 1704.000 1401.430 1704.280 ;
        RECT 1402.270 1704.000 1403.270 1704.280 ;
        RECT 1404.110 1704.000 1404.650 1704.280 ;
        RECT 1405.490 1704.000 1406.490 1704.280 ;
        RECT 1407.330 1704.000 1407.870 1704.280 ;
        RECT 1408.710 1704.000 1409.710 1704.280 ;
        RECT 1410.550 1704.000 1411.090 1704.280 ;
        RECT 1411.930 1704.000 1412.930 1704.280 ;
        RECT 1413.770 1704.000 1414.310 1704.280 ;
        RECT 1415.150 1704.000 1416.150 1704.280 ;
        RECT 1416.990 1704.000 1417.990 1704.280 ;
        RECT 1418.830 1704.000 1419.370 1704.280 ;
        RECT 1420.210 1704.000 1421.210 1704.280 ;
        RECT 1422.050 1704.000 1422.590 1704.280 ;
        RECT 1423.430 1704.000 1424.430 1704.280 ;
        RECT 1425.270 1704.000 1425.810 1704.280 ;
        RECT 1426.650 1704.000 1427.650 1704.280 ;
        RECT 1428.490 1704.000 1429.030 1704.280 ;
        RECT 1429.870 1704.000 1430.870 1704.280 ;
        RECT 1431.710 1704.000 1432.250 1704.280 ;
        RECT 1433.090 1704.000 1434.090 1704.280 ;
        RECT 1434.930 1704.000 1435.470 1704.280 ;
        RECT 1436.310 1704.000 1437.310 1704.280 ;
        RECT 1438.150 1704.000 1438.690 1704.280 ;
        RECT 1439.530 1704.000 1440.530 1704.280 ;
        RECT 1441.370 1704.000 1441.910 1704.280 ;
        RECT 1442.750 1704.000 1443.750 1704.280 ;
        RECT 1444.590 1704.000 1445.130 1704.280 ;
        RECT 1445.970 1704.000 1446.970 1704.280 ;
        RECT 1447.810 1704.000 1448.350 1704.280 ;
        RECT 1449.190 1704.000 1450.190 1704.280 ;
        RECT 1451.030 1704.000 1451.570 1704.280 ;
        RECT 1452.410 1704.000 1453.410 1704.280 ;
        RECT 1454.250 1704.000 1454.790 1704.280 ;
        RECT 1455.630 1704.000 1456.630 1704.280 ;
        RECT 1457.470 1704.000 1458.010 1704.280 ;
        RECT 1458.850 1704.000 1459.850 1704.280 ;
        RECT 1460.690 1704.000 1461.230 1704.280 ;
        RECT 1462.070 1704.000 1463.070 1704.280 ;
        RECT 1463.910 1704.000 1464.450 1704.280 ;
        RECT 1465.290 1704.000 1466.290 1704.280 ;
        RECT 1467.130 1704.000 1467.670 1704.280 ;
        RECT 1468.510 1704.000 1469.510 1704.280 ;
        RECT 1470.350 1704.000 1470.890 1704.280 ;
        RECT 1471.730 1704.000 1472.730 1704.280 ;
        RECT 1473.570 1704.000 1474.110 1704.280 ;
        RECT 1474.950 1704.000 1475.950 1704.280 ;
        RECT 1476.790 1704.000 1477.330 1704.280 ;
        RECT 1478.170 1704.000 1479.170 1704.280 ;
        RECT 1480.010 1704.000 1480.550 1704.280 ;
        RECT 1481.390 1704.000 1482.390 1704.280 ;
        RECT 1483.230 1704.000 1483.770 1704.280 ;
        RECT 1484.610 1704.000 1485.610 1704.280 ;
        RECT 1486.450 1704.000 1486.990 1704.280 ;
        RECT 1487.830 1704.000 1488.830 1704.280 ;
        RECT 1489.670 1704.000 1490.210 1704.280 ;
        RECT 1491.050 1704.000 1492.050 1704.280 ;
        RECT 1492.890 1704.000 1493.430 1704.280 ;
        RECT 1494.270 1704.000 1495.270 1704.280 ;
        RECT 1496.110 1704.000 1496.650 1704.280 ;
        RECT 1497.490 1704.000 1498.490 1704.280 ;
        RECT 1499.330 1704.000 1499.870 1704.280 ;
        RECT 1500.710 1704.000 1501.710 1704.280 ;
        RECT 1502.550 1704.000 1503.090 1704.280 ;
        RECT 1503.930 1704.000 1504.930 1704.280 ;
        RECT 1505.770 1704.000 1506.310 1704.280 ;
        RECT 1507.150 1704.000 1508.150 1704.280 ;
        RECT 1508.990 1704.000 1509.530 1704.280 ;
        RECT 1510.370 1704.000 1511.370 1704.280 ;
        RECT 1512.210 1704.000 1512.750 1704.280 ;
        RECT 1513.590 1704.000 1514.590 1704.280 ;
        RECT 1515.430 1704.000 1515.970 1704.280 ;
        RECT 1516.810 1704.000 1517.810 1704.280 ;
        RECT 1518.650 1704.000 1519.190 1704.280 ;
        RECT 1520.030 1704.000 1521.030 1704.280 ;
        RECT 1521.870 1704.000 1522.410 1704.280 ;
        RECT 1523.250 1704.000 1524.250 1704.280 ;
        RECT 1525.090 1704.000 1525.630 1704.280 ;
        RECT 1526.470 1704.000 1527.470 1704.280 ;
        RECT 1528.310 1704.000 1528.850 1704.280 ;
        RECT 1529.690 1704.000 1530.690 1704.280 ;
        RECT 1531.530 1704.000 1532.070 1704.280 ;
        RECT 1532.910 1704.000 1533.910 1704.280 ;
        RECT 1534.750 1704.000 1535.290 1704.280 ;
        RECT 1536.130 1704.000 1537.130 1704.280 ;
        RECT 1537.970 1704.000 1538.510 1704.280 ;
        RECT 1539.350 1704.000 1540.350 1704.280 ;
        RECT 1541.190 1704.000 1541.730 1704.280 ;
        RECT 1542.570 1704.000 1543.570 1704.280 ;
        RECT 1544.410 1704.000 1544.950 1704.280 ;
        RECT 1545.790 1704.000 1546.790 1704.280 ;
        RECT 1547.630 1704.000 1548.170 1704.280 ;
        RECT 1549.010 1704.000 1550.010 1704.280 ;
        RECT 1550.850 1704.000 1551.850 1704.280 ;
        RECT 1552.690 1704.000 1553.230 1704.280 ;
        RECT 1554.070 1704.000 1555.070 1704.280 ;
        RECT 1555.910 1704.000 1556.450 1704.280 ;
        RECT 1557.290 1704.000 1558.290 1704.280 ;
        RECT 1559.130 1704.000 1559.670 1704.280 ;
        RECT 1560.510 1704.000 1561.510 1704.280 ;
        RECT 1562.350 1704.000 1562.890 1704.280 ;
        RECT 1563.730 1704.000 1564.730 1704.280 ;
        RECT 1565.570 1704.000 1566.110 1704.280 ;
        RECT 1566.950 1704.000 1567.950 1704.280 ;
        RECT 1568.790 1704.000 1569.330 1704.280 ;
        RECT 1570.170 1704.000 1571.170 1704.280 ;
        RECT 1572.010 1704.000 1572.550 1704.280 ;
        RECT 1573.390 1704.000 1574.390 1704.280 ;
        RECT 1575.230 1704.000 1575.770 1704.280 ;
        RECT 1576.610 1704.000 1577.610 1704.280 ;
        RECT 1578.450 1704.000 1578.990 1704.280 ;
        RECT 1579.830 1704.000 1580.830 1704.280 ;
        RECT 1581.670 1704.000 1582.210 1704.280 ;
        RECT 1583.050 1704.000 1584.050 1704.280 ;
        RECT 1584.890 1704.000 1585.430 1704.280 ;
        RECT 1586.270 1704.000 1587.270 1704.280 ;
        RECT 1588.110 1704.000 1588.650 1704.280 ;
        RECT 1589.490 1704.000 1590.490 1704.280 ;
        RECT 1591.330 1704.000 1591.870 1704.280 ;
        RECT 1592.710 1704.000 1593.710 1704.280 ;
        RECT 1594.550 1704.000 1595.090 1704.280 ;
        RECT 1595.930 1704.000 1596.930 1704.280 ;
        RECT 1597.770 1704.000 1598.310 1704.280 ;
        RECT 1599.150 1704.000 1600.150 1704.280 ;
        RECT 1600.990 1704.000 1601.530 1704.280 ;
        RECT 1602.370 1704.000 1603.370 1704.280 ;
        RECT 1604.210 1704.000 1604.750 1704.280 ;
        RECT 1605.590 1704.000 1606.590 1704.280 ;
        RECT 1607.430 1704.000 1607.970 1704.280 ;
        RECT 1608.810 1704.000 1609.810 1704.280 ;
        RECT 1610.650 1704.000 1611.190 1704.280 ;
        RECT 1612.030 1704.000 1613.030 1704.280 ;
        RECT 1613.870 1704.000 1614.410 1704.280 ;
        RECT 1615.250 1704.000 1616.250 1704.280 ;
        RECT 1617.090 1704.000 1617.630 1704.280 ;
        RECT 1618.470 1704.000 1619.470 1704.280 ;
        RECT 1620.310 1704.000 1620.850 1704.280 ;
        RECT 1621.690 1704.000 1622.690 1704.280 ;
        RECT 1623.530 1704.000 1624.070 1704.280 ;
        RECT 1624.910 1704.000 1625.910 1704.280 ;
        RECT 1626.750 1704.000 1627.290 1704.280 ;
        RECT 1628.130 1704.000 1629.130 1704.280 ;
        RECT 1629.970 1704.000 1630.510 1704.280 ;
        RECT 1631.350 1704.000 1632.350 1704.280 ;
        RECT 1633.190 1704.000 1633.730 1704.280 ;
        RECT 1634.570 1704.000 1635.570 1704.280 ;
        RECT 1636.410 1704.000 1636.950 1704.280 ;
        RECT 1637.790 1704.000 1638.790 1704.280 ;
        RECT 1639.630 1704.000 1640.170 1704.280 ;
        RECT 1641.010 1704.000 1642.010 1704.280 ;
        RECT 1642.850 1704.000 1643.390 1704.280 ;
        RECT 1644.230 1704.000 1645.230 1704.280 ;
        RECT 1646.070 1704.000 1646.610 1704.280 ;
        RECT 1647.450 1704.000 1648.450 1704.280 ;
        RECT 1649.290 1704.000 1649.830 1704.280 ;
        RECT 1650.670 1704.000 1651.670 1704.280 ;
        RECT 1652.510 1704.000 1653.050 1704.280 ;
        RECT 1653.890 1704.000 1654.890 1704.280 ;
        RECT 1655.730 1704.000 1656.270 1704.280 ;
        RECT 1657.110 1704.000 1658.110 1704.280 ;
        RECT 1658.950 1704.000 1659.490 1704.280 ;
        RECT 1660.330 1704.000 1661.330 1704.280 ;
        RECT 1662.170 1704.000 1662.710 1704.280 ;
        RECT 1663.550 1704.000 1664.550 1704.280 ;
        RECT 1665.390 1704.000 1665.930 1704.280 ;
        RECT 1666.770 1704.000 1667.770 1704.280 ;
        RECT 1668.610 1704.000 1669.150 1704.280 ;
        RECT 1669.990 1704.000 1670.990 1704.280 ;
        RECT 1671.830 1704.000 1672.370 1704.280 ;
        RECT 1673.210 1704.000 1674.210 1704.280 ;
        RECT 1675.050 1704.000 1675.590 1704.280 ;
        RECT 1676.430 1704.000 1677.430 1704.280 ;
        RECT 1678.270 1704.000 1678.810 1704.280 ;
        RECT 1679.650 1704.000 1680.650 1704.280 ;
        RECT 1681.490 1704.000 1682.030 1704.280 ;
        RECT 1682.870 1704.000 1683.870 1704.280 ;
        RECT 1684.710 1704.000 1685.710 1704.280 ;
        RECT 1686.550 1704.000 1687.090 1704.280 ;
        RECT 1687.930 1704.000 1688.930 1704.280 ;
        RECT 1689.770 1704.000 1690.310 1704.280 ;
        RECT 1691.150 1704.000 1692.150 1704.280 ;
        RECT 1692.990 1704.000 1693.530 1704.280 ;
        RECT 1694.370 1704.000 1695.370 1704.280 ;
        RECT 1696.210 1704.000 1696.750 1704.280 ;
        RECT 1697.590 1704.000 1698.590 1704.280 ;
        RECT 1699.430 1704.000 1699.970 1704.280 ;
        RECT 1700.810 1704.000 1701.810 1704.280 ;
        RECT 1702.650 1704.000 1703.190 1704.280 ;
        RECT 1704.030 1704.000 1705.030 1704.280 ;
        RECT 1705.870 1704.000 1706.410 1704.280 ;
        RECT 1707.250 1704.000 1708.250 1704.280 ;
        RECT 1709.090 1704.000 1709.630 1704.280 ;
        RECT 1710.470 1704.000 1711.470 1704.280 ;
        RECT 1712.310 1704.000 1712.850 1704.280 ;
        RECT 1713.690 1704.000 1714.690 1704.280 ;
        RECT 1715.530 1704.000 1716.070 1704.280 ;
        RECT 1716.910 1704.000 1717.910 1704.280 ;
        RECT 1718.750 1704.000 1719.290 1704.280 ;
        RECT 1720.130 1704.000 1721.130 1704.280 ;
        RECT 1721.970 1704.000 1722.510 1704.280 ;
        RECT 1723.350 1704.000 1724.350 1704.280 ;
        RECT 1725.190 1704.000 1725.730 1704.280 ;
        RECT 1726.570 1704.000 1727.570 1704.280 ;
        RECT 1728.410 1704.000 1728.950 1704.280 ;
        RECT 1729.790 1704.000 1730.790 1704.280 ;
        RECT 1731.630 1704.000 1732.170 1704.280 ;
        RECT 1733.010 1704.000 1734.010 1704.280 ;
        RECT 1734.850 1704.000 1735.390 1704.280 ;
        RECT 1736.230 1704.000 1737.230 1704.280 ;
        RECT 1738.070 1704.000 1738.610 1704.280 ;
        RECT 1739.450 1704.000 1740.450 1704.280 ;
        RECT 1741.290 1704.000 1741.830 1704.280 ;
        RECT 1742.670 1704.000 1743.670 1704.280 ;
        RECT 1744.510 1704.000 1745.050 1704.280 ;
        RECT 1745.890 1704.000 1746.890 1704.280 ;
        RECT 1747.730 1704.000 1748.270 1704.280 ;
        RECT 1749.110 1704.000 1750.110 1704.280 ;
        RECT 1750.950 1704.000 1751.490 1704.280 ;
        RECT 1752.330 1704.000 1753.330 1704.280 ;
        RECT 1754.170 1704.000 1754.710 1704.280 ;
        RECT 1755.550 1704.000 1756.550 1704.280 ;
        RECT 1757.390 1704.000 1757.930 1704.280 ;
        RECT 1758.770 1704.000 1759.770 1704.280 ;
        RECT 1760.610 1704.000 1761.150 1704.280 ;
        RECT 1761.990 1704.000 1762.990 1704.280 ;
        RECT 1763.830 1704.000 1764.370 1704.280 ;
        RECT 1765.210 1704.000 1766.210 1704.280 ;
        RECT 1767.050 1704.000 1767.590 1704.280 ;
        RECT 1768.430 1704.000 1769.430 1704.280 ;
        RECT 1770.270 1704.000 1770.810 1704.280 ;
        RECT 1771.650 1704.000 1772.650 1704.280 ;
        RECT 1773.490 1704.000 1774.030 1704.280 ;
        RECT 1774.870 1704.000 1775.870 1704.280 ;
        RECT 1776.710 1704.000 1777.250 1704.280 ;
        RECT 1778.090 1704.000 1779.090 1704.280 ;
        RECT 1779.930 1704.000 1780.470 1704.280 ;
        RECT 1781.310 1704.000 1782.310 1704.280 ;
        RECT 1783.150 1704.000 1783.690 1704.280 ;
        RECT 1784.530 1704.000 1785.530 1704.280 ;
        RECT 1786.370 1704.000 1786.910 1704.280 ;
        RECT 1787.750 1704.000 1788.750 1704.280 ;
        RECT 1789.590 1704.000 1790.130 1704.280 ;
        RECT 1790.970 1704.000 1791.970 1704.280 ;
        RECT 1792.810 1704.000 1793.350 1704.280 ;
        RECT 1794.190 1704.000 1795.190 1704.280 ;
        RECT 1796.030 1704.000 1796.570 1704.280 ;
        RECT 1797.410 1704.000 1798.410 1704.280 ;
        RECT 1799.250 1704.000 1799.790 1704.280 ;
        RECT 1800.630 1704.000 1801.630 1704.280 ;
        RECT 1802.470 1704.000 1803.010 1704.280 ;
        RECT 1803.850 1704.000 1804.850 1704.280 ;
        RECT 1805.690 1704.000 1806.230 1704.280 ;
        RECT 1807.070 1704.000 1808.070 1704.280 ;
        RECT 1808.910 1704.000 1809.450 1704.280 ;
        RECT 1810.290 1704.000 1811.290 1704.280 ;
        RECT 1812.130 1704.000 1812.670 1704.280 ;
        RECT 1813.510 1704.000 1814.510 1704.280 ;
        RECT 1815.350 1704.000 1815.890 1704.280 ;
        RECT 1816.730 1704.000 1817.730 1704.280 ;
        RECT 1818.570 1704.000 1819.570 1704.280 ;
        RECT 1820.410 1704.000 1820.950 1704.280 ;
        RECT 1821.790 1704.000 1822.790 1704.280 ;
        RECT 1823.630 1704.000 1824.170 1704.280 ;
        RECT 1825.010 1704.000 1826.010 1704.280 ;
        RECT 1826.850 1704.000 1827.390 1704.280 ;
        RECT 1828.230 1704.000 1829.230 1704.280 ;
        RECT 1830.070 1704.000 1830.610 1704.280 ;
        RECT 1831.450 1704.000 1832.450 1704.280 ;
        RECT 1833.290 1704.000 1833.830 1704.280 ;
        RECT 1834.670 1704.000 1835.670 1704.280 ;
        RECT 1836.510 1704.000 1837.050 1704.280 ;
        RECT 1837.890 1704.000 1838.890 1704.280 ;
        RECT 1839.730 1704.000 1840.270 1704.280 ;
        RECT 1841.110 1704.000 1842.110 1704.280 ;
        RECT 1842.950 1704.000 1843.490 1704.280 ;
        RECT 1844.330 1704.000 1845.330 1704.280 ;
        RECT 1846.170 1704.000 1846.710 1704.280 ;
        RECT 1847.550 1704.000 1848.550 1704.280 ;
        RECT 1849.390 1704.000 1849.930 1704.280 ;
        RECT 1850.770 1704.000 1851.770 1704.280 ;
        RECT 1852.610 1704.000 1853.150 1704.280 ;
        RECT 1853.990 1704.000 1854.990 1704.280 ;
        RECT 1855.830 1704.000 1856.370 1704.280 ;
        RECT 1857.210 1704.000 1858.210 1704.280 ;
        RECT 1859.050 1704.000 1859.590 1704.280 ;
        RECT 1860.430 1704.000 1861.430 1704.280 ;
        RECT 1862.270 1704.000 1862.810 1704.280 ;
        RECT 1863.650 1704.000 1864.650 1704.280 ;
        RECT 1865.490 1704.000 1866.030 1704.280 ;
        RECT 1866.870 1704.000 1867.870 1704.280 ;
        RECT 1868.710 1704.000 1869.250 1704.280 ;
        RECT 1870.090 1704.000 1871.090 1704.280 ;
        RECT 1871.930 1704.000 1872.470 1704.280 ;
        RECT 1873.310 1704.000 1874.310 1704.280 ;
        RECT 1875.150 1704.000 1875.690 1704.280 ;
        RECT 1876.530 1704.000 1877.530 1704.280 ;
        RECT 1878.370 1704.000 1878.910 1704.280 ;
        RECT 1879.750 1704.000 1880.750 1704.280 ;
        RECT 1881.590 1704.000 1882.130 1704.280 ;
        RECT 1882.970 1704.000 1883.970 1704.280 ;
        RECT 1884.810 1704.000 1885.350 1704.280 ;
        RECT 1886.190 1704.000 1887.190 1704.280 ;
        RECT 1888.030 1704.000 1888.570 1704.280 ;
        RECT 1889.410 1704.000 1890.410 1704.280 ;
        RECT 1891.250 1704.000 1891.790 1704.280 ;
        RECT 1892.630 1704.000 1893.630 1704.280 ;
        RECT 1894.470 1704.000 1895.010 1704.280 ;
        RECT 1895.850 1704.000 1896.850 1704.280 ;
        RECT 1897.690 1704.000 1898.230 1704.280 ;
        RECT 1899.070 1704.000 1900.070 1704.280 ;
        RECT 1900.910 1704.000 1901.450 1704.280 ;
        RECT 1902.290 1704.000 1903.290 1704.280 ;
        RECT 1904.130 1704.000 1904.670 1704.280 ;
        RECT 1905.510 1704.000 1906.510 1704.280 ;
        RECT 1907.350 1704.000 1907.890 1704.280 ;
        RECT 1908.730 1704.000 1909.730 1704.280 ;
        RECT 1910.570 1704.000 1911.110 1704.280 ;
        RECT 1911.950 1704.000 1912.950 1704.280 ;
        RECT 1913.790 1704.000 1914.330 1704.280 ;
        RECT 1915.170 1704.000 1916.170 1704.280 ;
        RECT 1917.010 1704.000 1917.550 1704.280 ;
        RECT 1918.390 1704.000 1919.390 1704.280 ;
        RECT 1920.230 1704.000 1920.770 1704.280 ;
        RECT 1921.610 1704.000 1922.610 1704.280 ;
        RECT 1923.450 1704.000 1923.990 1704.280 ;
        RECT 1924.830 1704.000 1925.830 1704.280 ;
        RECT 1926.670 1704.000 1927.210 1704.280 ;
        RECT 1928.050 1704.000 1929.050 1704.280 ;
        RECT 1929.890 1704.000 1930.430 1704.280 ;
        RECT 1931.270 1704.000 1932.270 1704.280 ;
        RECT 1933.110 1704.000 1933.650 1704.280 ;
        RECT 1934.490 1704.000 1935.490 1704.280 ;
        RECT 1936.330 1704.000 1936.870 1704.280 ;
        RECT 1937.710 1704.000 1938.710 1704.280 ;
        RECT 1939.550 1704.000 1940.090 1704.280 ;
      LAYER met3 ;
        RECT 1150.525 2455.840 1940.640 2488.965 ;
        RECT 1154.400 2454.440 1940.640 2455.840 ;
        RECT 1150.525 2366.760 1940.640 2454.440 ;
        RECT 1154.400 2365.360 1940.640 2366.760 ;
        RECT 1150.525 2278.360 1940.640 2365.360 ;
        RECT 1154.400 2276.960 1940.640 2278.360 ;
        RECT 1150.525 2189.280 1940.640 2276.960 ;
        RECT 1154.400 2187.880 1940.640 2189.280 ;
        RECT 1150.525 2100.200 1940.640 2187.880 ;
        RECT 1154.400 2098.800 1940.640 2100.200 ;
        RECT 1150.525 2011.800 1940.640 2098.800 ;
        RECT 1154.400 2010.400 1940.640 2011.800 ;
        RECT 1150.525 1922.720 1940.640 2010.400 ;
        RECT 1154.400 1921.320 1940.640 1922.720 ;
        RECT 1150.525 1833.640 1940.640 1921.320 ;
        RECT 1154.400 1832.240 1940.640 1833.640 ;
        RECT 1150.525 1745.240 1940.640 1832.240 ;
        RECT 1154.400 1743.840 1940.640 1745.240 ;
        RECT 1150.525 1704.255 1940.640 1743.840 ;
      LAYER met4 ;
        RECT 1171.040 1710.640 1172.640 2489.040 ;
        RECT 1247.840 1710.640 1249.440 2489.040 ;
      LAYER met4 ;
        RECT 1303.020 1710.640 1318.020 2489.040 ;
        RECT 1321.020 1710.640 1354.020 2489.040 ;
        RECT 1357.020 1710.640 1372.020 2489.040 ;
        RECT 1375.020 1710.640 1390.020 2489.040 ;
        RECT 1393.020 1710.640 1408.020 2489.040 ;
        RECT 1411.020 1710.640 1444.020 2489.040 ;
        RECT 1447.020 1710.640 1462.020 2489.040 ;
        RECT 1465.020 1710.640 1480.020 2489.040 ;
        RECT 1483.020 1710.640 1498.020 2489.040 ;
        RECT 1501.020 1710.640 1534.020 2489.040 ;
        RECT 1537.020 1710.640 1552.020 2489.040 ;
        RECT 1555.020 1710.640 1570.020 2489.040 ;
        RECT 1573.020 1710.640 1588.020 2489.040 ;
        RECT 1591.020 1710.640 1624.020 2489.040 ;
        RECT 1627.020 1710.640 1642.020 2489.040 ;
        RECT 1645.020 1710.640 1660.020 2489.040 ;
        RECT 1663.020 1710.640 1678.020 2489.040 ;
        RECT 1681.020 1710.640 1714.020 2489.040 ;
        RECT 1717.020 1710.640 1732.020 2489.040 ;
        RECT 1735.020 1710.640 1750.020 2489.040 ;
        RECT 1753.020 1710.640 1768.020 2489.040 ;
        RECT 1771.020 1710.640 1804.020 2489.040 ;
        RECT 1807.020 1710.640 1822.020 2489.040 ;
        RECT 1825.020 1710.640 1840.020 2489.040 ;
        RECT 1843.020 1710.640 1858.020 2489.040 ;
        RECT 1861.020 1710.640 1894.020 2489.040 ;
        RECT 1897.020 1710.640 1912.020 2489.040 ;
        RECT 1915.020 1710.640 1930.020 2489.040 ;
        RECT 1933.020 1710.640 1940.640 2489.040 ;
>>>>>>> Latest run - not LVS matched yet
  END
END user_project_wrapper
END LIBRARY

