magic
tech sky130A
magscale 1 2
timestamp 1608129410
<< obsli1 >>
rect 1104 2159 278852 237745
<< obsm1 >>
rect 1104 1232 278852 237776
<< metal2 >>
rect 1122 239200 1178 240000
rect 3422 239200 3478 240000
rect 5722 239200 5778 240000
rect 8114 239200 8170 240000
rect 10414 239200 10470 240000
rect 12714 239200 12770 240000
rect 15106 239200 15162 240000
rect 17406 239200 17462 240000
rect 19706 239200 19762 240000
rect 22098 239200 22154 240000
rect 24398 239200 24454 240000
rect 26698 239200 26754 240000
rect 29090 239200 29146 240000
rect 31390 239200 31446 240000
rect 33782 239200 33838 240000
rect 36082 239200 36138 240000
rect 38382 239200 38438 240000
rect 40774 239200 40830 240000
rect 43074 239200 43130 240000
rect 45374 239200 45430 240000
rect 47766 239200 47822 240000
rect 50066 239200 50122 240000
rect 52366 239200 52422 240000
rect 54758 239200 54814 240000
rect 57058 239200 57114 240000
rect 59358 239200 59414 240000
rect 61750 239200 61806 240000
rect 64050 239200 64106 240000
rect 66442 239200 66498 240000
rect 68742 239200 68798 240000
rect 71042 239200 71098 240000
rect 73434 239200 73490 240000
rect 75734 239200 75790 240000
rect 78034 239200 78090 240000
rect 80426 239200 80482 240000
rect 82726 239200 82782 240000
rect 85026 239200 85082 240000
rect 87418 239200 87474 240000
rect 89718 239200 89774 240000
rect 92018 239200 92074 240000
rect 94410 239200 94466 240000
rect 96710 239200 96766 240000
rect 99102 239200 99158 240000
rect 101402 239200 101458 240000
rect 103702 239200 103758 240000
rect 106094 239200 106150 240000
rect 108394 239200 108450 240000
rect 110694 239200 110750 240000
rect 113086 239200 113142 240000
rect 115386 239200 115442 240000
rect 117686 239200 117742 240000
rect 120078 239200 120134 240000
rect 122378 239200 122434 240000
rect 124678 239200 124734 240000
rect 127070 239200 127126 240000
rect 129370 239200 129426 240000
rect 131762 239200 131818 240000
rect 134062 239200 134118 240000
rect 136362 239200 136418 240000
rect 138754 239200 138810 240000
rect 141054 239200 141110 240000
rect 143354 239200 143410 240000
rect 145746 239200 145802 240000
rect 148046 239200 148102 240000
rect 150346 239200 150402 240000
rect 152738 239200 152794 240000
rect 155038 239200 155094 240000
rect 157430 239200 157486 240000
rect 159730 239200 159786 240000
rect 162030 239200 162086 240000
rect 164422 239200 164478 240000
rect 166722 239200 166778 240000
rect 169022 239200 169078 240000
rect 171414 239200 171470 240000
rect 173714 239200 173770 240000
rect 176014 239200 176070 240000
rect 178406 239200 178462 240000
rect 180706 239200 180762 240000
rect 183006 239200 183062 240000
rect 185398 239200 185454 240000
rect 187698 239200 187754 240000
rect 190090 239200 190146 240000
rect 192390 239200 192446 240000
rect 194690 239200 194746 240000
rect 197082 239200 197138 240000
rect 199382 239200 199438 240000
rect 201682 239200 201738 240000
rect 204074 239200 204130 240000
rect 206374 239200 206430 240000
rect 208674 239200 208730 240000
rect 211066 239200 211122 240000
rect 213366 239200 213422 240000
rect 215666 239200 215722 240000
rect 218058 239200 218114 240000
rect 220358 239200 220414 240000
rect 222750 239200 222806 240000
rect 225050 239200 225106 240000
rect 227350 239200 227406 240000
rect 229742 239200 229798 240000
rect 232042 239200 232098 240000
rect 234342 239200 234398 240000
rect 236734 239200 236790 240000
rect 239034 239200 239090 240000
rect 241334 239200 241390 240000
rect 243726 239200 243782 240000
rect 246026 239200 246082 240000
rect 248326 239200 248382 240000
rect 250718 239200 250774 240000
rect 253018 239200 253074 240000
rect 255410 239200 255466 240000
rect 257710 239200 257766 240000
rect 260010 239200 260066 240000
rect 262402 239200 262458 240000
rect 264702 239200 264758 240000
rect 267002 239200 267058 240000
rect 269394 239200 269450 240000
rect 271694 239200 271750 240000
rect 273994 239200 274050 240000
rect 276386 239200 276442 240000
rect 278686 239200 278742 240000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6366 0 6422 800
rect 6918 0 6974 800
rect 7470 0 7526 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 11978 0 12034 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17590 0 17646 800
rect 18142 0 18198 800
rect 18694 0 18750 800
rect 19246 0 19302 800
rect 19798 0 19854 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21454 0 21510 800
rect 22006 0 22062 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23754 0 23810 800
rect 24306 0 24362 800
rect 24858 0 24914 800
rect 25410 0 25466 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 27066 0 27122 800
rect 27618 0 27674 800
rect 28170 0 28226 800
rect 28722 0 28778 800
rect 29274 0 29330 800
rect 29826 0 29882 800
rect 30378 0 30434 800
rect 31022 0 31078 800
rect 31574 0 31630 800
rect 32126 0 32182 800
rect 32678 0 32734 800
rect 33230 0 33286 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 35438 0 35494 800
rect 35990 0 36046 800
rect 36542 0 36598 800
rect 37094 0 37150 800
rect 37646 0 37702 800
rect 38290 0 38346 800
rect 38842 0 38898 800
rect 39394 0 39450 800
rect 39946 0 40002 800
rect 40498 0 40554 800
rect 41050 0 41106 800
rect 41602 0 41658 800
rect 42154 0 42210 800
rect 42706 0 42762 800
rect 43258 0 43314 800
rect 43810 0 43866 800
rect 44362 0 44418 800
rect 44914 0 44970 800
rect 45466 0 45522 800
rect 46110 0 46166 800
rect 46662 0 46718 800
rect 47214 0 47270 800
rect 47766 0 47822 800
rect 48318 0 48374 800
rect 48870 0 48926 800
rect 49422 0 49478 800
rect 49974 0 50030 800
rect 50526 0 50582 800
rect 51078 0 51134 800
rect 51630 0 51686 800
rect 52182 0 52238 800
rect 52734 0 52790 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54482 0 54538 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58898 0 58954 800
rect 59450 0 59506 800
rect 60002 0 60058 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62854 0 62910 800
rect 63406 0 63462 800
rect 63958 0 64014 800
rect 64510 0 64566 800
rect 65062 0 65118 800
rect 65614 0 65670 800
rect 66166 0 66222 800
rect 66718 0 66774 800
rect 67270 0 67326 800
rect 67822 0 67878 800
rect 68466 0 68522 800
rect 69018 0 69074 800
rect 69570 0 69626 800
rect 70122 0 70178 800
rect 70674 0 70730 800
rect 71226 0 71282 800
rect 71778 0 71834 800
rect 72330 0 72386 800
rect 72882 0 72938 800
rect 73434 0 73490 800
rect 73986 0 74042 800
rect 74538 0 74594 800
rect 75090 0 75146 800
rect 75642 0 75698 800
rect 76286 0 76342 800
rect 76838 0 76894 800
rect 77390 0 77446 800
rect 77942 0 77998 800
rect 78494 0 78550 800
rect 79046 0 79102 800
rect 79598 0 79654 800
rect 80150 0 80206 800
rect 80702 0 80758 800
rect 81254 0 81310 800
rect 81806 0 81862 800
rect 82358 0 82414 800
rect 82910 0 82966 800
rect 83554 0 83610 800
rect 84106 0 84162 800
rect 84658 0 84714 800
rect 85210 0 85266 800
rect 85762 0 85818 800
rect 86314 0 86370 800
rect 86866 0 86922 800
rect 87418 0 87474 800
rect 87970 0 88026 800
rect 88522 0 88578 800
rect 89074 0 89130 800
rect 89626 0 89682 800
rect 90178 0 90234 800
rect 90730 0 90786 800
rect 91374 0 91430 800
rect 91926 0 91982 800
rect 92478 0 92534 800
rect 93030 0 93086 800
rect 93582 0 93638 800
rect 94134 0 94190 800
rect 94686 0 94742 800
rect 95238 0 95294 800
rect 95790 0 95846 800
rect 96342 0 96398 800
rect 96894 0 96950 800
rect 97446 0 97502 800
rect 97998 0 98054 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99746 0 99802 800
rect 100298 0 100354 800
rect 100850 0 100906 800
rect 101402 0 101458 800
rect 101954 0 102010 800
rect 102506 0 102562 800
rect 103058 0 103114 800
rect 103610 0 103666 800
rect 104162 0 104218 800
rect 104714 0 104770 800
rect 105266 0 105322 800
rect 105818 0 105874 800
rect 106462 0 106518 800
rect 107014 0 107070 800
rect 107566 0 107622 800
rect 108118 0 108174 800
rect 108670 0 108726 800
rect 109222 0 109278 800
rect 109774 0 109830 800
rect 110326 0 110382 800
rect 110878 0 110934 800
rect 111430 0 111486 800
rect 111982 0 112038 800
rect 112534 0 112590 800
rect 113086 0 113142 800
rect 113638 0 113694 800
rect 114282 0 114338 800
rect 114834 0 114890 800
rect 115386 0 115442 800
rect 115938 0 115994 800
rect 116490 0 116546 800
rect 117042 0 117098 800
rect 117594 0 117650 800
rect 118146 0 118202 800
rect 118698 0 118754 800
rect 119250 0 119306 800
rect 119802 0 119858 800
rect 120354 0 120410 800
rect 120906 0 120962 800
rect 121550 0 121606 800
rect 122102 0 122158 800
rect 122654 0 122710 800
rect 123206 0 123262 800
rect 123758 0 123814 800
rect 124310 0 124366 800
rect 124862 0 124918 800
rect 125414 0 125470 800
rect 125966 0 126022 800
rect 126518 0 126574 800
rect 127070 0 127126 800
rect 127622 0 127678 800
rect 128174 0 128230 800
rect 128726 0 128782 800
rect 129370 0 129426 800
rect 129922 0 129978 800
rect 130474 0 130530 800
rect 131026 0 131082 800
rect 131578 0 131634 800
rect 132130 0 132186 800
rect 132682 0 132738 800
rect 133234 0 133290 800
rect 133786 0 133842 800
rect 134338 0 134394 800
rect 134890 0 134946 800
rect 135442 0 135498 800
rect 135994 0 136050 800
rect 136638 0 136694 800
rect 137190 0 137246 800
rect 137742 0 137798 800
rect 138294 0 138350 800
rect 138846 0 138902 800
rect 139398 0 139454 800
rect 139950 0 140006 800
rect 140502 0 140558 800
rect 141054 0 141110 800
rect 141606 0 141662 800
rect 142158 0 142214 800
rect 142710 0 142766 800
rect 143262 0 143318 800
rect 143814 0 143870 800
rect 144458 0 144514 800
rect 145010 0 145066 800
rect 145562 0 145618 800
rect 146114 0 146170 800
rect 146666 0 146722 800
rect 147218 0 147274 800
rect 147770 0 147826 800
rect 148322 0 148378 800
rect 148874 0 148930 800
rect 149426 0 149482 800
rect 149978 0 150034 800
rect 150530 0 150586 800
rect 151082 0 151138 800
rect 151726 0 151782 800
rect 152278 0 152334 800
rect 152830 0 152886 800
rect 153382 0 153438 800
rect 153934 0 153990 800
rect 154486 0 154542 800
rect 155038 0 155094 800
rect 155590 0 155646 800
rect 156142 0 156198 800
rect 156694 0 156750 800
rect 157246 0 157302 800
rect 157798 0 157854 800
rect 158350 0 158406 800
rect 158902 0 158958 800
rect 159546 0 159602 800
rect 160098 0 160154 800
rect 160650 0 160706 800
rect 161202 0 161258 800
rect 161754 0 161810 800
rect 162306 0 162362 800
rect 162858 0 162914 800
rect 163410 0 163466 800
rect 163962 0 164018 800
rect 164514 0 164570 800
rect 165066 0 165122 800
rect 165618 0 165674 800
rect 166170 0 166226 800
rect 166814 0 166870 800
rect 167366 0 167422 800
rect 167918 0 167974 800
rect 168470 0 168526 800
rect 169022 0 169078 800
rect 169574 0 169630 800
rect 170126 0 170182 800
rect 170678 0 170734 800
rect 171230 0 171286 800
rect 171782 0 171838 800
rect 172334 0 172390 800
rect 172886 0 172942 800
rect 173438 0 173494 800
rect 173990 0 174046 800
rect 174634 0 174690 800
rect 175186 0 175242 800
rect 175738 0 175794 800
rect 176290 0 176346 800
rect 176842 0 176898 800
rect 177394 0 177450 800
rect 177946 0 178002 800
rect 178498 0 178554 800
rect 179050 0 179106 800
rect 179602 0 179658 800
rect 180154 0 180210 800
rect 180706 0 180762 800
rect 181258 0 181314 800
rect 181902 0 181958 800
rect 182454 0 182510 800
rect 183006 0 183062 800
rect 183558 0 183614 800
rect 184110 0 184166 800
rect 184662 0 184718 800
rect 185214 0 185270 800
rect 185766 0 185822 800
rect 186318 0 186374 800
rect 186870 0 186926 800
rect 187422 0 187478 800
rect 187974 0 188030 800
rect 188526 0 188582 800
rect 189078 0 189134 800
rect 189722 0 189778 800
rect 190274 0 190330 800
rect 190826 0 190882 800
rect 191378 0 191434 800
rect 191930 0 191986 800
rect 192482 0 192538 800
rect 193034 0 193090 800
rect 193586 0 193642 800
rect 194138 0 194194 800
rect 194690 0 194746 800
rect 195242 0 195298 800
rect 195794 0 195850 800
rect 196346 0 196402 800
rect 196898 0 196954 800
rect 197542 0 197598 800
rect 198094 0 198150 800
rect 198646 0 198702 800
rect 199198 0 199254 800
rect 199750 0 199806 800
rect 200302 0 200358 800
rect 200854 0 200910 800
rect 201406 0 201462 800
rect 201958 0 202014 800
rect 202510 0 202566 800
rect 203062 0 203118 800
rect 203614 0 203670 800
rect 204166 0 204222 800
rect 204810 0 204866 800
rect 205362 0 205418 800
rect 205914 0 205970 800
rect 206466 0 206522 800
rect 207018 0 207074 800
rect 207570 0 207626 800
rect 208122 0 208178 800
rect 208674 0 208730 800
rect 209226 0 209282 800
rect 209778 0 209834 800
rect 210330 0 210386 800
rect 210882 0 210938 800
rect 211434 0 211490 800
rect 211986 0 212042 800
rect 212630 0 212686 800
rect 213182 0 213238 800
rect 213734 0 213790 800
rect 214286 0 214342 800
rect 214838 0 214894 800
rect 215390 0 215446 800
rect 215942 0 215998 800
rect 216494 0 216550 800
rect 217046 0 217102 800
rect 217598 0 217654 800
rect 218150 0 218206 800
rect 218702 0 218758 800
rect 219254 0 219310 800
rect 219898 0 219954 800
rect 220450 0 220506 800
rect 221002 0 221058 800
rect 221554 0 221610 800
rect 222106 0 222162 800
rect 222658 0 222714 800
rect 223210 0 223266 800
rect 223762 0 223818 800
rect 224314 0 224370 800
rect 224866 0 224922 800
rect 225418 0 225474 800
rect 225970 0 226026 800
rect 226522 0 226578 800
rect 227074 0 227130 800
rect 227718 0 227774 800
rect 228270 0 228326 800
rect 228822 0 228878 800
rect 229374 0 229430 800
rect 229926 0 229982 800
rect 230478 0 230534 800
rect 231030 0 231086 800
rect 231582 0 231638 800
rect 232134 0 232190 800
rect 232686 0 232742 800
rect 233238 0 233294 800
rect 233790 0 233846 800
rect 234342 0 234398 800
rect 234986 0 235042 800
rect 235538 0 235594 800
rect 236090 0 236146 800
rect 236642 0 236698 800
rect 237194 0 237250 800
rect 237746 0 237802 800
rect 238298 0 238354 800
rect 238850 0 238906 800
rect 239402 0 239458 800
rect 239954 0 240010 800
rect 240506 0 240562 800
rect 241058 0 241114 800
rect 241610 0 241666 800
rect 242162 0 242218 800
rect 242806 0 242862 800
rect 243358 0 243414 800
rect 243910 0 243966 800
rect 244462 0 244518 800
rect 245014 0 245070 800
rect 245566 0 245622 800
rect 246118 0 246174 800
rect 246670 0 246726 800
rect 247222 0 247278 800
rect 247774 0 247830 800
rect 248326 0 248382 800
rect 248878 0 248934 800
rect 249430 0 249486 800
rect 250074 0 250130 800
rect 250626 0 250682 800
rect 251178 0 251234 800
rect 251730 0 251786 800
rect 252282 0 252338 800
rect 252834 0 252890 800
rect 253386 0 253442 800
rect 253938 0 253994 800
rect 254490 0 254546 800
rect 255042 0 255098 800
rect 255594 0 255650 800
rect 256146 0 256202 800
rect 256698 0 256754 800
rect 257250 0 257306 800
rect 257894 0 257950 800
rect 258446 0 258502 800
rect 258998 0 259054 800
rect 259550 0 259606 800
rect 260102 0 260158 800
rect 260654 0 260710 800
rect 261206 0 261262 800
rect 261758 0 261814 800
rect 262310 0 262366 800
rect 262862 0 262918 800
rect 263414 0 263470 800
rect 263966 0 264022 800
rect 264518 0 264574 800
rect 265162 0 265218 800
rect 265714 0 265770 800
rect 266266 0 266322 800
rect 266818 0 266874 800
rect 267370 0 267426 800
rect 267922 0 267978 800
rect 268474 0 268530 800
rect 269026 0 269082 800
rect 269578 0 269634 800
rect 270130 0 270186 800
rect 270682 0 270738 800
rect 271234 0 271290 800
rect 271786 0 271842 800
rect 272338 0 272394 800
rect 272982 0 273038 800
rect 273534 0 273590 800
rect 274086 0 274142 800
rect 274638 0 274694 800
rect 275190 0 275246 800
rect 275742 0 275798 800
rect 276294 0 276350 800
rect 276846 0 276902 800
rect 277398 0 277454 800
rect 277950 0 278006 800
rect 278502 0 278558 800
rect 279054 0 279110 800
rect 279606 0 279662 800
<< obsm2 >>
rect 294 239144 1066 239200
rect 1234 239144 3366 239200
rect 3534 239144 5666 239200
rect 5834 239144 8058 239200
rect 8226 239144 10358 239200
rect 10526 239144 12658 239200
rect 12826 239144 15050 239200
rect 15218 239144 17350 239200
rect 17518 239144 19650 239200
rect 19818 239144 22042 239200
rect 22210 239144 24342 239200
rect 24510 239144 26642 239200
rect 26810 239144 29034 239200
rect 29202 239144 31334 239200
rect 31502 239144 33726 239200
rect 33894 239144 36026 239200
rect 36194 239144 38326 239200
rect 38494 239144 40718 239200
rect 40886 239144 43018 239200
rect 43186 239144 45318 239200
rect 45486 239144 47710 239200
rect 47878 239144 50010 239200
rect 50178 239144 52310 239200
rect 52478 239144 54702 239200
rect 54870 239144 57002 239200
rect 57170 239144 59302 239200
rect 59470 239144 61694 239200
rect 61862 239144 63994 239200
rect 64162 239144 66386 239200
rect 66554 239144 68686 239200
rect 68854 239144 70986 239200
rect 71154 239144 73378 239200
rect 73546 239144 75678 239200
rect 75846 239144 77978 239200
rect 78146 239144 80370 239200
rect 80538 239144 82670 239200
rect 82838 239144 84970 239200
rect 85138 239144 87362 239200
rect 87530 239144 89662 239200
rect 89830 239144 91962 239200
rect 92130 239144 94354 239200
rect 94522 239144 96654 239200
rect 96822 239144 99046 239200
rect 99214 239144 101346 239200
rect 101514 239144 103646 239200
rect 103814 239144 106038 239200
rect 106206 239144 108338 239200
rect 108506 239144 110638 239200
rect 110806 239144 113030 239200
rect 113198 239144 115330 239200
rect 115498 239144 117630 239200
rect 117798 239144 120022 239200
rect 120190 239144 122322 239200
rect 122490 239144 124622 239200
rect 124790 239144 127014 239200
rect 127182 239144 129314 239200
rect 129482 239144 131706 239200
rect 131874 239144 134006 239200
rect 134174 239144 136306 239200
rect 136474 239144 138698 239200
rect 138866 239144 140998 239200
rect 141166 239144 143298 239200
rect 143466 239144 145690 239200
rect 145858 239144 147990 239200
rect 148158 239144 150290 239200
rect 150458 239144 152682 239200
rect 152850 239144 154982 239200
rect 155150 239144 157374 239200
rect 157542 239144 159674 239200
rect 159842 239144 161974 239200
rect 162142 239144 164366 239200
rect 164534 239144 166666 239200
rect 166834 239144 168966 239200
rect 169134 239144 171358 239200
rect 171526 239144 173658 239200
rect 173826 239144 175958 239200
rect 176126 239144 178350 239200
rect 178518 239144 180650 239200
rect 180818 239144 182950 239200
rect 183118 239144 185342 239200
rect 185510 239144 187642 239200
rect 187810 239144 190034 239200
rect 190202 239144 192334 239200
rect 192502 239144 194634 239200
rect 194802 239144 197026 239200
rect 197194 239144 199326 239200
rect 199494 239144 201626 239200
rect 201794 239144 204018 239200
rect 204186 239144 206318 239200
rect 206486 239144 208618 239200
rect 208786 239144 211010 239200
rect 211178 239144 213310 239200
rect 213478 239144 215610 239200
rect 215778 239144 218002 239200
rect 218170 239144 220302 239200
rect 220470 239144 222694 239200
rect 222862 239144 224994 239200
rect 225162 239144 227294 239200
rect 227462 239144 229686 239200
rect 229854 239144 231986 239200
rect 232154 239144 234286 239200
rect 234454 239144 236678 239200
rect 236846 239144 238978 239200
rect 239146 239144 241278 239200
rect 241446 239144 243670 239200
rect 243838 239144 245970 239200
rect 246138 239144 248270 239200
rect 248438 239144 250662 239200
rect 250830 239144 252962 239200
rect 253130 239144 255354 239200
rect 255522 239144 257654 239200
rect 257822 239144 259954 239200
rect 260122 239144 262346 239200
rect 262514 239144 264646 239200
rect 264814 239144 266946 239200
rect 267114 239144 269338 239200
rect 269506 239144 271638 239200
rect 271806 239144 273938 239200
rect 274106 239144 276330 239200
rect 276498 239144 278630 239200
rect 278798 239144 279662 239200
rect 294 856 279662 239144
rect 406 800 790 856
rect 958 800 1342 856
rect 1510 800 1894 856
rect 2062 800 2446 856
rect 2614 800 2998 856
rect 3166 800 3550 856
rect 3718 800 4102 856
rect 4270 800 4654 856
rect 4822 800 5206 856
rect 5374 800 5758 856
rect 5926 800 6310 856
rect 6478 800 6862 856
rect 7030 800 7414 856
rect 7582 800 8058 856
rect 8226 800 8610 856
rect 8778 800 9162 856
rect 9330 800 9714 856
rect 9882 800 10266 856
rect 10434 800 10818 856
rect 10986 800 11370 856
rect 11538 800 11922 856
rect 12090 800 12474 856
rect 12642 800 13026 856
rect 13194 800 13578 856
rect 13746 800 14130 856
rect 14298 800 14682 856
rect 14850 800 15234 856
rect 15402 800 15878 856
rect 16046 800 16430 856
rect 16598 800 16982 856
rect 17150 800 17534 856
rect 17702 800 18086 856
rect 18254 800 18638 856
rect 18806 800 19190 856
rect 19358 800 19742 856
rect 19910 800 20294 856
rect 20462 800 20846 856
rect 21014 800 21398 856
rect 21566 800 21950 856
rect 22118 800 22502 856
rect 22670 800 23146 856
rect 23314 800 23698 856
rect 23866 800 24250 856
rect 24418 800 24802 856
rect 24970 800 25354 856
rect 25522 800 25906 856
rect 26074 800 26458 856
rect 26626 800 27010 856
rect 27178 800 27562 856
rect 27730 800 28114 856
rect 28282 800 28666 856
rect 28834 800 29218 856
rect 29386 800 29770 856
rect 29938 800 30322 856
rect 30490 800 30966 856
rect 31134 800 31518 856
rect 31686 800 32070 856
rect 32238 800 32622 856
rect 32790 800 33174 856
rect 33342 800 33726 856
rect 33894 800 34278 856
rect 34446 800 34830 856
rect 34998 800 35382 856
rect 35550 800 35934 856
rect 36102 800 36486 856
rect 36654 800 37038 856
rect 37206 800 37590 856
rect 37758 800 38234 856
rect 38402 800 38786 856
rect 38954 800 39338 856
rect 39506 800 39890 856
rect 40058 800 40442 856
rect 40610 800 40994 856
rect 41162 800 41546 856
rect 41714 800 42098 856
rect 42266 800 42650 856
rect 42818 800 43202 856
rect 43370 800 43754 856
rect 43922 800 44306 856
rect 44474 800 44858 856
rect 45026 800 45410 856
rect 45578 800 46054 856
rect 46222 800 46606 856
rect 46774 800 47158 856
rect 47326 800 47710 856
rect 47878 800 48262 856
rect 48430 800 48814 856
rect 48982 800 49366 856
rect 49534 800 49918 856
rect 50086 800 50470 856
rect 50638 800 51022 856
rect 51190 800 51574 856
rect 51742 800 52126 856
rect 52294 800 52678 856
rect 52846 800 53322 856
rect 53490 800 53874 856
rect 54042 800 54426 856
rect 54594 800 54978 856
rect 55146 800 55530 856
rect 55698 800 56082 856
rect 56250 800 56634 856
rect 56802 800 57186 856
rect 57354 800 57738 856
rect 57906 800 58290 856
rect 58458 800 58842 856
rect 59010 800 59394 856
rect 59562 800 59946 856
rect 60114 800 60498 856
rect 60666 800 61142 856
rect 61310 800 61694 856
rect 61862 800 62246 856
rect 62414 800 62798 856
rect 62966 800 63350 856
rect 63518 800 63902 856
rect 64070 800 64454 856
rect 64622 800 65006 856
rect 65174 800 65558 856
rect 65726 800 66110 856
rect 66278 800 66662 856
rect 66830 800 67214 856
rect 67382 800 67766 856
rect 67934 800 68410 856
rect 68578 800 68962 856
rect 69130 800 69514 856
rect 69682 800 70066 856
rect 70234 800 70618 856
rect 70786 800 71170 856
rect 71338 800 71722 856
rect 71890 800 72274 856
rect 72442 800 72826 856
rect 72994 800 73378 856
rect 73546 800 73930 856
rect 74098 800 74482 856
rect 74650 800 75034 856
rect 75202 800 75586 856
rect 75754 800 76230 856
rect 76398 800 76782 856
rect 76950 800 77334 856
rect 77502 800 77886 856
rect 78054 800 78438 856
rect 78606 800 78990 856
rect 79158 800 79542 856
rect 79710 800 80094 856
rect 80262 800 80646 856
rect 80814 800 81198 856
rect 81366 800 81750 856
rect 81918 800 82302 856
rect 82470 800 82854 856
rect 83022 800 83498 856
rect 83666 800 84050 856
rect 84218 800 84602 856
rect 84770 800 85154 856
rect 85322 800 85706 856
rect 85874 800 86258 856
rect 86426 800 86810 856
rect 86978 800 87362 856
rect 87530 800 87914 856
rect 88082 800 88466 856
rect 88634 800 89018 856
rect 89186 800 89570 856
rect 89738 800 90122 856
rect 90290 800 90674 856
rect 90842 800 91318 856
rect 91486 800 91870 856
rect 92038 800 92422 856
rect 92590 800 92974 856
rect 93142 800 93526 856
rect 93694 800 94078 856
rect 94246 800 94630 856
rect 94798 800 95182 856
rect 95350 800 95734 856
rect 95902 800 96286 856
rect 96454 800 96838 856
rect 97006 800 97390 856
rect 97558 800 97942 856
rect 98110 800 98494 856
rect 98662 800 99138 856
rect 99306 800 99690 856
rect 99858 800 100242 856
rect 100410 800 100794 856
rect 100962 800 101346 856
rect 101514 800 101898 856
rect 102066 800 102450 856
rect 102618 800 103002 856
rect 103170 800 103554 856
rect 103722 800 104106 856
rect 104274 800 104658 856
rect 104826 800 105210 856
rect 105378 800 105762 856
rect 105930 800 106406 856
rect 106574 800 106958 856
rect 107126 800 107510 856
rect 107678 800 108062 856
rect 108230 800 108614 856
rect 108782 800 109166 856
rect 109334 800 109718 856
rect 109886 800 110270 856
rect 110438 800 110822 856
rect 110990 800 111374 856
rect 111542 800 111926 856
rect 112094 800 112478 856
rect 112646 800 113030 856
rect 113198 800 113582 856
rect 113750 800 114226 856
rect 114394 800 114778 856
rect 114946 800 115330 856
rect 115498 800 115882 856
rect 116050 800 116434 856
rect 116602 800 116986 856
rect 117154 800 117538 856
rect 117706 800 118090 856
rect 118258 800 118642 856
rect 118810 800 119194 856
rect 119362 800 119746 856
rect 119914 800 120298 856
rect 120466 800 120850 856
rect 121018 800 121494 856
rect 121662 800 122046 856
rect 122214 800 122598 856
rect 122766 800 123150 856
rect 123318 800 123702 856
rect 123870 800 124254 856
rect 124422 800 124806 856
rect 124974 800 125358 856
rect 125526 800 125910 856
rect 126078 800 126462 856
rect 126630 800 127014 856
rect 127182 800 127566 856
rect 127734 800 128118 856
rect 128286 800 128670 856
rect 128838 800 129314 856
rect 129482 800 129866 856
rect 130034 800 130418 856
rect 130586 800 130970 856
rect 131138 800 131522 856
rect 131690 800 132074 856
rect 132242 800 132626 856
rect 132794 800 133178 856
rect 133346 800 133730 856
rect 133898 800 134282 856
rect 134450 800 134834 856
rect 135002 800 135386 856
rect 135554 800 135938 856
rect 136106 800 136582 856
rect 136750 800 137134 856
rect 137302 800 137686 856
rect 137854 800 138238 856
rect 138406 800 138790 856
rect 138958 800 139342 856
rect 139510 800 139894 856
rect 140062 800 140446 856
rect 140614 800 140998 856
rect 141166 800 141550 856
rect 141718 800 142102 856
rect 142270 800 142654 856
rect 142822 800 143206 856
rect 143374 800 143758 856
rect 143926 800 144402 856
rect 144570 800 144954 856
rect 145122 800 145506 856
rect 145674 800 146058 856
rect 146226 800 146610 856
rect 146778 800 147162 856
rect 147330 800 147714 856
rect 147882 800 148266 856
rect 148434 800 148818 856
rect 148986 800 149370 856
rect 149538 800 149922 856
rect 150090 800 150474 856
rect 150642 800 151026 856
rect 151194 800 151670 856
rect 151838 800 152222 856
rect 152390 800 152774 856
rect 152942 800 153326 856
rect 153494 800 153878 856
rect 154046 800 154430 856
rect 154598 800 154982 856
rect 155150 800 155534 856
rect 155702 800 156086 856
rect 156254 800 156638 856
rect 156806 800 157190 856
rect 157358 800 157742 856
rect 157910 800 158294 856
rect 158462 800 158846 856
rect 159014 800 159490 856
rect 159658 800 160042 856
rect 160210 800 160594 856
rect 160762 800 161146 856
rect 161314 800 161698 856
rect 161866 800 162250 856
rect 162418 800 162802 856
rect 162970 800 163354 856
rect 163522 800 163906 856
rect 164074 800 164458 856
rect 164626 800 165010 856
rect 165178 800 165562 856
rect 165730 800 166114 856
rect 166282 800 166758 856
rect 166926 800 167310 856
rect 167478 800 167862 856
rect 168030 800 168414 856
rect 168582 800 168966 856
rect 169134 800 169518 856
rect 169686 800 170070 856
rect 170238 800 170622 856
rect 170790 800 171174 856
rect 171342 800 171726 856
rect 171894 800 172278 856
rect 172446 800 172830 856
rect 172998 800 173382 856
rect 173550 800 173934 856
rect 174102 800 174578 856
rect 174746 800 175130 856
rect 175298 800 175682 856
rect 175850 800 176234 856
rect 176402 800 176786 856
rect 176954 800 177338 856
rect 177506 800 177890 856
rect 178058 800 178442 856
rect 178610 800 178994 856
rect 179162 800 179546 856
rect 179714 800 180098 856
rect 180266 800 180650 856
rect 180818 800 181202 856
rect 181370 800 181846 856
rect 182014 800 182398 856
rect 182566 800 182950 856
rect 183118 800 183502 856
rect 183670 800 184054 856
rect 184222 800 184606 856
rect 184774 800 185158 856
rect 185326 800 185710 856
rect 185878 800 186262 856
rect 186430 800 186814 856
rect 186982 800 187366 856
rect 187534 800 187918 856
rect 188086 800 188470 856
rect 188638 800 189022 856
rect 189190 800 189666 856
rect 189834 800 190218 856
rect 190386 800 190770 856
rect 190938 800 191322 856
rect 191490 800 191874 856
rect 192042 800 192426 856
rect 192594 800 192978 856
rect 193146 800 193530 856
rect 193698 800 194082 856
rect 194250 800 194634 856
rect 194802 800 195186 856
rect 195354 800 195738 856
rect 195906 800 196290 856
rect 196458 800 196842 856
rect 197010 800 197486 856
rect 197654 800 198038 856
rect 198206 800 198590 856
rect 198758 800 199142 856
rect 199310 800 199694 856
rect 199862 800 200246 856
rect 200414 800 200798 856
rect 200966 800 201350 856
rect 201518 800 201902 856
rect 202070 800 202454 856
rect 202622 800 203006 856
rect 203174 800 203558 856
rect 203726 800 204110 856
rect 204278 800 204754 856
rect 204922 800 205306 856
rect 205474 800 205858 856
rect 206026 800 206410 856
rect 206578 800 206962 856
rect 207130 800 207514 856
rect 207682 800 208066 856
rect 208234 800 208618 856
rect 208786 800 209170 856
rect 209338 800 209722 856
rect 209890 800 210274 856
rect 210442 800 210826 856
rect 210994 800 211378 856
rect 211546 800 211930 856
rect 212098 800 212574 856
rect 212742 800 213126 856
rect 213294 800 213678 856
rect 213846 800 214230 856
rect 214398 800 214782 856
rect 214950 800 215334 856
rect 215502 800 215886 856
rect 216054 800 216438 856
rect 216606 800 216990 856
rect 217158 800 217542 856
rect 217710 800 218094 856
rect 218262 800 218646 856
rect 218814 800 219198 856
rect 219366 800 219842 856
rect 220010 800 220394 856
rect 220562 800 220946 856
rect 221114 800 221498 856
rect 221666 800 222050 856
rect 222218 800 222602 856
rect 222770 800 223154 856
rect 223322 800 223706 856
rect 223874 800 224258 856
rect 224426 800 224810 856
rect 224978 800 225362 856
rect 225530 800 225914 856
rect 226082 800 226466 856
rect 226634 800 227018 856
rect 227186 800 227662 856
rect 227830 800 228214 856
rect 228382 800 228766 856
rect 228934 800 229318 856
rect 229486 800 229870 856
rect 230038 800 230422 856
rect 230590 800 230974 856
rect 231142 800 231526 856
rect 231694 800 232078 856
rect 232246 800 232630 856
rect 232798 800 233182 856
rect 233350 800 233734 856
rect 233902 800 234286 856
rect 234454 800 234930 856
rect 235098 800 235482 856
rect 235650 800 236034 856
rect 236202 800 236586 856
rect 236754 800 237138 856
rect 237306 800 237690 856
rect 237858 800 238242 856
rect 238410 800 238794 856
rect 238962 800 239346 856
rect 239514 800 239898 856
rect 240066 800 240450 856
rect 240618 800 241002 856
rect 241170 800 241554 856
rect 241722 800 242106 856
rect 242274 800 242750 856
rect 242918 800 243302 856
rect 243470 800 243854 856
rect 244022 800 244406 856
rect 244574 800 244958 856
rect 245126 800 245510 856
rect 245678 800 246062 856
rect 246230 800 246614 856
rect 246782 800 247166 856
rect 247334 800 247718 856
rect 247886 800 248270 856
rect 248438 800 248822 856
rect 248990 800 249374 856
rect 249542 800 250018 856
rect 250186 800 250570 856
rect 250738 800 251122 856
rect 251290 800 251674 856
rect 251842 800 252226 856
rect 252394 800 252778 856
rect 252946 800 253330 856
rect 253498 800 253882 856
rect 254050 800 254434 856
rect 254602 800 254986 856
rect 255154 800 255538 856
rect 255706 800 256090 856
rect 256258 800 256642 856
rect 256810 800 257194 856
rect 257362 800 257838 856
rect 258006 800 258390 856
rect 258558 800 258942 856
rect 259110 800 259494 856
rect 259662 800 260046 856
rect 260214 800 260598 856
rect 260766 800 261150 856
rect 261318 800 261702 856
rect 261870 800 262254 856
rect 262422 800 262806 856
rect 262974 800 263358 856
rect 263526 800 263910 856
rect 264078 800 264462 856
rect 264630 800 265106 856
rect 265274 800 265658 856
rect 265826 800 266210 856
rect 266378 800 266762 856
rect 266930 800 267314 856
rect 267482 800 267866 856
rect 268034 800 268418 856
rect 268586 800 268970 856
rect 269138 800 269522 856
rect 269690 800 270074 856
rect 270242 800 270626 856
rect 270794 800 271178 856
rect 271346 800 271730 856
rect 271898 800 272282 856
rect 272450 800 272926 856
rect 273094 800 273478 856
rect 273646 800 274030 856
rect 274198 800 274582 856
rect 274750 800 275134 856
rect 275302 800 275686 856
rect 275854 800 276238 856
rect 276406 800 276790 856
rect 276958 800 277342 856
rect 277510 800 277894 856
rect 278062 800 278446 856
rect 278614 800 278998 856
rect 279166 800 279550 856
<< metal3 >>
rect 0 224952 800 225072
rect 279200 219920 280000 220040
rect 0 194896 800 195016
rect 279200 179936 280000 180056
rect 0 164976 800 165096
rect 279200 139952 280000 140072
rect 0 134920 800 135040
rect 0 104864 800 104984
rect 279200 99968 280000 100088
rect 0 74944 800 75064
rect 279200 59984 280000 60104
rect 0 44888 800 45008
rect 279200 20000 280000 20120
rect 0 14968 800 15088
<< obsm3 >>
rect 289 225152 279667 237761
rect 880 224872 279667 225152
rect 289 220120 279667 224872
rect 289 219840 279120 220120
rect 289 195096 279667 219840
rect 880 194816 279667 195096
rect 289 180136 279667 194816
rect 289 179856 279120 180136
rect 289 165176 279667 179856
rect 880 164896 279667 165176
rect 289 140152 279667 164896
rect 289 139872 279120 140152
rect 289 135120 279667 139872
rect 880 134840 279667 135120
rect 289 105064 279667 134840
rect 880 104784 279667 105064
rect 289 100168 279667 104784
rect 289 99888 279120 100168
rect 289 75144 279667 99888
rect 880 74864 279667 75144
rect 289 60184 279667 74864
rect 289 59904 279120 60184
rect 289 45088 279667 59904
rect 880 44808 279667 45088
rect 289 20200 279667 44808
rect 289 19920 279120 20200
rect 289 15168 279667 19920
rect 880 14888 279667 15168
rect 289 2143 279667 14888
<< metal4 >>
rect 4208 2128 4528 237776
rect 19568 2128 19888 237776
rect 34928 2128 35248 237776
rect 50288 2128 50608 237776
rect 65648 2128 65968 237776
rect 81008 2128 81328 237776
rect 96368 2128 96688 237776
rect 111728 2128 112048 237776
rect 127088 2128 127408 237776
rect 142448 2128 142768 237776
rect 157808 2128 158128 237776
rect 173168 2128 173488 237776
rect 188528 2128 188848 237776
rect 203888 2128 204208 237776
rect 219248 2128 219568 237776
rect 234608 2128 234928 237776
rect 249968 2128 250288 237776
rect 265328 2128 265648 237776
<< obsm4 >>
rect 64091 144875 65568 212533
rect 66048 144875 80928 212533
rect 81408 144875 96288 212533
rect 96768 144875 111648 212533
rect 112128 144875 127008 212533
rect 127488 144875 142368 212533
rect 142848 144875 157728 212533
rect 158208 144875 165909 212533
<< labels >>
rlabel metal2 s 267002 239200 267058 240000 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 0 74944 800 75064 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 276846 0 276902 800 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 271694 239200 271750 240000 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 273994 239200 274050 240000 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 276386 239200 276442 240000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 0 104864 800 104984 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal3 s 279200 59984 280000 60104 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 277398 0 277454 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 277950 0 278006 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 278502 0 278558 800 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 274086 0 274142 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 279200 99968 280000 100088 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 134920 800 135040 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 279200 139952 280000 140072 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 279054 0 279110 800 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 164976 800 165096 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 279606 0 279662 800 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 194896 800 195016 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal2 s 278686 239200 278742 240000 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 279200 179936 280000 180056 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 279200 219920 280000 220040 6 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal2 s 274638 0 274694 800 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s 0 224952 800 225072 6 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal2 s 275190 0 275246 800 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 279200 20000 280000 20120 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal3 s 0 14968 800 15088 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal3 s 0 44888 800 45008 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal2 s 275742 0 275798 800 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal2 s 276294 0 276350 800 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 269394 239200 269450 240000 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 1122 239200 1178 240000 6 io_in[0]
port 32 nsew signal input
rlabel metal2 s 71042 239200 71098 240000 6 io_in[10]
port 33 nsew signal input
rlabel metal2 s 78034 239200 78090 240000 6 io_in[11]
port 34 nsew signal input
rlabel metal2 s 85026 239200 85082 240000 6 io_in[12]
port 35 nsew signal input
rlabel metal2 s 92018 239200 92074 240000 6 io_in[13]
port 36 nsew signal input
rlabel metal2 s 99102 239200 99158 240000 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 106094 239200 106150 240000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 113086 239200 113142 240000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 120078 239200 120134 240000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 127070 239200 127126 240000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 134062 239200 134118 240000 6 io_in[19]
port 42 nsew signal input
rlabel metal2 s 8114 239200 8170 240000 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 141054 239200 141110 240000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 148046 239200 148102 240000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 155038 239200 155094 240000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 162030 239200 162086 240000 6 io_in[23]
port 47 nsew signal input
rlabel metal2 s 169022 239200 169078 240000 6 io_in[24]
port 48 nsew signal input
rlabel metal2 s 176014 239200 176070 240000 6 io_in[25]
port 49 nsew signal input
rlabel metal2 s 183006 239200 183062 240000 6 io_in[26]
port 50 nsew signal input
rlabel metal2 s 190090 239200 190146 240000 6 io_in[27]
port 51 nsew signal input
rlabel metal2 s 197082 239200 197138 240000 6 io_in[28]
port 52 nsew signal input
rlabel metal2 s 204074 239200 204130 240000 6 io_in[29]
port 53 nsew signal input
rlabel metal2 s 15106 239200 15162 240000 6 io_in[2]
port 54 nsew signal input
rlabel metal2 s 211066 239200 211122 240000 6 io_in[30]
port 55 nsew signal input
rlabel metal2 s 218058 239200 218114 240000 6 io_in[31]
port 56 nsew signal input
rlabel metal2 s 225050 239200 225106 240000 6 io_in[32]
port 57 nsew signal input
rlabel metal2 s 232042 239200 232098 240000 6 io_in[33]
port 58 nsew signal input
rlabel metal2 s 239034 239200 239090 240000 6 io_in[34]
port 59 nsew signal input
rlabel metal2 s 246026 239200 246082 240000 6 io_in[35]
port 60 nsew signal input
rlabel metal2 s 253018 239200 253074 240000 6 io_in[36]
port 61 nsew signal input
rlabel metal2 s 260010 239200 260066 240000 6 io_in[37]
port 62 nsew signal input
rlabel metal2 s 22098 239200 22154 240000 6 io_in[3]
port 63 nsew signal input
rlabel metal2 s 29090 239200 29146 240000 6 io_in[4]
port 64 nsew signal input
rlabel metal2 s 36082 239200 36138 240000 6 io_in[5]
port 65 nsew signal input
rlabel metal2 s 43074 239200 43130 240000 6 io_in[6]
port 66 nsew signal input
rlabel metal2 s 50066 239200 50122 240000 6 io_in[7]
port 67 nsew signal input
rlabel metal2 s 57058 239200 57114 240000 6 io_in[8]
port 68 nsew signal input
rlabel metal2 s 64050 239200 64106 240000 6 io_in[9]
port 69 nsew signal input
rlabel metal2 s 3422 239200 3478 240000 6 io_oeb[0]
port 70 nsew signal output
rlabel metal2 s 73434 239200 73490 240000 6 io_oeb[10]
port 71 nsew signal output
rlabel metal2 s 80426 239200 80482 240000 6 io_oeb[11]
port 72 nsew signal output
rlabel metal2 s 87418 239200 87474 240000 6 io_oeb[12]
port 73 nsew signal output
rlabel metal2 s 94410 239200 94466 240000 6 io_oeb[13]
port 74 nsew signal output
rlabel metal2 s 101402 239200 101458 240000 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 108394 239200 108450 240000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 115386 239200 115442 240000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 122378 239200 122434 240000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 129370 239200 129426 240000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 136362 239200 136418 240000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal2 s 10414 239200 10470 240000 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 143354 239200 143410 240000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 150346 239200 150402 240000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 157430 239200 157486 240000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 164422 239200 164478 240000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal2 s 171414 239200 171470 240000 6 io_oeb[24]
port 86 nsew signal output
rlabel metal2 s 178406 239200 178462 240000 6 io_oeb[25]
port 87 nsew signal output
rlabel metal2 s 185398 239200 185454 240000 6 io_oeb[26]
port 88 nsew signal output
rlabel metal2 s 192390 239200 192446 240000 6 io_oeb[27]
port 89 nsew signal output
rlabel metal2 s 199382 239200 199438 240000 6 io_oeb[28]
port 90 nsew signal output
rlabel metal2 s 206374 239200 206430 240000 6 io_oeb[29]
port 91 nsew signal output
rlabel metal2 s 17406 239200 17462 240000 6 io_oeb[2]
port 92 nsew signal output
rlabel metal2 s 213366 239200 213422 240000 6 io_oeb[30]
port 93 nsew signal output
rlabel metal2 s 220358 239200 220414 240000 6 io_oeb[31]
port 94 nsew signal output
rlabel metal2 s 227350 239200 227406 240000 6 io_oeb[32]
port 95 nsew signal output
rlabel metal2 s 234342 239200 234398 240000 6 io_oeb[33]
port 96 nsew signal output
rlabel metal2 s 241334 239200 241390 240000 6 io_oeb[34]
port 97 nsew signal output
rlabel metal2 s 248326 239200 248382 240000 6 io_oeb[35]
port 98 nsew signal output
rlabel metal2 s 255410 239200 255466 240000 6 io_oeb[36]
port 99 nsew signal output
rlabel metal2 s 262402 239200 262458 240000 6 io_oeb[37]
port 100 nsew signal output
rlabel metal2 s 24398 239200 24454 240000 6 io_oeb[3]
port 101 nsew signal output
rlabel metal2 s 31390 239200 31446 240000 6 io_oeb[4]
port 102 nsew signal output
rlabel metal2 s 38382 239200 38438 240000 6 io_oeb[5]
port 103 nsew signal output
rlabel metal2 s 45374 239200 45430 240000 6 io_oeb[6]
port 104 nsew signal output
rlabel metal2 s 52366 239200 52422 240000 6 io_oeb[7]
port 105 nsew signal output
rlabel metal2 s 59358 239200 59414 240000 6 io_oeb[8]
port 106 nsew signal output
rlabel metal2 s 66442 239200 66498 240000 6 io_oeb[9]
port 107 nsew signal output
rlabel metal2 s 5722 239200 5778 240000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 75734 239200 75790 240000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 82726 239200 82782 240000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 89718 239200 89774 240000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 96710 239200 96766 240000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 103702 239200 103758 240000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 110694 239200 110750 240000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 117686 239200 117742 240000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 124678 239200 124734 240000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 131762 239200 131818 240000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 138754 239200 138810 240000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 12714 239200 12770 240000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 145746 239200 145802 240000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 152738 239200 152794 240000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 159730 239200 159786 240000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 166722 239200 166778 240000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 173714 239200 173770 240000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 180706 239200 180762 240000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 187698 239200 187754 240000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 194690 239200 194746 240000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 201682 239200 201738 240000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 208674 239200 208730 240000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 19706 239200 19762 240000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 215666 239200 215722 240000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 222750 239200 222806 240000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 229742 239200 229798 240000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 236734 239200 236790 240000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 243726 239200 243782 240000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 250718 239200 250774 240000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 257710 239200 257766 240000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 264702 239200 264758 240000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 26698 239200 26754 240000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 33782 239200 33838 240000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 40774 239200 40830 240000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 47766 239200 47822 240000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 54758 239200 54814 240000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 61750 239200 61806 240000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 68742 239200 68798 240000 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 227074 0 227130 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 230478 0 230534 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 235538 0 235594 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 237194 0 237250 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 240506 0 240562 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 242162 0 242218 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 243910 0 243966 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 247222 0 247278 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 248878 0 248934 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 250626 0 250682 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 252282 0 252338 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 253938 0 253994 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 255594 0 255650 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 258998 0 259054 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 260654 0 260710 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 262310 0 262366 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 263966 0 264022 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 265714 0 265770 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 267370 0 267426 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 269026 0 269082 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 270682 0 270738 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 272338 0 272394 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 186870 0 186926 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 193586 0 193642 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 198646 0 198702 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 201958 0 202014 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 205362 0 205418 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 213734 0 213790 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 223762 0 223818 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 227718 0 227774 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 229374 0 229430 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 231030 0 231086 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 232686 0 232742 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 234342 0 234398 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 236090 0 236146 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 237746 0 237802 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 239402 0 239458 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 241058 0 241114 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 242806 0 242862 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 244462 0 244518 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 246118 0 246174 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 247774 0 247830 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 249430 0 249486 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 251178 0 251234 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 252834 0 252890 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 254490 0 254546 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 256146 0 256202 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 257894 0 257950 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 259550 0 259606 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 261206 0 261262 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 262862 0 262918 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 264518 0 264574 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 266266 0 266322 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 267922 0 267978 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 269578 0 269634 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 271234 0 271290 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 272982 0 273038 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 108670 0 108726 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 110326 0 110382 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 120354 0 120410 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 133786 0 133842 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 167366 0 167422 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 169022 0 169078 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 172334 0 172390 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 173990 0 174046 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 177394 0 177450 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 179050 0 179106 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 180706 0 180762 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 182454 0 182510 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 184110 0 184166 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 185766 0 185822 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 187422 0 187478 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 189078 0 189134 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 190826 0 190882 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 192482 0 192538 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 194138 0 194194 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 197542 0 197598 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 200854 0 200910 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 202510 0 202566 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 205914 0 205970 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 207570 0 207626 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 209226 0 209282 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 212630 0 212686 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 214286 0 214342 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 215942 0 215998 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 217598 0 217654 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 219254 0 219310 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 221002 0 221058 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 222658 0 222714 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 224314 0 224370 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 225970 0 226026 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 234986 0 235042 800 6 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 238298 0 238354 800 6 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 239954 0 240010 800 6 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 241610 0 241666 800 6 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 245014 0 245070 800 6 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 248326 0 248382 800 6 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 250074 0 250130 800 6 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 251730 0 251786 800 6 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 255042 0 255098 800 6 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 256698 0 256754 800 6 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 258446 0 258502 800 6 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 261758 0 261814 800 6 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 263414 0 263470 800 6 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 265162 0 265218 800 6 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 266818 0 266874 800 6 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 268474 0 268530 800 6 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 270130 0 270186 800 6 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 271786 0 271842 800 6 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 273534 0 273590 800 6 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 181258 0 181314 800 6 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 183006 0 183062 800 6 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 184662 0 184718 800 6 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 187974 0 188030 800 6 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 189722 0 189778 800 6 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 194690 0 194746 800 6 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 196346 0 196402 800 6 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 201406 0 201462 800 6 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 206466 0 206522 800 6 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 208122 0 208178 800 6 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 211434 0 211490 800 6 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 214838 0 214894 800 6 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 218150 0 218206 800 6 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 223210 0 223266 800 6 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 224866 0 224922 800 6 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 226522 0 226578 800 6 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 530 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 531 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 532 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 wbs_adr_i[0]
port 533 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[10]
port 534 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_adr_i[11]
port 535 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[12]
port 536 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_adr_i[13]
port 537 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[14]
port 538 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[15]
port 539 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_adr_i[16]
port 540 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_adr_i[17]
port 541 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_adr_i[18]
port 542 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[19]
port 543 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[1]
port 544 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_adr_i[20]
port 545 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_adr_i[21]
port 546 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 wbs_adr_i[22]
port 547 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 wbs_adr_i[23]
port 548 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wbs_adr_i[24]
port 549 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 wbs_adr_i[25]
port 550 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_adr_i[26]
port 551 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_adr_i[27]
port 552 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_adr_i[28]
port 553 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 wbs_adr_i[29]
port 554 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[2]
port 555 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 wbs_adr_i[30]
port 556 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 wbs_adr_i[31]
port 557 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[3]
port 558 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[4]
port 559 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[5]
port 560 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[6]
port 561 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[7]
port 562 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[8]
port 563 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[9]
port 564 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_cyc_i
port 565 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_i[0]
port 566 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[10]
port 567 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[11]
port 568 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_i[12]
port 569 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_i[13]
port 570 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_i[14]
port 571 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[15]
port 572 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[16]
port 573 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_i[17]
port 574 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_i[18]
port 575 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[19]
port 576 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_i[1]
port 577 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_i[20]
port 578 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_i[21]
port 579 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_dat_i[22]
port 580 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_i[23]
port 581 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_i[24]
port 582 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[25]
port 583 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wbs_dat_i[26]
port 584 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_i[27]
port 585 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_i[28]
port 586 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_i[29]
port 587 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_i[2]
port 588 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_i[30]
port 589 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_i[31]
port 590 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[3]
port 591 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[4]
port 592 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_i[5]
port 593 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[6]
port 594 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[7]
port 595 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[8]
port 596 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[9]
port 597 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_o[0]
port 598 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_o[10]
port 599 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[11]
port 600 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_o[12]
port 601 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[13]
port 602 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[14]
port 603 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[15]
port 604 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[16]
port 605 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_o[17]
port 606 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_o[18]
port 607 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_o[19]
port 608 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_o[1]
port 609 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_o[20]
port 610 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_o[21]
port 611 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 wbs_dat_o[22]
port 612 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_o[23]
port 613 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 wbs_dat_o[24]
port 614 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 wbs_dat_o[25]
port 615 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_o[26]
port 616 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_o[27]
port 617 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_o[28]
port 618 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 wbs_dat_o[29]
port 619 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[2]
port 620 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_o[30]
port 621 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_o[31]
port 622 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[3]
port 623 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_o[4]
port 624 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[5]
port 625 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[6]
port 626 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[7]
port 627 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[8]
port 628 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[9]
port 629 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 wbs_sel_i[0]
port 630 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_sel_i[1]
port 631 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_sel_i[2]
port 632 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_sel_i[3]
port 633 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_stb_i
port 634 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_we_i
port 635 nsew signal input
rlabel metal4 s 249968 2128 250288 237776 6 VPWR
port 636 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 237776 6 VPWR
port 637 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 237776 6 VPWR
port 638 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 237776 6 VPWR
port 639 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 237776 6 VPWR
port 640 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 237776 6 VPWR
port 641 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 237776 6 VPWR
port 642 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 237776 6 VPWR
port 643 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 237776 6 VPWR
port 644 nsew power bidirectional
rlabel metal4 s 265328 2128 265648 237776 6 VGND
port 645 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 237776 6 VGND
port 646 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 237776 6 VGND
port 647 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 237776 6 VGND
port 648 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 237776 6 VGND
port 649 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 237776 6 VGND
port 650 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 237776 6 VGND
port 651 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 237776 6 VGND
port 652 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 237776 6 VGND
port 653 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 280000 240000
string LEFview TRUE
<< end >>
