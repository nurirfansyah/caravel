magic
tech sky130A
magscale 1 2
timestamp 1608262846
<< obsli1 >>
rect 1104 2159 278852 237745
<< obsm1 >>
rect 290 1912 279114 237776
<< metal2 >>
rect 1122 239200 1178 240000
rect 3330 239200 3386 240000
rect 5630 239200 5686 240000
rect 7930 239200 7986 240000
rect 10138 239200 10194 240000
rect 12438 239200 12494 240000
rect 14738 239200 14794 240000
rect 17038 239200 17094 240000
rect 19246 239200 19302 240000
rect 21546 239200 21602 240000
rect 23846 239200 23902 240000
rect 26146 239200 26202 240000
rect 28354 239200 28410 240000
rect 30654 239200 30710 240000
rect 32954 239200 33010 240000
rect 35254 239200 35310 240000
rect 37462 239200 37518 240000
rect 39762 239200 39818 240000
rect 42062 239200 42118 240000
rect 44362 239200 44418 240000
rect 46570 239200 46626 240000
rect 48870 239200 48926 240000
rect 51170 239200 51226 240000
rect 53470 239200 53526 240000
rect 55678 239200 55734 240000
rect 57978 239200 58034 240000
rect 60278 239200 60334 240000
rect 62486 239200 62542 240000
rect 64786 239200 64842 240000
rect 67086 239200 67142 240000
rect 69386 239200 69442 240000
rect 71594 239200 71650 240000
rect 73894 239200 73950 240000
rect 76194 239200 76250 240000
rect 78494 239200 78550 240000
rect 80702 239200 80758 240000
rect 83002 239200 83058 240000
rect 85302 239200 85358 240000
rect 87602 239200 87658 240000
rect 89810 239200 89866 240000
rect 92110 239200 92166 240000
rect 94410 239200 94466 240000
rect 96710 239200 96766 240000
rect 98918 239200 98974 240000
rect 101218 239200 101274 240000
rect 103518 239200 103574 240000
rect 105818 239200 105874 240000
rect 108026 239200 108082 240000
rect 110326 239200 110382 240000
rect 112626 239200 112682 240000
rect 114834 239200 114890 240000
rect 117134 239200 117190 240000
rect 119434 239200 119490 240000
rect 121734 239200 121790 240000
rect 123942 239200 123998 240000
rect 126242 239200 126298 240000
rect 128542 239200 128598 240000
rect 130842 239200 130898 240000
rect 133050 239200 133106 240000
rect 135350 239200 135406 240000
rect 137650 239200 137706 240000
rect 139950 239200 140006 240000
rect 142158 239200 142214 240000
rect 144458 239200 144514 240000
rect 146758 239200 146814 240000
rect 149058 239200 149114 240000
rect 151266 239200 151322 240000
rect 153566 239200 153622 240000
rect 155866 239200 155922 240000
rect 158166 239200 158222 240000
rect 160374 239200 160430 240000
rect 162674 239200 162730 240000
rect 164974 239200 165030 240000
rect 167274 239200 167330 240000
rect 169482 239200 169538 240000
rect 171782 239200 171838 240000
rect 174082 239200 174138 240000
rect 176290 239200 176346 240000
rect 178590 239200 178646 240000
rect 180890 239200 180946 240000
rect 183190 239200 183246 240000
rect 185398 239200 185454 240000
rect 187698 239200 187754 240000
rect 189998 239200 190054 240000
rect 192298 239200 192354 240000
rect 194506 239200 194562 240000
rect 196806 239200 196862 240000
rect 199106 239200 199162 240000
rect 201406 239200 201462 240000
rect 203614 239200 203670 240000
rect 205914 239200 205970 240000
rect 208214 239200 208270 240000
rect 210514 239200 210570 240000
rect 212722 239200 212778 240000
rect 215022 239200 215078 240000
rect 217322 239200 217378 240000
rect 219622 239200 219678 240000
rect 221830 239200 221886 240000
rect 224130 239200 224186 240000
rect 226430 239200 226486 240000
rect 228638 239200 228694 240000
rect 230938 239200 230994 240000
rect 233238 239200 233294 240000
rect 235538 239200 235594 240000
rect 237746 239200 237802 240000
rect 240046 239200 240102 240000
rect 242346 239200 242402 240000
rect 244646 239200 244702 240000
rect 246854 239200 246910 240000
rect 249154 239200 249210 240000
rect 251454 239200 251510 240000
rect 253754 239200 253810 240000
rect 255962 239200 256018 240000
rect 258262 239200 258318 240000
rect 260562 239200 260618 240000
rect 262862 239200 262918 240000
rect 265070 239200 265126 240000
rect 267370 239200 267426 240000
rect 269670 239200 269726 240000
rect 271970 239200 272026 240000
rect 274178 239200 274234 240000
rect 276478 239200 276534 240000
rect 278778 239200 278834 240000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8206 0 8262 800
rect 8758 0 8814 800
rect 9310 0 9366 800
rect 9862 0 9918 800
rect 10414 0 10470 800
rect 10966 0 11022 800
rect 11518 0 11574 800
rect 12162 0 12218 800
rect 12714 0 12770 800
rect 13266 0 13322 800
rect 13818 0 13874 800
rect 14370 0 14426 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17222 0 17278 800
rect 17774 0 17830 800
rect 18326 0 18382 800
rect 18878 0 18934 800
rect 19522 0 19578 800
rect 20074 0 20130 800
rect 20626 0 20682 800
rect 21178 0 21234 800
rect 21730 0 21786 800
rect 22282 0 22338 800
rect 22834 0 22890 800
rect 23478 0 23534 800
rect 24030 0 24086 800
rect 24582 0 24638 800
rect 25134 0 25190 800
rect 25686 0 25742 800
rect 26238 0 26294 800
rect 26790 0 26846 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29642 0 29698 800
rect 30194 0 30250 800
rect 30746 0 30802 800
rect 31390 0 31446 800
rect 31942 0 31998 800
rect 32494 0 32550 800
rect 33046 0 33102 800
rect 33598 0 33654 800
rect 34150 0 34206 800
rect 34702 0 34758 800
rect 35346 0 35402 800
rect 35898 0 35954 800
rect 36450 0 36506 800
rect 37002 0 37058 800
rect 37554 0 37610 800
rect 38106 0 38162 800
rect 38750 0 38806 800
rect 39302 0 39358 800
rect 39854 0 39910 800
rect 40406 0 40462 800
rect 40958 0 41014 800
rect 41510 0 41566 800
rect 42062 0 42118 800
rect 42706 0 42762 800
rect 43258 0 43314 800
rect 43810 0 43866 800
rect 44362 0 44418 800
rect 44914 0 44970 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46662 0 46718 800
rect 47214 0 47270 800
rect 47766 0 47822 800
rect 48318 0 48374 800
rect 48870 0 48926 800
rect 49422 0 49478 800
rect 49974 0 50030 800
rect 50618 0 50674 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 53378 0 53434 800
rect 54022 0 54078 800
rect 54574 0 54630 800
rect 55126 0 55182 800
rect 55678 0 55734 800
rect 56230 0 56286 800
rect 56782 0 56838 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58530 0 58586 800
rect 59082 0 59138 800
rect 59634 0 59690 800
rect 60186 0 60242 800
rect 60738 0 60794 800
rect 61290 0 61346 800
rect 61934 0 61990 800
rect 62486 0 62542 800
rect 63038 0 63094 800
rect 63590 0 63646 800
rect 64142 0 64198 800
rect 64694 0 64750 800
rect 65246 0 65302 800
rect 65890 0 65946 800
rect 66442 0 66498 800
rect 66994 0 67050 800
rect 67546 0 67602 800
rect 68098 0 68154 800
rect 68650 0 68706 800
rect 69202 0 69258 800
rect 69846 0 69902 800
rect 70398 0 70454 800
rect 70950 0 71006 800
rect 71502 0 71558 800
rect 72054 0 72110 800
rect 72606 0 72662 800
rect 73250 0 73306 800
rect 73802 0 73858 800
rect 74354 0 74410 800
rect 74906 0 74962 800
rect 75458 0 75514 800
rect 76010 0 76066 800
rect 76562 0 76618 800
rect 77206 0 77262 800
rect 77758 0 77814 800
rect 78310 0 78366 800
rect 78862 0 78918 800
rect 79414 0 79470 800
rect 79966 0 80022 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81714 0 81770 800
rect 82266 0 82322 800
rect 82818 0 82874 800
rect 83370 0 83426 800
rect 83922 0 83978 800
rect 84474 0 84530 800
rect 85118 0 85174 800
rect 85670 0 85726 800
rect 86222 0 86278 800
rect 86774 0 86830 800
rect 87326 0 87382 800
rect 87878 0 87934 800
rect 88522 0 88578 800
rect 89074 0 89130 800
rect 89626 0 89682 800
rect 90178 0 90234 800
rect 90730 0 90786 800
rect 91282 0 91338 800
rect 91834 0 91890 800
rect 92478 0 92534 800
rect 93030 0 93086 800
rect 93582 0 93638 800
rect 94134 0 94190 800
rect 94686 0 94742 800
rect 95238 0 95294 800
rect 95790 0 95846 800
rect 96434 0 96490 800
rect 96986 0 97042 800
rect 97538 0 97594 800
rect 98090 0 98146 800
rect 98642 0 98698 800
rect 99194 0 99250 800
rect 99746 0 99802 800
rect 100390 0 100446 800
rect 100942 0 100998 800
rect 101494 0 101550 800
rect 102046 0 102102 800
rect 102598 0 102654 800
rect 103150 0 103206 800
rect 103702 0 103758 800
rect 104346 0 104402 800
rect 104898 0 104954 800
rect 105450 0 105506 800
rect 106002 0 106058 800
rect 106554 0 106610 800
rect 107106 0 107162 800
rect 107750 0 107806 800
rect 108302 0 108358 800
rect 108854 0 108910 800
rect 109406 0 109462 800
rect 109958 0 110014 800
rect 110510 0 110566 800
rect 111062 0 111118 800
rect 111706 0 111762 800
rect 112258 0 112314 800
rect 112810 0 112866 800
rect 113362 0 113418 800
rect 113914 0 113970 800
rect 114466 0 114522 800
rect 115018 0 115074 800
rect 115662 0 115718 800
rect 116214 0 116270 800
rect 116766 0 116822 800
rect 117318 0 117374 800
rect 117870 0 117926 800
rect 118422 0 118478 800
rect 118974 0 119030 800
rect 119618 0 119674 800
rect 120170 0 120226 800
rect 120722 0 120778 800
rect 121274 0 121330 800
rect 121826 0 121882 800
rect 122378 0 122434 800
rect 123022 0 123078 800
rect 123574 0 123630 800
rect 124126 0 124182 800
rect 124678 0 124734 800
rect 125230 0 125286 800
rect 125782 0 125838 800
rect 126334 0 126390 800
rect 126978 0 127034 800
rect 127530 0 127586 800
rect 128082 0 128138 800
rect 128634 0 128690 800
rect 129186 0 129242 800
rect 129738 0 129794 800
rect 130290 0 130346 800
rect 130934 0 130990 800
rect 131486 0 131542 800
rect 132038 0 132094 800
rect 132590 0 132646 800
rect 133142 0 133198 800
rect 133694 0 133750 800
rect 134246 0 134302 800
rect 134890 0 134946 800
rect 135442 0 135498 800
rect 135994 0 136050 800
rect 136546 0 136602 800
rect 137098 0 137154 800
rect 137650 0 137706 800
rect 138202 0 138258 800
rect 138846 0 138902 800
rect 139398 0 139454 800
rect 139950 0 140006 800
rect 140502 0 140558 800
rect 141054 0 141110 800
rect 141606 0 141662 800
rect 142250 0 142306 800
rect 142802 0 142858 800
rect 143354 0 143410 800
rect 143906 0 143962 800
rect 144458 0 144514 800
rect 145010 0 145066 800
rect 145562 0 145618 800
rect 146206 0 146262 800
rect 146758 0 146814 800
rect 147310 0 147366 800
rect 147862 0 147918 800
rect 148414 0 148470 800
rect 148966 0 149022 800
rect 149518 0 149574 800
rect 150162 0 150218 800
rect 150714 0 150770 800
rect 151266 0 151322 800
rect 151818 0 151874 800
rect 152370 0 152426 800
rect 152922 0 152978 800
rect 153474 0 153530 800
rect 154118 0 154174 800
rect 154670 0 154726 800
rect 155222 0 155278 800
rect 155774 0 155830 800
rect 156326 0 156382 800
rect 156878 0 156934 800
rect 157430 0 157486 800
rect 158074 0 158130 800
rect 158626 0 158682 800
rect 159178 0 159234 800
rect 159730 0 159786 800
rect 160282 0 160338 800
rect 160834 0 160890 800
rect 161478 0 161534 800
rect 162030 0 162086 800
rect 162582 0 162638 800
rect 163134 0 163190 800
rect 163686 0 163742 800
rect 164238 0 164294 800
rect 164790 0 164846 800
rect 165434 0 165490 800
rect 165986 0 166042 800
rect 166538 0 166594 800
rect 167090 0 167146 800
rect 167642 0 167698 800
rect 168194 0 168250 800
rect 168746 0 168802 800
rect 169390 0 169446 800
rect 169942 0 169998 800
rect 170494 0 170550 800
rect 171046 0 171102 800
rect 171598 0 171654 800
rect 172150 0 172206 800
rect 172702 0 172758 800
rect 173346 0 173402 800
rect 173898 0 173954 800
rect 174450 0 174506 800
rect 175002 0 175058 800
rect 175554 0 175610 800
rect 176106 0 176162 800
rect 176750 0 176806 800
rect 177302 0 177358 800
rect 177854 0 177910 800
rect 178406 0 178462 800
rect 178958 0 179014 800
rect 179510 0 179566 800
rect 180062 0 180118 800
rect 180706 0 180762 800
rect 181258 0 181314 800
rect 181810 0 181866 800
rect 182362 0 182418 800
rect 182914 0 182970 800
rect 183466 0 183522 800
rect 184018 0 184074 800
rect 184662 0 184718 800
rect 185214 0 185270 800
rect 185766 0 185822 800
rect 186318 0 186374 800
rect 186870 0 186926 800
rect 187422 0 187478 800
rect 187974 0 188030 800
rect 188618 0 188674 800
rect 189170 0 189226 800
rect 189722 0 189778 800
rect 190274 0 190330 800
rect 190826 0 190882 800
rect 191378 0 191434 800
rect 191930 0 191986 800
rect 192574 0 192630 800
rect 193126 0 193182 800
rect 193678 0 193734 800
rect 194230 0 194286 800
rect 194782 0 194838 800
rect 195334 0 195390 800
rect 195978 0 196034 800
rect 196530 0 196586 800
rect 197082 0 197138 800
rect 197634 0 197690 800
rect 198186 0 198242 800
rect 198738 0 198794 800
rect 199290 0 199346 800
rect 199934 0 199990 800
rect 200486 0 200542 800
rect 201038 0 201094 800
rect 201590 0 201646 800
rect 202142 0 202198 800
rect 202694 0 202750 800
rect 203246 0 203302 800
rect 203890 0 203946 800
rect 204442 0 204498 800
rect 204994 0 205050 800
rect 205546 0 205602 800
rect 206098 0 206154 800
rect 206650 0 206706 800
rect 207202 0 207258 800
rect 207846 0 207902 800
rect 208398 0 208454 800
rect 208950 0 209006 800
rect 209502 0 209558 800
rect 210054 0 210110 800
rect 210606 0 210662 800
rect 211250 0 211306 800
rect 211802 0 211858 800
rect 212354 0 212410 800
rect 212906 0 212962 800
rect 213458 0 213514 800
rect 214010 0 214066 800
rect 214562 0 214618 800
rect 215206 0 215262 800
rect 215758 0 215814 800
rect 216310 0 216366 800
rect 216862 0 216918 800
rect 217414 0 217470 800
rect 217966 0 218022 800
rect 218518 0 218574 800
rect 219162 0 219218 800
rect 219714 0 219770 800
rect 220266 0 220322 800
rect 220818 0 220874 800
rect 221370 0 221426 800
rect 221922 0 221978 800
rect 222474 0 222530 800
rect 223118 0 223174 800
rect 223670 0 223726 800
rect 224222 0 224278 800
rect 224774 0 224830 800
rect 225326 0 225382 800
rect 225878 0 225934 800
rect 226430 0 226486 800
rect 227074 0 227130 800
rect 227626 0 227682 800
rect 228178 0 228234 800
rect 228730 0 228786 800
rect 229282 0 229338 800
rect 229834 0 229890 800
rect 230478 0 230534 800
rect 231030 0 231086 800
rect 231582 0 231638 800
rect 232134 0 232190 800
rect 232686 0 232742 800
rect 233238 0 233294 800
rect 233790 0 233846 800
rect 234434 0 234490 800
rect 234986 0 235042 800
rect 235538 0 235594 800
rect 236090 0 236146 800
rect 236642 0 236698 800
rect 237194 0 237250 800
rect 237746 0 237802 800
rect 238390 0 238446 800
rect 238942 0 238998 800
rect 239494 0 239550 800
rect 240046 0 240102 800
rect 240598 0 240654 800
rect 241150 0 241206 800
rect 241702 0 241758 800
rect 242346 0 242402 800
rect 242898 0 242954 800
rect 243450 0 243506 800
rect 244002 0 244058 800
rect 244554 0 244610 800
rect 245106 0 245162 800
rect 245750 0 245806 800
rect 246302 0 246358 800
rect 246854 0 246910 800
rect 247406 0 247462 800
rect 247958 0 248014 800
rect 248510 0 248566 800
rect 249062 0 249118 800
rect 249706 0 249762 800
rect 250258 0 250314 800
rect 250810 0 250866 800
rect 251362 0 251418 800
rect 251914 0 251970 800
rect 252466 0 252522 800
rect 253018 0 253074 800
rect 253662 0 253718 800
rect 254214 0 254270 800
rect 254766 0 254822 800
rect 255318 0 255374 800
rect 255870 0 255926 800
rect 256422 0 256478 800
rect 256974 0 257030 800
rect 257618 0 257674 800
rect 258170 0 258226 800
rect 258722 0 258778 800
rect 259274 0 259330 800
rect 259826 0 259882 800
rect 260378 0 260434 800
rect 260930 0 260986 800
rect 261574 0 261630 800
rect 262126 0 262182 800
rect 262678 0 262734 800
rect 263230 0 263286 800
rect 263782 0 263838 800
rect 264334 0 264390 800
rect 264978 0 265034 800
rect 265530 0 265586 800
rect 266082 0 266138 800
rect 266634 0 266690 800
rect 267186 0 267242 800
rect 267738 0 267794 800
rect 268290 0 268346 800
rect 268934 0 268990 800
rect 269486 0 269542 800
rect 270038 0 270094 800
rect 270590 0 270646 800
rect 271142 0 271198 800
rect 271694 0 271750 800
rect 272246 0 272302 800
rect 272890 0 272946 800
rect 273442 0 273498 800
rect 273994 0 274050 800
rect 274546 0 274602 800
rect 275098 0 275154 800
rect 275650 0 275706 800
rect 276202 0 276258 800
rect 276846 0 276902 800
rect 277398 0 277454 800
rect 277950 0 278006 800
rect 278502 0 278558 800
rect 279054 0 279110 800
rect 279606 0 279662 800
<< obsm2 >>
rect 296 239144 1066 239200
rect 1234 239144 3274 239200
rect 3442 239144 5574 239200
rect 5742 239144 7874 239200
rect 8042 239144 10082 239200
rect 10250 239144 12382 239200
rect 12550 239144 14682 239200
rect 14850 239144 16982 239200
rect 17150 239144 19190 239200
rect 19358 239144 21490 239200
rect 21658 239144 23790 239200
rect 23958 239144 26090 239200
rect 26258 239144 28298 239200
rect 28466 239144 30598 239200
rect 30766 239144 32898 239200
rect 33066 239144 35198 239200
rect 35366 239144 37406 239200
rect 37574 239144 39706 239200
rect 39874 239144 42006 239200
rect 42174 239144 44306 239200
rect 44474 239144 46514 239200
rect 46682 239144 48814 239200
rect 48982 239144 51114 239200
rect 51282 239144 53414 239200
rect 53582 239144 55622 239200
rect 55790 239144 57922 239200
rect 58090 239144 60222 239200
rect 60390 239144 62430 239200
rect 62598 239144 64730 239200
rect 64898 239144 67030 239200
rect 67198 239144 69330 239200
rect 69498 239144 71538 239200
rect 71706 239144 73838 239200
rect 74006 239144 76138 239200
rect 76306 239144 78438 239200
rect 78606 239144 80646 239200
rect 80814 239144 82946 239200
rect 83114 239144 85246 239200
rect 85414 239144 87546 239200
rect 87714 239144 89754 239200
rect 89922 239144 92054 239200
rect 92222 239144 94354 239200
rect 94522 239144 96654 239200
rect 96822 239144 98862 239200
rect 99030 239144 101162 239200
rect 101330 239144 103462 239200
rect 103630 239144 105762 239200
rect 105930 239144 107970 239200
rect 108138 239144 110270 239200
rect 110438 239144 112570 239200
rect 112738 239144 114778 239200
rect 114946 239144 117078 239200
rect 117246 239144 119378 239200
rect 119546 239144 121678 239200
rect 121846 239144 123886 239200
rect 124054 239144 126186 239200
rect 126354 239144 128486 239200
rect 128654 239144 130786 239200
rect 130954 239144 132994 239200
rect 133162 239144 135294 239200
rect 135462 239144 137594 239200
rect 137762 239144 139894 239200
rect 140062 239144 142102 239200
rect 142270 239144 144402 239200
rect 144570 239144 146702 239200
rect 146870 239144 149002 239200
rect 149170 239144 151210 239200
rect 151378 239144 153510 239200
rect 153678 239144 155810 239200
rect 155978 239144 158110 239200
rect 158278 239144 160318 239200
rect 160486 239144 162618 239200
rect 162786 239144 164918 239200
rect 165086 239144 167218 239200
rect 167386 239144 169426 239200
rect 169594 239144 171726 239200
rect 171894 239144 174026 239200
rect 174194 239144 176234 239200
rect 176402 239144 178534 239200
rect 178702 239144 180834 239200
rect 181002 239144 183134 239200
rect 183302 239144 185342 239200
rect 185510 239144 187642 239200
rect 187810 239144 189942 239200
rect 190110 239144 192242 239200
rect 192410 239144 194450 239200
rect 194618 239144 196750 239200
rect 196918 239144 199050 239200
rect 199218 239144 201350 239200
rect 201518 239144 203558 239200
rect 203726 239144 205858 239200
rect 206026 239144 208158 239200
rect 208326 239144 210458 239200
rect 210626 239144 212666 239200
rect 212834 239144 214966 239200
rect 215134 239144 217266 239200
rect 217434 239144 219566 239200
rect 219734 239144 221774 239200
rect 221942 239144 224074 239200
rect 224242 239144 226374 239200
rect 226542 239144 228582 239200
rect 228750 239144 230882 239200
rect 231050 239144 233182 239200
rect 233350 239144 235482 239200
rect 235650 239144 237690 239200
rect 237858 239144 239990 239200
rect 240158 239144 242290 239200
rect 242458 239144 244590 239200
rect 244758 239144 246798 239200
rect 246966 239144 249098 239200
rect 249266 239144 251398 239200
rect 251566 239144 253698 239200
rect 253866 239144 255906 239200
rect 256074 239144 258206 239200
rect 258374 239144 260506 239200
rect 260674 239144 262806 239200
rect 262974 239144 265014 239200
rect 265182 239144 267314 239200
rect 267482 239144 269614 239200
rect 269782 239144 271914 239200
rect 272082 239144 274122 239200
rect 274290 239144 276422 239200
rect 276590 239144 278722 239200
rect 278890 239144 279108 239200
rect 296 856 279108 239144
rect 406 800 790 856
rect 958 800 1342 856
rect 1510 800 1894 856
rect 2062 800 2446 856
rect 2614 800 2998 856
rect 3166 800 3550 856
rect 3718 800 4194 856
rect 4362 800 4746 856
rect 4914 800 5298 856
rect 5466 800 5850 856
rect 6018 800 6402 856
rect 6570 800 6954 856
rect 7122 800 7506 856
rect 7674 800 8150 856
rect 8318 800 8702 856
rect 8870 800 9254 856
rect 9422 800 9806 856
rect 9974 800 10358 856
rect 10526 800 10910 856
rect 11078 800 11462 856
rect 11630 800 12106 856
rect 12274 800 12658 856
rect 12826 800 13210 856
rect 13378 800 13762 856
rect 13930 800 14314 856
rect 14482 800 14866 856
rect 15034 800 15418 856
rect 15586 800 16062 856
rect 16230 800 16614 856
rect 16782 800 17166 856
rect 17334 800 17718 856
rect 17886 800 18270 856
rect 18438 800 18822 856
rect 18990 800 19466 856
rect 19634 800 20018 856
rect 20186 800 20570 856
rect 20738 800 21122 856
rect 21290 800 21674 856
rect 21842 800 22226 856
rect 22394 800 22778 856
rect 22946 800 23422 856
rect 23590 800 23974 856
rect 24142 800 24526 856
rect 24694 800 25078 856
rect 25246 800 25630 856
rect 25798 800 26182 856
rect 26350 800 26734 856
rect 26902 800 27378 856
rect 27546 800 27930 856
rect 28098 800 28482 856
rect 28650 800 29034 856
rect 29202 800 29586 856
rect 29754 800 30138 856
rect 30306 800 30690 856
rect 30858 800 31334 856
rect 31502 800 31886 856
rect 32054 800 32438 856
rect 32606 800 32990 856
rect 33158 800 33542 856
rect 33710 800 34094 856
rect 34262 800 34646 856
rect 34814 800 35290 856
rect 35458 800 35842 856
rect 36010 800 36394 856
rect 36562 800 36946 856
rect 37114 800 37498 856
rect 37666 800 38050 856
rect 38218 800 38694 856
rect 38862 800 39246 856
rect 39414 800 39798 856
rect 39966 800 40350 856
rect 40518 800 40902 856
rect 41070 800 41454 856
rect 41622 800 42006 856
rect 42174 800 42650 856
rect 42818 800 43202 856
rect 43370 800 43754 856
rect 43922 800 44306 856
rect 44474 800 44858 856
rect 45026 800 45410 856
rect 45578 800 45962 856
rect 46130 800 46606 856
rect 46774 800 47158 856
rect 47326 800 47710 856
rect 47878 800 48262 856
rect 48430 800 48814 856
rect 48982 800 49366 856
rect 49534 800 49918 856
rect 50086 800 50562 856
rect 50730 800 51114 856
rect 51282 800 51666 856
rect 51834 800 52218 856
rect 52386 800 52770 856
rect 52938 800 53322 856
rect 53490 800 53966 856
rect 54134 800 54518 856
rect 54686 800 55070 856
rect 55238 800 55622 856
rect 55790 800 56174 856
rect 56342 800 56726 856
rect 56894 800 57278 856
rect 57446 800 57922 856
rect 58090 800 58474 856
rect 58642 800 59026 856
rect 59194 800 59578 856
rect 59746 800 60130 856
rect 60298 800 60682 856
rect 60850 800 61234 856
rect 61402 800 61878 856
rect 62046 800 62430 856
rect 62598 800 62982 856
rect 63150 800 63534 856
rect 63702 800 64086 856
rect 64254 800 64638 856
rect 64806 800 65190 856
rect 65358 800 65834 856
rect 66002 800 66386 856
rect 66554 800 66938 856
rect 67106 800 67490 856
rect 67658 800 68042 856
rect 68210 800 68594 856
rect 68762 800 69146 856
rect 69314 800 69790 856
rect 69958 800 70342 856
rect 70510 800 70894 856
rect 71062 800 71446 856
rect 71614 800 71998 856
rect 72166 800 72550 856
rect 72718 800 73194 856
rect 73362 800 73746 856
rect 73914 800 74298 856
rect 74466 800 74850 856
rect 75018 800 75402 856
rect 75570 800 75954 856
rect 76122 800 76506 856
rect 76674 800 77150 856
rect 77318 800 77702 856
rect 77870 800 78254 856
rect 78422 800 78806 856
rect 78974 800 79358 856
rect 79526 800 79910 856
rect 80078 800 80462 856
rect 80630 800 81106 856
rect 81274 800 81658 856
rect 81826 800 82210 856
rect 82378 800 82762 856
rect 82930 800 83314 856
rect 83482 800 83866 856
rect 84034 800 84418 856
rect 84586 800 85062 856
rect 85230 800 85614 856
rect 85782 800 86166 856
rect 86334 800 86718 856
rect 86886 800 87270 856
rect 87438 800 87822 856
rect 87990 800 88466 856
rect 88634 800 89018 856
rect 89186 800 89570 856
rect 89738 800 90122 856
rect 90290 800 90674 856
rect 90842 800 91226 856
rect 91394 800 91778 856
rect 91946 800 92422 856
rect 92590 800 92974 856
rect 93142 800 93526 856
rect 93694 800 94078 856
rect 94246 800 94630 856
rect 94798 800 95182 856
rect 95350 800 95734 856
rect 95902 800 96378 856
rect 96546 800 96930 856
rect 97098 800 97482 856
rect 97650 800 98034 856
rect 98202 800 98586 856
rect 98754 800 99138 856
rect 99306 800 99690 856
rect 99858 800 100334 856
rect 100502 800 100886 856
rect 101054 800 101438 856
rect 101606 800 101990 856
rect 102158 800 102542 856
rect 102710 800 103094 856
rect 103262 800 103646 856
rect 103814 800 104290 856
rect 104458 800 104842 856
rect 105010 800 105394 856
rect 105562 800 105946 856
rect 106114 800 106498 856
rect 106666 800 107050 856
rect 107218 800 107694 856
rect 107862 800 108246 856
rect 108414 800 108798 856
rect 108966 800 109350 856
rect 109518 800 109902 856
rect 110070 800 110454 856
rect 110622 800 111006 856
rect 111174 800 111650 856
rect 111818 800 112202 856
rect 112370 800 112754 856
rect 112922 800 113306 856
rect 113474 800 113858 856
rect 114026 800 114410 856
rect 114578 800 114962 856
rect 115130 800 115606 856
rect 115774 800 116158 856
rect 116326 800 116710 856
rect 116878 800 117262 856
rect 117430 800 117814 856
rect 117982 800 118366 856
rect 118534 800 118918 856
rect 119086 800 119562 856
rect 119730 800 120114 856
rect 120282 800 120666 856
rect 120834 800 121218 856
rect 121386 800 121770 856
rect 121938 800 122322 856
rect 122490 800 122966 856
rect 123134 800 123518 856
rect 123686 800 124070 856
rect 124238 800 124622 856
rect 124790 800 125174 856
rect 125342 800 125726 856
rect 125894 800 126278 856
rect 126446 800 126922 856
rect 127090 800 127474 856
rect 127642 800 128026 856
rect 128194 800 128578 856
rect 128746 800 129130 856
rect 129298 800 129682 856
rect 129850 800 130234 856
rect 130402 800 130878 856
rect 131046 800 131430 856
rect 131598 800 131982 856
rect 132150 800 132534 856
rect 132702 800 133086 856
rect 133254 800 133638 856
rect 133806 800 134190 856
rect 134358 800 134834 856
rect 135002 800 135386 856
rect 135554 800 135938 856
rect 136106 800 136490 856
rect 136658 800 137042 856
rect 137210 800 137594 856
rect 137762 800 138146 856
rect 138314 800 138790 856
rect 138958 800 139342 856
rect 139510 800 139894 856
rect 140062 800 140446 856
rect 140614 800 140998 856
rect 141166 800 141550 856
rect 141718 800 142194 856
rect 142362 800 142746 856
rect 142914 800 143298 856
rect 143466 800 143850 856
rect 144018 800 144402 856
rect 144570 800 144954 856
rect 145122 800 145506 856
rect 145674 800 146150 856
rect 146318 800 146702 856
rect 146870 800 147254 856
rect 147422 800 147806 856
rect 147974 800 148358 856
rect 148526 800 148910 856
rect 149078 800 149462 856
rect 149630 800 150106 856
rect 150274 800 150658 856
rect 150826 800 151210 856
rect 151378 800 151762 856
rect 151930 800 152314 856
rect 152482 800 152866 856
rect 153034 800 153418 856
rect 153586 800 154062 856
rect 154230 800 154614 856
rect 154782 800 155166 856
rect 155334 800 155718 856
rect 155886 800 156270 856
rect 156438 800 156822 856
rect 156990 800 157374 856
rect 157542 800 158018 856
rect 158186 800 158570 856
rect 158738 800 159122 856
rect 159290 800 159674 856
rect 159842 800 160226 856
rect 160394 800 160778 856
rect 160946 800 161422 856
rect 161590 800 161974 856
rect 162142 800 162526 856
rect 162694 800 163078 856
rect 163246 800 163630 856
rect 163798 800 164182 856
rect 164350 800 164734 856
rect 164902 800 165378 856
rect 165546 800 165930 856
rect 166098 800 166482 856
rect 166650 800 167034 856
rect 167202 800 167586 856
rect 167754 800 168138 856
rect 168306 800 168690 856
rect 168858 800 169334 856
rect 169502 800 169886 856
rect 170054 800 170438 856
rect 170606 800 170990 856
rect 171158 800 171542 856
rect 171710 800 172094 856
rect 172262 800 172646 856
rect 172814 800 173290 856
rect 173458 800 173842 856
rect 174010 800 174394 856
rect 174562 800 174946 856
rect 175114 800 175498 856
rect 175666 800 176050 856
rect 176218 800 176694 856
rect 176862 800 177246 856
rect 177414 800 177798 856
rect 177966 800 178350 856
rect 178518 800 178902 856
rect 179070 800 179454 856
rect 179622 800 180006 856
rect 180174 800 180650 856
rect 180818 800 181202 856
rect 181370 800 181754 856
rect 181922 800 182306 856
rect 182474 800 182858 856
rect 183026 800 183410 856
rect 183578 800 183962 856
rect 184130 800 184606 856
rect 184774 800 185158 856
rect 185326 800 185710 856
rect 185878 800 186262 856
rect 186430 800 186814 856
rect 186982 800 187366 856
rect 187534 800 187918 856
rect 188086 800 188562 856
rect 188730 800 189114 856
rect 189282 800 189666 856
rect 189834 800 190218 856
rect 190386 800 190770 856
rect 190938 800 191322 856
rect 191490 800 191874 856
rect 192042 800 192518 856
rect 192686 800 193070 856
rect 193238 800 193622 856
rect 193790 800 194174 856
rect 194342 800 194726 856
rect 194894 800 195278 856
rect 195446 800 195922 856
rect 196090 800 196474 856
rect 196642 800 197026 856
rect 197194 800 197578 856
rect 197746 800 198130 856
rect 198298 800 198682 856
rect 198850 800 199234 856
rect 199402 800 199878 856
rect 200046 800 200430 856
rect 200598 800 200982 856
rect 201150 800 201534 856
rect 201702 800 202086 856
rect 202254 800 202638 856
rect 202806 800 203190 856
rect 203358 800 203834 856
rect 204002 800 204386 856
rect 204554 800 204938 856
rect 205106 800 205490 856
rect 205658 800 206042 856
rect 206210 800 206594 856
rect 206762 800 207146 856
rect 207314 800 207790 856
rect 207958 800 208342 856
rect 208510 800 208894 856
rect 209062 800 209446 856
rect 209614 800 209998 856
rect 210166 800 210550 856
rect 210718 800 211194 856
rect 211362 800 211746 856
rect 211914 800 212298 856
rect 212466 800 212850 856
rect 213018 800 213402 856
rect 213570 800 213954 856
rect 214122 800 214506 856
rect 214674 800 215150 856
rect 215318 800 215702 856
rect 215870 800 216254 856
rect 216422 800 216806 856
rect 216974 800 217358 856
rect 217526 800 217910 856
rect 218078 800 218462 856
rect 218630 800 219106 856
rect 219274 800 219658 856
rect 219826 800 220210 856
rect 220378 800 220762 856
rect 220930 800 221314 856
rect 221482 800 221866 856
rect 222034 800 222418 856
rect 222586 800 223062 856
rect 223230 800 223614 856
rect 223782 800 224166 856
rect 224334 800 224718 856
rect 224886 800 225270 856
rect 225438 800 225822 856
rect 225990 800 226374 856
rect 226542 800 227018 856
rect 227186 800 227570 856
rect 227738 800 228122 856
rect 228290 800 228674 856
rect 228842 800 229226 856
rect 229394 800 229778 856
rect 229946 800 230422 856
rect 230590 800 230974 856
rect 231142 800 231526 856
rect 231694 800 232078 856
rect 232246 800 232630 856
rect 232798 800 233182 856
rect 233350 800 233734 856
rect 233902 800 234378 856
rect 234546 800 234930 856
rect 235098 800 235482 856
rect 235650 800 236034 856
rect 236202 800 236586 856
rect 236754 800 237138 856
rect 237306 800 237690 856
rect 237858 800 238334 856
rect 238502 800 238886 856
rect 239054 800 239438 856
rect 239606 800 239990 856
rect 240158 800 240542 856
rect 240710 800 241094 856
rect 241262 800 241646 856
rect 241814 800 242290 856
rect 242458 800 242842 856
rect 243010 800 243394 856
rect 243562 800 243946 856
rect 244114 800 244498 856
rect 244666 800 245050 856
rect 245218 800 245694 856
rect 245862 800 246246 856
rect 246414 800 246798 856
rect 246966 800 247350 856
rect 247518 800 247902 856
rect 248070 800 248454 856
rect 248622 800 249006 856
rect 249174 800 249650 856
rect 249818 800 250202 856
rect 250370 800 250754 856
rect 250922 800 251306 856
rect 251474 800 251858 856
rect 252026 800 252410 856
rect 252578 800 252962 856
rect 253130 800 253606 856
rect 253774 800 254158 856
rect 254326 800 254710 856
rect 254878 800 255262 856
rect 255430 800 255814 856
rect 255982 800 256366 856
rect 256534 800 256918 856
rect 257086 800 257562 856
rect 257730 800 258114 856
rect 258282 800 258666 856
rect 258834 800 259218 856
rect 259386 800 259770 856
rect 259938 800 260322 856
rect 260490 800 260874 856
rect 261042 800 261518 856
rect 261686 800 262070 856
rect 262238 800 262622 856
rect 262790 800 263174 856
rect 263342 800 263726 856
rect 263894 800 264278 856
rect 264446 800 264922 856
rect 265090 800 265474 856
rect 265642 800 266026 856
rect 266194 800 266578 856
rect 266746 800 267130 856
rect 267298 800 267682 856
rect 267850 800 268234 856
rect 268402 800 268878 856
rect 269046 800 269430 856
rect 269598 800 269982 856
rect 270150 800 270534 856
rect 270702 800 271086 856
rect 271254 800 271638 856
rect 271806 800 272190 856
rect 272358 800 272834 856
rect 273002 800 273386 856
rect 273554 800 273938 856
rect 274106 800 274490 856
rect 274658 800 275042 856
rect 275210 800 275594 856
rect 275762 800 276146 856
rect 276314 800 276790 856
rect 276958 800 277342 856
rect 277510 800 277894 856
rect 278062 800 278446 856
rect 278614 800 278998 856
<< metal3 >>
rect 0 215976 800 216096
rect 0 167968 800 168088
rect 0 119960 800 120080
rect 0 71952 800 72072
rect 0 23944 800 24064
rect 279200 229848 280000 229968
rect 279200 209856 280000 209976
rect 279200 189864 280000 189984
rect 279200 169872 280000 169992
rect 279200 149880 280000 150000
rect 279200 129888 280000 130008
rect 279200 109896 280000 110016
rect 279200 89904 280000 90024
rect 279200 69912 280000 70032
rect 279200 49920 280000 50040
rect 279200 29928 280000 30048
rect 279200 9936 280000 10056
<< obsm3 >>
rect 4208 851 273871 237761
<< metal4 >>
rect 4208 2128 4528 237776
rect 19568 2128 19888 237776
rect 34928 2128 35248 237776
rect 50288 2128 50608 237776
rect 65648 2128 65968 237776
rect 81008 2128 81328 237776
rect 96368 2128 96688 237776
rect 111728 2128 112048 237776
rect 127088 2128 127408 237776
rect 142448 2128 142768 237776
rect 157808 2128 158128 237776
rect 173168 2128 173488 237776
rect 188528 2128 188848 237776
rect 203888 2128 204208 237776
rect 219248 2128 219568 237776
rect 234608 2128 234928 237776
rect 249968 2128 250288 237776
rect 265328 2128 265648 237776
<< obsm4 >>
rect 46979 5475 50208 235925
rect 50688 5475 65568 235925
rect 66048 5475 80928 235925
rect 81408 5475 96288 235925
rect 96768 5475 111648 235925
rect 112128 5475 127008 235925
rect 127488 5475 142368 235925
rect 142848 5475 144834 235925
<< obsm5 >>
rect 134436 96740 144876 100460
<< labels >>
rlabel metal2 s 260562 239200 260618 240000 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 267370 239200 267426 240000 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 0 167968 800 168088 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 279200 49920 280000 50040 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 278502 0 278558 800 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 279200 69912 280000 70032 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 279200 89904 280000 90024 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal3 s 279200 109896 280000 110016 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 279200 129888 280000 130008 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 279200 149880 280000 150000 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 279200 169872 280000 169992 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 0 23944 800 24064 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 269670 239200 269726 240000 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 215976 800 216096 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 279200 189864 280000 189984 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 271970 239200 272026 240000 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 274178 239200 274234 240000 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 279054 0 279110 800 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 276478 239200 276534 240000 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal2 s 278778 239200 278834 240000 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 279200 209856 280000 209976 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 279200 229848 280000 229968 6 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal2 s 262862 239200 262918 240000 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 279606 0 279662 800 6 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal3 s 0 71952 800 72072 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 279200 9936 280000 10056 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal2 s 277398 0 277454 800 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal2 s 265070 239200 265126 240000 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal3 s 0 119960 800 120080 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal3 s 279200 29928 280000 30048 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 277950 0 278006 800 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 1122 239200 1178 240000 6 io_in[0]
port 32 nsew signal input
rlabel metal2 s 69386 239200 69442 240000 6 io_in[10]
port 33 nsew signal input
rlabel metal2 s 76194 239200 76250 240000 6 io_in[11]
port 34 nsew signal input
rlabel metal2 s 83002 239200 83058 240000 6 io_in[12]
port 35 nsew signal input
rlabel metal2 s 89810 239200 89866 240000 6 io_in[13]
port 36 nsew signal input
rlabel metal2 s 96710 239200 96766 240000 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 103518 239200 103574 240000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 110326 239200 110382 240000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 117134 239200 117190 240000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 123942 239200 123998 240000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 130842 239200 130898 240000 6 io_in[19]
port 42 nsew signal input
rlabel metal2 s 7930 239200 7986 240000 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 137650 239200 137706 240000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 144458 239200 144514 240000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 151266 239200 151322 240000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 158166 239200 158222 240000 6 io_in[23]
port 47 nsew signal input
rlabel metal2 s 164974 239200 165030 240000 6 io_in[24]
port 48 nsew signal input
rlabel metal2 s 171782 239200 171838 240000 6 io_in[25]
port 49 nsew signal input
rlabel metal2 s 178590 239200 178646 240000 6 io_in[26]
port 50 nsew signal input
rlabel metal2 s 185398 239200 185454 240000 6 io_in[27]
port 51 nsew signal input
rlabel metal2 s 192298 239200 192354 240000 6 io_in[28]
port 52 nsew signal input
rlabel metal2 s 199106 239200 199162 240000 6 io_in[29]
port 53 nsew signal input
rlabel metal2 s 14738 239200 14794 240000 6 io_in[2]
port 54 nsew signal input
rlabel metal2 s 205914 239200 205970 240000 6 io_in[30]
port 55 nsew signal input
rlabel metal2 s 212722 239200 212778 240000 6 io_in[31]
port 56 nsew signal input
rlabel metal2 s 219622 239200 219678 240000 6 io_in[32]
port 57 nsew signal input
rlabel metal2 s 226430 239200 226486 240000 6 io_in[33]
port 58 nsew signal input
rlabel metal2 s 233238 239200 233294 240000 6 io_in[34]
port 59 nsew signal input
rlabel metal2 s 240046 239200 240102 240000 6 io_in[35]
port 60 nsew signal input
rlabel metal2 s 246854 239200 246910 240000 6 io_in[36]
port 61 nsew signal input
rlabel metal2 s 253754 239200 253810 240000 6 io_in[37]
port 62 nsew signal input
rlabel metal2 s 21546 239200 21602 240000 6 io_in[3]
port 63 nsew signal input
rlabel metal2 s 28354 239200 28410 240000 6 io_in[4]
port 64 nsew signal input
rlabel metal2 s 35254 239200 35310 240000 6 io_in[5]
port 65 nsew signal input
rlabel metal2 s 42062 239200 42118 240000 6 io_in[6]
port 66 nsew signal input
rlabel metal2 s 48870 239200 48926 240000 6 io_in[7]
port 67 nsew signal input
rlabel metal2 s 55678 239200 55734 240000 6 io_in[8]
port 68 nsew signal input
rlabel metal2 s 62486 239200 62542 240000 6 io_in[9]
port 69 nsew signal input
rlabel metal2 s 3330 239200 3386 240000 6 io_oeb[0]
port 70 nsew signal output
rlabel metal2 s 71594 239200 71650 240000 6 io_oeb[10]
port 71 nsew signal output
rlabel metal2 s 78494 239200 78550 240000 6 io_oeb[11]
port 72 nsew signal output
rlabel metal2 s 85302 239200 85358 240000 6 io_oeb[12]
port 73 nsew signal output
rlabel metal2 s 92110 239200 92166 240000 6 io_oeb[13]
port 74 nsew signal output
rlabel metal2 s 98918 239200 98974 240000 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 105818 239200 105874 240000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 112626 239200 112682 240000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 119434 239200 119490 240000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 126242 239200 126298 240000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 133050 239200 133106 240000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal2 s 10138 239200 10194 240000 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 139950 239200 140006 240000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 146758 239200 146814 240000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 153566 239200 153622 240000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 160374 239200 160430 240000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal2 s 167274 239200 167330 240000 6 io_oeb[24]
port 86 nsew signal output
rlabel metal2 s 174082 239200 174138 240000 6 io_oeb[25]
port 87 nsew signal output
rlabel metal2 s 180890 239200 180946 240000 6 io_oeb[26]
port 88 nsew signal output
rlabel metal2 s 187698 239200 187754 240000 6 io_oeb[27]
port 89 nsew signal output
rlabel metal2 s 194506 239200 194562 240000 6 io_oeb[28]
port 90 nsew signal output
rlabel metal2 s 201406 239200 201462 240000 6 io_oeb[29]
port 91 nsew signal output
rlabel metal2 s 17038 239200 17094 240000 6 io_oeb[2]
port 92 nsew signal output
rlabel metal2 s 208214 239200 208270 240000 6 io_oeb[30]
port 93 nsew signal output
rlabel metal2 s 215022 239200 215078 240000 6 io_oeb[31]
port 94 nsew signal output
rlabel metal2 s 221830 239200 221886 240000 6 io_oeb[32]
port 95 nsew signal output
rlabel metal2 s 228638 239200 228694 240000 6 io_oeb[33]
port 96 nsew signal output
rlabel metal2 s 235538 239200 235594 240000 6 io_oeb[34]
port 97 nsew signal output
rlabel metal2 s 242346 239200 242402 240000 6 io_oeb[35]
port 98 nsew signal output
rlabel metal2 s 249154 239200 249210 240000 6 io_oeb[36]
port 99 nsew signal output
rlabel metal2 s 255962 239200 256018 240000 6 io_oeb[37]
port 100 nsew signal output
rlabel metal2 s 23846 239200 23902 240000 6 io_oeb[3]
port 101 nsew signal output
rlabel metal2 s 30654 239200 30710 240000 6 io_oeb[4]
port 102 nsew signal output
rlabel metal2 s 37462 239200 37518 240000 6 io_oeb[5]
port 103 nsew signal output
rlabel metal2 s 44362 239200 44418 240000 6 io_oeb[6]
port 104 nsew signal output
rlabel metal2 s 51170 239200 51226 240000 6 io_oeb[7]
port 105 nsew signal output
rlabel metal2 s 57978 239200 58034 240000 6 io_oeb[8]
port 106 nsew signal output
rlabel metal2 s 64786 239200 64842 240000 6 io_oeb[9]
port 107 nsew signal output
rlabel metal2 s 5630 239200 5686 240000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 73894 239200 73950 240000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 80702 239200 80758 240000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 87602 239200 87658 240000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 94410 239200 94466 240000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 101218 239200 101274 240000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 108026 239200 108082 240000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 114834 239200 114890 240000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 121734 239200 121790 240000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 128542 239200 128598 240000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 135350 239200 135406 240000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 12438 239200 12494 240000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 142158 239200 142214 240000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 149058 239200 149114 240000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 155866 239200 155922 240000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 162674 239200 162730 240000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 169482 239200 169538 240000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 176290 239200 176346 240000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 183190 239200 183246 240000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 189998 239200 190054 240000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 196806 239200 196862 240000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 203614 239200 203670 240000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 19246 239200 19302 240000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 210514 239200 210570 240000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 217322 239200 217378 240000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 224130 239200 224186 240000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 230938 239200 230994 240000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 237746 239200 237802 240000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 244646 239200 244702 240000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 251454 239200 251510 240000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 258262 239200 258318 240000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 26146 239200 26202 240000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 32954 239200 33010 240000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 39762 239200 39818 240000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 46570 239200 46626 240000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 53470 239200 53526 240000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 60278 239200 60334 240000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 67086 239200 67142 240000 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 229834 0 229890 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 234986 0 235042 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 238390 0 238446 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 240046 0 240102 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 243450 0 243506 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 245106 0 245162 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 246854 0 246910 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 248510 0 248566 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 250258 0 250314 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 251914 0 251970 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 253662 0 253718 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 255318 0 255374 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 256974 0 257030 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 258722 0 258778 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 260378 0 260434 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 262126 0 262182 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 263782 0 263838 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 265530 0 265586 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 267186 0 267242 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 268934 0 268990 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 270590 0 270646 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 272246 0 272302 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 273994 0 274050 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 275650 0 275706 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 170494 0 170550 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 178958 0 179014 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 180706 0 180762 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 182362 0 182418 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 184018 0 184074 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 185766 0 185822 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 189170 0 189226 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 194230 0 194286 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 202694 0 202750 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 204442 0 204498 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 207846 0 207902 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 209502 0 209558 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 211250 0 211306 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 214562 0 214618 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 216310 0 216366 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 217966 0 218022 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 219714 0 219770 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 221370 0 221426 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 226430 0 226486 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 228178 0 228234 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 230478 0 230534 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 232134 0 232190 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 233790 0 233846 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 235538 0 235594 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 237194 0 237250 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 238942 0 238998 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 240598 0 240654 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 242346 0 242402 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 244002 0 244058 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 245750 0 245806 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 247406 0 247462 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 249062 0 249118 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 250810 0 250866 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 252466 0 252522 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 254214 0 254270 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 255870 0 255926 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 257618 0 257674 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 259274 0 259330 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 260930 0 260986 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 262678 0 262734 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 264334 0 264390 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 266082 0 266138 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 267738 0 267794 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 269486 0 269542 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 271142 0 271198 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 272890 0 272946 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 274546 0 274602 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 276202 0 276258 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 99746 0 99802 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 126978 0 127034 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 142250 0 142306 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 143906 0 143962 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 147310 0 147366 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 148966 0 149022 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 152370 0 152426 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 154118 0 154174 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 155774 0 155830 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 160834 0 160890 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 162582 0 162638 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 165986 0 166042 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 171046 0 171102 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 174450 0 174506 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 176106 0 176162 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 177854 0 177910 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 179510 0 179566 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 182914 0 182970 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 184662 0 184718 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 186318 0 186374 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 187974 0 188030 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 189722 0 189778 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 191378 0 191434 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 193126 0 193182 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 194782 0 194838 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 196530 0 196586 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 198186 0 198242 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 199934 0 199990 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 201590 0 201646 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 203246 0 203302 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 204994 0 205050 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 206650 0 206706 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 208398 0 208454 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 210054 0 210110 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 211802 0 211858 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 213458 0 213514 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 215206 0 215262 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 216862 0 216918 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 218518 0 218574 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 220266 0 220322 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 221922 0 221978 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 223670 0 223726 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 225326 0 225382 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 227074 0 227130 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 228730 0 228786 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 231030 0 231086 800 6 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 232686 0 232742 800 6 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 234434 0 234490 800 6 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 236090 0 236146 800 6 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 237746 0 237802 800 6 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 239494 0 239550 800 6 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 241150 0 241206 800 6 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 242898 0 242954 800 6 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 244554 0 244610 800 6 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 246302 0 246358 800 6 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 247958 0 248014 800 6 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 249706 0 249762 800 6 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 251362 0 251418 800 6 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 253018 0 253074 800 6 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 254766 0 254822 800 6 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 256422 0 256478 800 6 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 258170 0 258226 800 6 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 259826 0 259882 800 6 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 261574 0 261630 800 6 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 263230 0 263286 800 6 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 264978 0 265034 800 6 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 266634 0 266690 800 6 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 268290 0 268346 800 6 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 270038 0 270094 800 6 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 271694 0 271750 800 6 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 273442 0 273498 800 6 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 275098 0 275154 800 6 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 276846 0 276902 800 6 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 181810 0 181866 800 6 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 186870 0 186926 800 6 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 193678 0 193734 800 6 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 195334 0 195390 800 6 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 197082 0 197138 800 6 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 198738 0 198794 800 6 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 200486 0 200542 800 6 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 202142 0 202198 800 6 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 203890 0 203946 800 6 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 205546 0 205602 800 6 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 208950 0 209006 800 6 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 210606 0 210662 800 6 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 212354 0 212410 800 6 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 214010 0 214066 800 6 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 217414 0 217470 800 6 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 219162 0 219218 800 6 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 220818 0 220874 800 6 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 224222 0 224278 800 6 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 225878 0 225934 800 6 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 227626 0 227682 800 6 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 530 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 531 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 532 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 wbs_adr_i[0]
port 533 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_adr_i[10]
port 534 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[11]
port 535 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[12]
port 536 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[13]
port 537 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[14]
port 538 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[15]
port 539 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_adr_i[16]
port 540 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_adr_i[17]
port 541 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_adr_i[18]
port 542 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_adr_i[19]
port 543 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[1]
port 544 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_adr_i[20]
port 545 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wbs_adr_i[21]
port 546 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_adr_i[22]
port 547 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_adr_i[23]
port 548 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 wbs_adr_i[24]
port 549 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_adr_i[25]
port 550 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wbs_adr_i[26]
port 551 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 wbs_adr_i[27]
port 552 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_adr_i[28]
port 553 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_adr_i[29]
port 554 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[2]
port 555 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 wbs_adr_i[30]
port 556 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_adr_i[31]
port 557 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[3]
port 558 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[4]
port 559 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_adr_i[5]
port 560 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[6]
port 561 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[7]
port 562 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_adr_i[8]
port 563 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[9]
port 564 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_cyc_i
port 565 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_i[0]
port 566 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_i[10]
port 567 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_i[11]
port 568 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_i[12]
port 569 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[13]
port 570 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[14]
port 571 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_i[15]
port 572 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_i[16]
port 573 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_i[17]
port 574 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_i[18]
port 575 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_i[19]
port 576 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[1]
port 577 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_i[20]
port 578 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_dat_i[21]
port 579 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_dat_i[22]
port 580 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_i[23]
port 581 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 wbs_dat_i[24]
port 582 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 wbs_dat_i[25]
port 583 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_i[26]
port 584 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 wbs_dat_i[27]
port 585 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_i[28]
port 586 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_dat_i[29]
port 587 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[2]
port 588 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_dat_i[30]
port 589 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 wbs_dat_i[31]
port 590 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[3]
port 591 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[4]
port 592 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[5]
port 593 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[6]
port 594 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_i[7]
port 595 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_i[8]
port 596 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[9]
port 597 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_o[0]
port 598 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[10]
port 599 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_o[11]
port 600 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_o[12]
port 601 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[13]
port 602 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[14]
port 603 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_o[15]
port 604 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_o[16]
port 605 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_o[17]
port 606 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_o[18]
port 607 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[19]
port 608 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_o[1]
port 609 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_o[20]
port 610 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_o[21]
port 611 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 wbs_dat_o[22]
port 612 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[23]
port 613 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 wbs_dat_o[24]
port 614 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_o[25]
port 615 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_o[26]
port 616 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_o[27]
port 617 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 wbs_dat_o[28]
port 618 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 wbs_dat_o[29]
port 619 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_o[2]
port 620 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 wbs_dat_o[30]
port 621 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 wbs_dat_o[31]
port 622 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_o[3]
port 623 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_o[4]
port 624 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[5]
port 625 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[6]
port 626 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[7]
port 627 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[8]
port 628 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[9]
port 629 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 wbs_sel_i[0]
port 630 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_sel_i[1]
port 631 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_sel_i[2]
port 632 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_sel_i[3]
port 633 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_stb_i
port 634 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_we_i
port 635 nsew signal input
rlabel metal4 s 249968 2128 250288 237776 6 VPWR
port 636 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 237776 6 VPWR
port 637 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 237776 6 VPWR
port 638 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 237776 6 VPWR
port 639 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 237776 6 VPWR
port 640 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 237776 6 VPWR
port 641 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 237776 6 VPWR
port 642 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 237776 6 VPWR
port 643 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 237776 6 VPWR
port 644 nsew power bidirectional
rlabel metal4 s 265328 2128 265648 237776 6 VGND
port 645 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 237776 6 VGND
port 646 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 237776 6 VGND
port 647 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 237776 6 VGND
port 648 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 237776 6 VGND
port 649 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 237776 6 VGND
port 650 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 237776 6 VGND
port 651 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 237776 6 VGND
port 652 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 237776 6 VGND
port 653 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 280000 240000
string LEFview TRUE
<< end >>
