magic
tech sky130A
magscale 1 2
timestamp 1611887857
<< obsli1 >>
rect 1104 2159 278852 237745
<< obsm1 >>
rect 290 2048 278852 237776
<< metal2 >>
rect 1122 239200 1178 240000
rect 3422 239200 3478 240000
rect 5814 239200 5870 240000
rect 8114 239200 8170 240000
rect 10506 239200 10562 240000
rect 12806 239200 12862 240000
rect 15198 239200 15254 240000
rect 17590 239200 17646 240000
rect 19890 239200 19946 240000
rect 22282 239200 22338 240000
rect 24582 239200 24638 240000
rect 26974 239200 27030 240000
rect 29274 239200 29330 240000
rect 31666 239200 31722 240000
rect 34058 239200 34114 240000
rect 36358 239200 36414 240000
rect 38750 239200 38806 240000
rect 41050 239200 41106 240000
rect 43442 239200 43498 240000
rect 45742 239200 45798 240000
rect 48134 239200 48190 240000
rect 50526 239200 50582 240000
rect 52826 239200 52882 240000
rect 55218 239200 55274 240000
rect 57518 239200 57574 240000
rect 59910 239200 59966 240000
rect 62210 239200 62266 240000
rect 64602 239200 64658 240000
rect 66994 239200 67050 240000
rect 69294 239200 69350 240000
rect 71686 239200 71742 240000
rect 73986 239200 74042 240000
rect 76378 239200 76434 240000
rect 78678 239200 78734 240000
rect 81070 239200 81126 240000
rect 83462 239200 83518 240000
rect 85762 239200 85818 240000
rect 88154 239200 88210 240000
rect 90454 239200 90510 240000
rect 92846 239200 92902 240000
rect 95146 239200 95202 240000
rect 97538 239200 97594 240000
rect 99930 239200 99986 240000
rect 102230 239200 102286 240000
rect 104622 239200 104678 240000
rect 106922 239200 106978 240000
rect 109314 239200 109370 240000
rect 111614 239200 111670 240000
rect 114006 239200 114062 240000
rect 116398 239200 116454 240000
rect 118698 239200 118754 240000
rect 121090 239200 121146 240000
rect 123390 239200 123446 240000
rect 125782 239200 125838 240000
rect 128082 239200 128138 240000
rect 130474 239200 130530 240000
rect 132866 239200 132922 240000
rect 135166 239200 135222 240000
rect 137558 239200 137614 240000
rect 139858 239200 139914 240000
rect 142250 239200 142306 240000
rect 144550 239200 144606 240000
rect 146942 239200 146998 240000
rect 149334 239200 149390 240000
rect 151634 239200 151690 240000
rect 154026 239200 154082 240000
rect 156326 239200 156382 240000
rect 158718 239200 158774 240000
rect 161018 239200 161074 240000
rect 163410 239200 163466 240000
rect 165802 239200 165858 240000
rect 168102 239200 168158 240000
rect 170494 239200 170550 240000
rect 172794 239200 172850 240000
rect 175186 239200 175242 240000
rect 177486 239200 177542 240000
rect 179878 239200 179934 240000
rect 182270 239200 182326 240000
rect 184570 239200 184626 240000
rect 186962 239200 187018 240000
rect 189262 239200 189318 240000
rect 191654 239200 191710 240000
rect 193954 239200 194010 240000
rect 196346 239200 196402 240000
rect 198738 239200 198794 240000
rect 201038 239200 201094 240000
rect 203430 239200 203486 240000
rect 205730 239200 205786 240000
rect 208122 239200 208178 240000
rect 210422 239200 210478 240000
rect 212814 239200 212870 240000
rect 215206 239200 215262 240000
rect 217506 239200 217562 240000
rect 219898 239200 219954 240000
rect 222198 239200 222254 240000
rect 224590 239200 224646 240000
rect 226890 239200 226946 240000
rect 229282 239200 229338 240000
rect 231674 239200 231730 240000
rect 233974 239200 234030 240000
rect 236366 239200 236422 240000
rect 238666 239200 238722 240000
rect 241058 239200 241114 240000
rect 243358 239200 243414 240000
rect 245750 239200 245806 240000
rect 248142 239200 248198 240000
rect 250442 239200 250498 240000
rect 252834 239200 252890 240000
rect 255134 239200 255190 240000
rect 257526 239200 257582 240000
rect 259826 239200 259882 240000
rect 262218 239200 262274 240000
rect 264610 239200 264666 240000
rect 266910 239200 266966 240000
rect 269302 239200 269358 240000
rect 271602 239200 271658 240000
rect 273994 239200 274050 240000
rect 276294 239200 276350 240000
rect 278686 239200 278742 240000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6366 0 6422 800
rect 6918 0 6974 800
rect 7470 0 7526 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 11978 0 12034 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17590 0 17646 800
rect 18142 0 18198 800
rect 18694 0 18750 800
rect 19246 0 19302 800
rect 19798 0 19854 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21454 0 21510 800
rect 22006 0 22062 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23754 0 23810 800
rect 24306 0 24362 800
rect 24858 0 24914 800
rect 25410 0 25466 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 27066 0 27122 800
rect 27618 0 27674 800
rect 28170 0 28226 800
rect 28722 0 28778 800
rect 29274 0 29330 800
rect 29826 0 29882 800
rect 30378 0 30434 800
rect 31022 0 31078 800
rect 31574 0 31630 800
rect 32126 0 32182 800
rect 32678 0 32734 800
rect 33230 0 33286 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 35438 0 35494 800
rect 35990 0 36046 800
rect 36542 0 36598 800
rect 37094 0 37150 800
rect 37646 0 37702 800
rect 38290 0 38346 800
rect 38842 0 38898 800
rect 39394 0 39450 800
rect 39946 0 40002 800
rect 40498 0 40554 800
rect 41050 0 41106 800
rect 41602 0 41658 800
rect 42154 0 42210 800
rect 42706 0 42762 800
rect 43258 0 43314 800
rect 43810 0 43866 800
rect 44362 0 44418 800
rect 44914 0 44970 800
rect 45466 0 45522 800
rect 46110 0 46166 800
rect 46662 0 46718 800
rect 47214 0 47270 800
rect 47766 0 47822 800
rect 48318 0 48374 800
rect 48870 0 48926 800
rect 49422 0 49478 800
rect 49974 0 50030 800
rect 50526 0 50582 800
rect 51078 0 51134 800
rect 51630 0 51686 800
rect 52182 0 52238 800
rect 52734 0 52790 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54482 0 54538 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58898 0 58954 800
rect 59450 0 59506 800
rect 60002 0 60058 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62854 0 62910 800
rect 63406 0 63462 800
rect 63958 0 64014 800
rect 64510 0 64566 800
rect 65062 0 65118 800
rect 65614 0 65670 800
rect 66166 0 66222 800
rect 66718 0 66774 800
rect 67270 0 67326 800
rect 67822 0 67878 800
rect 68466 0 68522 800
rect 69018 0 69074 800
rect 69570 0 69626 800
rect 70122 0 70178 800
rect 70674 0 70730 800
rect 71226 0 71282 800
rect 71778 0 71834 800
rect 72330 0 72386 800
rect 72882 0 72938 800
rect 73434 0 73490 800
rect 73986 0 74042 800
rect 74538 0 74594 800
rect 75090 0 75146 800
rect 75642 0 75698 800
rect 76286 0 76342 800
rect 76838 0 76894 800
rect 77390 0 77446 800
rect 77942 0 77998 800
rect 78494 0 78550 800
rect 79046 0 79102 800
rect 79598 0 79654 800
rect 80150 0 80206 800
rect 80702 0 80758 800
rect 81254 0 81310 800
rect 81806 0 81862 800
rect 82358 0 82414 800
rect 82910 0 82966 800
rect 83554 0 83610 800
rect 84106 0 84162 800
rect 84658 0 84714 800
rect 85210 0 85266 800
rect 85762 0 85818 800
rect 86314 0 86370 800
rect 86866 0 86922 800
rect 87418 0 87474 800
rect 87970 0 88026 800
rect 88522 0 88578 800
rect 89074 0 89130 800
rect 89626 0 89682 800
rect 90178 0 90234 800
rect 90730 0 90786 800
rect 91374 0 91430 800
rect 91926 0 91982 800
rect 92478 0 92534 800
rect 93030 0 93086 800
rect 93582 0 93638 800
rect 94134 0 94190 800
rect 94686 0 94742 800
rect 95238 0 95294 800
rect 95790 0 95846 800
rect 96342 0 96398 800
rect 96894 0 96950 800
rect 97446 0 97502 800
rect 97998 0 98054 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99746 0 99802 800
rect 100298 0 100354 800
rect 100850 0 100906 800
rect 101402 0 101458 800
rect 101954 0 102010 800
rect 102506 0 102562 800
rect 103058 0 103114 800
rect 103610 0 103666 800
rect 104162 0 104218 800
rect 104714 0 104770 800
rect 105266 0 105322 800
rect 105818 0 105874 800
rect 106462 0 106518 800
rect 107014 0 107070 800
rect 107566 0 107622 800
rect 108118 0 108174 800
rect 108670 0 108726 800
rect 109222 0 109278 800
rect 109774 0 109830 800
rect 110326 0 110382 800
rect 110878 0 110934 800
rect 111430 0 111486 800
rect 111982 0 112038 800
rect 112534 0 112590 800
rect 113086 0 113142 800
rect 113638 0 113694 800
rect 114282 0 114338 800
rect 114834 0 114890 800
rect 115386 0 115442 800
rect 115938 0 115994 800
rect 116490 0 116546 800
rect 117042 0 117098 800
rect 117594 0 117650 800
rect 118146 0 118202 800
rect 118698 0 118754 800
rect 119250 0 119306 800
rect 119802 0 119858 800
rect 120354 0 120410 800
rect 120906 0 120962 800
rect 121550 0 121606 800
rect 122102 0 122158 800
rect 122654 0 122710 800
rect 123206 0 123262 800
rect 123758 0 123814 800
rect 124310 0 124366 800
rect 124862 0 124918 800
rect 125414 0 125470 800
rect 125966 0 126022 800
rect 126518 0 126574 800
rect 127070 0 127126 800
rect 127622 0 127678 800
rect 128174 0 128230 800
rect 128726 0 128782 800
rect 129370 0 129426 800
rect 129922 0 129978 800
rect 130474 0 130530 800
rect 131026 0 131082 800
rect 131578 0 131634 800
rect 132130 0 132186 800
rect 132682 0 132738 800
rect 133234 0 133290 800
rect 133786 0 133842 800
rect 134338 0 134394 800
rect 134890 0 134946 800
rect 135442 0 135498 800
rect 135994 0 136050 800
rect 136638 0 136694 800
rect 137190 0 137246 800
rect 137742 0 137798 800
rect 138294 0 138350 800
rect 138846 0 138902 800
rect 139398 0 139454 800
rect 139950 0 140006 800
rect 140502 0 140558 800
rect 141054 0 141110 800
rect 141606 0 141662 800
rect 142158 0 142214 800
rect 142710 0 142766 800
rect 143262 0 143318 800
rect 143814 0 143870 800
rect 144458 0 144514 800
rect 145010 0 145066 800
rect 145562 0 145618 800
rect 146114 0 146170 800
rect 146666 0 146722 800
rect 147218 0 147274 800
rect 147770 0 147826 800
rect 148322 0 148378 800
rect 148874 0 148930 800
rect 149426 0 149482 800
rect 149978 0 150034 800
rect 150530 0 150586 800
rect 151082 0 151138 800
rect 151726 0 151782 800
rect 152278 0 152334 800
rect 152830 0 152886 800
rect 153382 0 153438 800
rect 153934 0 153990 800
rect 154486 0 154542 800
rect 155038 0 155094 800
rect 155590 0 155646 800
rect 156142 0 156198 800
rect 156694 0 156750 800
rect 157246 0 157302 800
rect 157798 0 157854 800
rect 158350 0 158406 800
rect 158902 0 158958 800
rect 159546 0 159602 800
rect 160098 0 160154 800
rect 160650 0 160706 800
rect 161202 0 161258 800
rect 161754 0 161810 800
rect 162306 0 162362 800
rect 162858 0 162914 800
rect 163410 0 163466 800
rect 163962 0 164018 800
rect 164514 0 164570 800
rect 165066 0 165122 800
rect 165618 0 165674 800
rect 166170 0 166226 800
rect 166814 0 166870 800
rect 167366 0 167422 800
rect 167918 0 167974 800
rect 168470 0 168526 800
rect 169022 0 169078 800
rect 169574 0 169630 800
rect 170126 0 170182 800
rect 170678 0 170734 800
rect 171230 0 171286 800
rect 171782 0 171838 800
rect 172334 0 172390 800
rect 172886 0 172942 800
rect 173438 0 173494 800
rect 173990 0 174046 800
rect 174634 0 174690 800
rect 175186 0 175242 800
rect 175738 0 175794 800
rect 176290 0 176346 800
rect 176842 0 176898 800
rect 177394 0 177450 800
rect 177946 0 178002 800
rect 178498 0 178554 800
rect 179050 0 179106 800
rect 179602 0 179658 800
rect 180154 0 180210 800
rect 180706 0 180762 800
rect 181258 0 181314 800
rect 181902 0 181958 800
rect 182454 0 182510 800
rect 183006 0 183062 800
rect 183558 0 183614 800
rect 184110 0 184166 800
rect 184662 0 184718 800
rect 185214 0 185270 800
rect 185766 0 185822 800
rect 186318 0 186374 800
rect 186870 0 186926 800
rect 187422 0 187478 800
rect 187974 0 188030 800
rect 188526 0 188582 800
rect 189078 0 189134 800
rect 189722 0 189778 800
rect 190274 0 190330 800
rect 190826 0 190882 800
rect 191378 0 191434 800
rect 191930 0 191986 800
rect 192482 0 192538 800
rect 193034 0 193090 800
rect 193586 0 193642 800
rect 194138 0 194194 800
rect 194690 0 194746 800
rect 195242 0 195298 800
rect 195794 0 195850 800
rect 196346 0 196402 800
rect 196898 0 196954 800
rect 197542 0 197598 800
rect 198094 0 198150 800
rect 198646 0 198702 800
rect 199198 0 199254 800
rect 199750 0 199806 800
rect 200302 0 200358 800
rect 200854 0 200910 800
rect 201406 0 201462 800
rect 201958 0 202014 800
rect 202510 0 202566 800
rect 203062 0 203118 800
rect 203614 0 203670 800
rect 204166 0 204222 800
rect 204810 0 204866 800
rect 205362 0 205418 800
rect 205914 0 205970 800
rect 206466 0 206522 800
rect 207018 0 207074 800
rect 207570 0 207626 800
rect 208122 0 208178 800
rect 208674 0 208730 800
rect 209226 0 209282 800
rect 209778 0 209834 800
rect 210330 0 210386 800
rect 210882 0 210938 800
rect 211434 0 211490 800
rect 211986 0 212042 800
rect 212630 0 212686 800
rect 213182 0 213238 800
rect 213734 0 213790 800
rect 214286 0 214342 800
rect 214838 0 214894 800
rect 215390 0 215446 800
rect 215942 0 215998 800
rect 216494 0 216550 800
rect 217046 0 217102 800
rect 217598 0 217654 800
rect 218150 0 218206 800
rect 218702 0 218758 800
rect 219254 0 219310 800
rect 219898 0 219954 800
rect 220450 0 220506 800
rect 221002 0 221058 800
rect 221554 0 221610 800
rect 222106 0 222162 800
rect 222658 0 222714 800
rect 223210 0 223266 800
rect 223762 0 223818 800
rect 224314 0 224370 800
rect 224866 0 224922 800
rect 225418 0 225474 800
rect 225970 0 226026 800
rect 226522 0 226578 800
rect 227074 0 227130 800
rect 227718 0 227774 800
rect 228270 0 228326 800
rect 228822 0 228878 800
rect 229374 0 229430 800
rect 229926 0 229982 800
rect 230478 0 230534 800
rect 231030 0 231086 800
rect 231582 0 231638 800
rect 232134 0 232190 800
rect 232686 0 232742 800
rect 233238 0 233294 800
rect 233790 0 233846 800
rect 234342 0 234398 800
rect 234986 0 235042 800
rect 235538 0 235594 800
rect 236090 0 236146 800
rect 236642 0 236698 800
rect 237194 0 237250 800
rect 237746 0 237802 800
rect 238298 0 238354 800
rect 238850 0 238906 800
rect 239402 0 239458 800
rect 239954 0 240010 800
rect 240506 0 240562 800
rect 241058 0 241114 800
rect 241610 0 241666 800
rect 242162 0 242218 800
rect 242806 0 242862 800
rect 243358 0 243414 800
rect 243910 0 243966 800
rect 244462 0 244518 800
rect 245014 0 245070 800
rect 245566 0 245622 800
rect 246118 0 246174 800
rect 246670 0 246726 800
rect 247222 0 247278 800
rect 247774 0 247830 800
rect 248326 0 248382 800
rect 248878 0 248934 800
rect 249430 0 249486 800
rect 250074 0 250130 800
rect 250626 0 250682 800
rect 251178 0 251234 800
rect 251730 0 251786 800
rect 252282 0 252338 800
rect 252834 0 252890 800
rect 253386 0 253442 800
rect 253938 0 253994 800
rect 254490 0 254546 800
rect 255042 0 255098 800
rect 255594 0 255650 800
rect 256146 0 256202 800
rect 256698 0 256754 800
rect 257250 0 257306 800
rect 257894 0 257950 800
rect 258446 0 258502 800
rect 258998 0 259054 800
rect 259550 0 259606 800
rect 260102 0 260158 800
rect 260654 0 260710 800
rect 261206 0 261262 800
rect 261758 0 261814 800
rect 262310 0 262366 800
rect 262862 0 262918 800
rect 263414 0 263470 800
rect 263966 0 264022 800
rect 264518 0 264574 800
rect 265162 0 265218 800
rect 265714 0 265770 800
rect 266266 0 266322 800
rect 266818 0 266874 800
rect 267370 0 267426 800
rect 267922 0 267978 800
rect 268474 0 268530 800
rect 269026 0 269082 800
rect 269578 0 269634 800
rect 270130 0 270186 800
rect 270682 0 270738 800
rect 271234 0 271290 800
rect 271786 0 271842 800
rect 272338 0 272394 800
rect 272982 0 273038 800
rect 273534 0 273590 800
rect 274086 0 274142 800
rect 274638 0 274694 800
rect 275190 0 275246 800
rect 275742 0 275798 800
rect 276294 0 276350 800
rect 276846 0 276902 800
rect 277398 0 277454 800
rect 277950 0 278006 800
rect 278502 0 278558 800
rect 279054 0 279110 800
rect 279606 0 279662 800
<< obsm2 >>
rect 296 239144 1066 239200
rect 1234 239144 3366 239200
rect 3534 239144 5758 239200
rect 5926 239144 8058 239200
rect 8226 239144 10450 239200
rect 10618 239144 12750 239200
rect 12918 239144 15142 239200
rect 15310 239144 17534 239200
rect 17702 239144 19834 239200
rect 20002 239144 22226 239200
rect 22394 239144 24526 239200
rect 24694 239144 26918 239200
rect 27086 239144 29218 239200
rect 29386 239144 31610 239200
rect 31778 239144 34002 239200
rect 34170 239144 36302 239200
rect 36470 239144 38694 239200
rect 38862 239144 40994 239200
rect 41162 239144 43386 239200
rect 43554 239144 45686 239200
rect 45854 239144 48078 239200
rect 48246 239144 50470 239200
rect 50638 239144 52770 239200
rect 52938 239144 55162 239200
rect 55330 239144 57462 239200
rect 57630 239144 59854 239200
rect 60022 239144 62154 239200
rect 62322 239144 64546 239200
rect 64714 239144 66938 239200
rect 67106 239144 69238 239200
rect 69406 239144 71630 239200
rect 71798 239144 73930 239200
rect 74098 239144 76322 239200
rect 76490 239144 78622 239200
rect 78790 239144 81014 239200
rect 81182 239144 83406 239200
rect 83574 239144 85706 239200
rect 85874 239144 88098 239200
rect 88266 239144 90398 239200
rect 90566 239144 92790 239200
rect 92958 239144 95090 239200
rect 95258 239144 97482 239200
rect 97650 239144 99874 239200
rect 100042 239144 102174 239200
rect 102342 239144 104566 239200
rect 104734 239144 106866 239200
rect 107034 239144 109258 239200
rect 109426 239144 111558 239200
rect 111726 239144 113950 239200
rect 114118 239144 116342 239200
rect 116510 239144 118642 239200
rect 118810 239144 121034 239200
rect 121202 239144 123334 239200
rect 123502 239144 125726 239200
rect 125894 239144 128026 239200
rect 128194 239144 130418 239200
rect 130586 239144 132810 239200
rect 132978 239144 135110 239200
rect 135278 239144 137502 239200
rect 137670 239144 139802 239200
rect 139970 239144 142194 239200
rect 142362 239144 144494 239200
rect 144662 239144 146886 239200
rect 147054 239144 149278 239200
rect 149446 239144 151578 239200
rect 151746 239144 153970 239200
rect 154138 239144 156270 239200
rect 156438 239144 158662 239200
rect 158830 239144 160962 239200
rect 161130 239144 163354 239200
rect 163522 239144 165746 239200
rect 165914 239144 168046 239200
rect 168214 239144 170438 239200
rect 170606 239144 172738 239200
rect 172906 239144 175130 239200
rect 175298 239144 177430 239200
rect 177598 239144 179822 239200
rect 179990 239144 182214 239200
rect 182382 239144 184514 239200
rect 184682 239144 186906 239200
rect 187074 239144 189206 239200
rect 189374 239144 191598 239200
rect 191766 239144 193898 239200
rect 194066 239144 196290 239200
rect 196458 239144 198682 239200
rect 198850 239144 200982 239200
rect 201150 239144 203374 239200
rect 203542 239144 205674 239200
rect 205842 239144 208066 239200
rect 208234 239144 210366 239200
rect 210534 239144 212758 239200
rect 212926 239144 215150 239200
rect 215318 239144 217450 239200
rect 217618 239144 219842 239200
rect 220010 239144 222142 239200
rect 222310 239144 224534 239200
rect 224702 239144 226834 239200
rect 227002 239144 229226 239200
rect 229394 239144 231618 239200
rect 231786 239144 233918 239200
rect 234086 239144 236310 239200
rect 236478 239144 238610 239200
rect 238778 239144 241002 239200
rect 241170 239144 243302 239200
rect 243470 239144 245694 239200
rect 245862 239144 248086 239200
rect 248254 239144 250386 239200
rect 250554 239144 252778 239200
rect 252946 239144 255078 239200
rect 255246 239144 257470 239200
rect 257638 239144 259770 239200
rect 259938 239144 262162 239200
rect 262330 239144 264554 239200
rect 264722 239144 266854 239200
rect 267022 239144 269246 239200
rect 269414 239144 271546 239200
rect 271714 239144 273938 239200
rect 274106 239144 276238 239200
rect 276406 239144 278630 239200
rect 296 856 278740 239144
rect 406 800 790 856
rect 958 800 1342 856
rect 1510 800 1894 856
rect 2062 800 2446 856
rect 2614 800 2998 856
rect 3166 800 3550 856
rect 3718 800 4102 856
rect 4270 800 4654 856
rect 4822 800 5206 856
rect 5374 800 5758 856
rect 5926 800 6310 856
rect 6478 800 6862 856
rect 7030 800 7414 856
rect 7582 800 8058 856
rect 8226 800 8610 856
rect 8778 800 9162 856
rect 9330 800 9714 856
rect 9882 800 10266 856
rect 10434 800 10818 856
rect 10986 800 11370 856
rect 11538 800 11922 856
rect 12090 800 12474 856
rect 12642 800 13026 856
rect 13194 800 13578 856
rect 13746 800 14130 856
rect 14298 800 14682 856
rect 14850 800 15234 856
rect 15402 800 15878 856
rect 16046 800 16430 856
rect 16598 800 16982 856
rect 17150 800 17534 856
rect 17702 800 18086 856
rect 18254 800 18638 856
rect 18806 800 19190 856
rect 19358 800 19742 856
rect 19910 800 20294 856
rect 20462 800 20846 856
rect 21014 800 21398 856
rect 21566 800 21950 856
rect 22118 800 22502 856
rect 22670 800 23146 856
rect 23314 800 23698 856
rect 23866 800 24250 856
rect 24418 800 24802 856
rect 24970 800 25354 856
rect 25522 800 25906 856
rect 26074 800 26458 856
rect 26626 800 27010 856
rect 27178 800 27562 856
rect 27730 800 28114 856
rect 28282 800 28666 856
rect 28834 800 29218 856
rect 29386 800 29770 856
rect 29938 800 30322 856
rect 30490 800 30966 856
rect 31134 800 31518 856
rect 31686 800 32070 856
rect 32238 800 32622 856
rect 32790 800 33174 856
rect 33342 800 33726 856
rect 33894 800 34278 856
rect 34446 800 34830 856
rect 34998 800 35382 856
rect 35550 800 35934 856
rect 36102 800 36486 856
rect 36654 800 37038 856
rect 37206 800 37590 856
rect 37758 800 38234 856
rect 38402 800 38786 856
rect 38954 800 39338 856
rect 39506 800 39890 856
rect 40058 800 40442 856
rect 40610 800 40994 856
rect 41162 800 41546 856
rect 41714 800 42098 856
rect 42266 800 42650 856
rect 42818 800 43202 856
rect 43370 800 43754 856
rect 43922 800 44306 856
rect 44474 800 44858 856
rect 45026 800 45410 856
rect 45578 800 46054 856
rect 46222 800 46606 856
rect 46774 800 47158 856
rect 47326 800 47710 856
rect 47878 800 48262 856
rect 48430 800 48814 856
rect 48982 800 49366 856
rect 49534 800 49918 856
rect 50086 800 50470 856
rect 50638 800 51022 856
rect 51190 800 51574 856
rect 51742 800 52126 856
rect 52294 800 52678 856
rect 52846 800 53322 856
rect 53490 800 53874 856
rect 54042 800 54426 856
rect 54594 800 54978 856
rect 55146 800 55530 856
rect 55698 800 56082 856
rect 56250 800 56634 856
rect 56802 800 57186 856
rect 57354 800 57738 856
rect 57906 800 58290 856
rect 58458 800 58842 856
rect 59010 800 59394 856
rect 59562 800 59946 856
rect 60114 800 60498 856
rect 60666 800 61142 856
rect 61310 800 61694 856
rect 61862 800 62246 856
rect 62414 800 62798 856
rect 62966 800 63350 856
rect 63518 800 63902 856
rect 64070 800 64454 856
rect 64622 800 65006 856
rect 65174 800 65558 856
rect 65726 800 66110 856
rect 66278 800 66662 856
rect 66830 800 67214 856
rect 67382 800 67766 856
rect 67934 800 68410 856
rect 68578 800 68962 856
rect 69130 800 69514 856
rect 69682 800 70066 856
rect 70234 800 70618 856
rect 70786 800 71170 856
rect 71338 800 71722 856
rect 71890 800 72274 856
rect 72442 800 72826 856
rect 72994 800 73378 856
rect 73546 800 73930 856
rect 74098 800 74482 856
rect 74650 800 75034 856
rect 75202 800 75586 856
rect 75754 800 76230 856
rect 76398 800 76782 856
rect 76950 800 77334 856
rect 77502 800 77886 856
rect 78054 800 78438 856
rect 78606 800 78990 856
rect 79158 800 79542 856
rect 79710 800 80094 856
rect 80262 800 80646 856
rect 80814 800 81198 856
rect 81366 800 81750 856
rect 81918 800 82302 856
rect 82470 800 82854 856
rect 83022 800 83498 856
rect 83666 800 84050 856
rect 84218 800 84602 856
rect 84770 800 85154 856
rect 85322 800 85706 856
rect 85874 800 86258 856
rect 86426 800 86810 856
rect 86978 800 87362 856
rect 87530 800 87914 856
rect 88082 800 88466 856
rect 88634 800 89018 856
rect 89186 800 89570 856
rect 89738 800 90122 856
rect 90290 800 90674 856
rect 90842 800 91318 856
rect 91486 800 91870 856
rect 92038 800 92422 856
rect 92590 800 92974 856
rect 93142 800 93526 856
rect 93694 800 94078 856
rect 94246 800 94630 856
rect 94798 800 95182 856
rect 95350 800 95734 856
rect 95902 800 96286 856
rect 96454 800 96838 856
rect 97006 800 97390 856
rect 97558 800 97942 856
rect 98110 800 98494 856
rect 98662 800 99138 856
rect 99306 800 99690 856
rect 99858 800 100242 856
rect 100410 800 100794 856
rect 100962 800 101346 856
rect 101514 800 101898 856
rect 102066 800 102450 856
rect 102618 800 103002 856
rect 103170 800 103554 856
rect 103722 800 104106 856
rect 104274 800 104658 856
rect 104826 800 105210 856
rect 105378 800 105762 856
rect 105930 800 106406 856
rect 106574 800 106958 856
rect 107126 800 107510 856
rect 107678 800 108062 856
rect 108230 800 108614 856
rect 108782 800 109166 856
rect 109334 800 109718 856
rect 109886 800 110270 856
rect 110438 800 110822 856
rect 110990 800 111374 856
rect 111542 800 111926 856
rect 112094 800 112478 856
rect 112646 800 113030 856
rect 113198 800 113582 856
rect 113750 800 114226 856
rect 114394 800 114778 856
rect 114946 800 115330 856
rect 115498 800 115882 856
rect 116050 800 116434 856
rect 116602 800 116986 856
rect 117154 800 117538 856
rect 117706 800 118090 856
rect 118258 800 118642 856
rect 118810 800 119194 856
rect 119362 800 119746 856
rect 119914 800 120298 856
rect 120466 800 120850 856
rect 121018 800 121494 856
rect 121662 800 122046 856
rect 122214 800 122598 856
rect 122766 800 123150 856
rect 123318 800 123702 856
rect 123870 800 124254 856
rect 124422 800 124806 856
rect 124974 800 125358 856
rect 125526 800 125910 856
rect 126078 800 126462 856
rect 126630 800 127014 856
rect 127182 800 127566 856
rect 127734 800 128118 856
rect 128286 800 128670 856
rect 128838 800 129314 856
rect 129482 800 129866 856
rect 130034 800 130418 856
rect 130586 800 130970 856
rect 131138 800 131522 856
rect 131690 800 132074 856
rect 132242 800 132626 856
rect 132794 800 133178 856
rect 133346 800 133730 856
rect 133898 800 134282 856
rect 134450 800 134834 856
rect 135002 800 135386 856
rect 135554 800 135938 856
rect 136106 800 136582 856
rect 136750 800 137134 856
rect 137302 800 137686 856
rect 137854 800 138238 856
rect 138406 800 138790 856
rect 138958 800 139342 856
rect 139510 800 139894 856
rect 140062 800 140446 856
rect 140614 800 140998 856
rect 141166 800 141550 856
rect 141718 800 142102 856
rect 142270 800 142654 856
rect 142822 800 143206 856
rect 143374 800 143758 856
rect 143926 800 144402 856
rect 144570 800 144954 856
rect 145122 800 145506 856
rect 145674 800 146058 856
rect 146226 800 146610 856
rect 146778 800 147162 856
rect 147330 800 147714 856
rect 147882 800 148266 856
rect 148434 800 148818 856
rect 148986 800 149370 856
rect 149538 800 149922 856
rect 150090 800 150474 856
rect 150642 800 151026 856
rect 151194 800 151670 856
rect 151838 800 152222 856
rect 152390 800 152774 856
rect 152942 800 153326 856
rect 153494 800 153878 856
rect 154046 800 154430 856
rect 154598 800 154982 856
rect 155150 800 155534 856
rect 155702 800 156086 856
rect 156254 800 156638 856
rect 156806 800 157190 856
rect 157358 800 157742 856
rect 157910 800 158294 856
rect 158462 800 158846 856
rect 159014 800 159490 856
rect 159658 800 160042 856
rect 160210 800 160594 856
rect 160762 800 161146 856
rect 161314 800 161698 856
rect 161866 800 162250 856
rect 162418 800 162802 856
rect 162970 800 163354 856
rect 163522 800 163906 856
rect 164074 800 164458 856
rect 164626 800 165010 856
rect 165178 800 165562 856
rect 165730 800 166114 856
rect 166282 800 166758 856
rect 166926 800 167310 856
rect 167478 800 167862 856
rect 168030 800 168414 856
rect 168582 800 168966 856
rect 169134 800 169518 856
rect 169686 800 170070 856
rect 170238 800 170622 856
rect 170790 800 171174 856
rect 171342 800 171726 856
rect 171894 800 172278 856
rect 172446 800 172830 856
rect 172998 800 173382 856
rect 173550 800 173934 856
rect 174102 800 174578 856
rect 174746 800 175130 856
rect 175298 800 175682 856
rect 175850 800 176234 856
rect 176402 800 176786 856
rect 176954 800 177338 856
rect 177506 800 177890 856
rect 178058 800 178442 856
rect 178610 800 178994 856
rect 179162 800 179546 856
rect 179714 800 180098 856
rect 180266 800 180650 856
rect 180818 800 181202 856
rect 181370 800 181846 856
rect 182014 800 182398 856
rect 182566 800 182950 856
rect 183118 800 183502 856
rect 183670 800 184054 856
rect 184222 800 184606 856
rect 184774 800 185158 856
rect 185326 800 185710 856
rect 185878 800 186262 856
rect 186430 800 186814 856
rect 186982 800 187366 856
rect 187534 800 187918 856
rect 188086 800 188470 856
rect 188638 800 189022 856
rect 189190 800 189666 856
rect 189834 800 190218 856
rect 190386 800 190770 856
rect 190938 800 191322 856
rect 191490 800 191874 856
rect 192042 800 192426 856
rect 192594 800 192978 856
rect 193146 800 193530 856
rect 193698 800 194082 856
rect 194250 800 194634 856
rect 194802 800 195186 856
rect 195354 800 195738 856
rect 195906 800 196290 856
rect 196458 800 196842 856
rect 197010 800 197486 856
rect 197654 800 198038 856
rect 198206 800 198590 856
rect 198758 800 199142 856
rect 199310 800 199694 856
rect 199862 800 200246 856
rect 200414 800 200798 856
rect 200966 800 201350 856
rect 201518 800 201902 856
rect 202070 800 202454 856
rect 202622 800 203006 856
rect 203174 800 203558 856
rect 203726 800 204110 856
rect 204278 800 204754 856
rect 204922 800 205306 856
rect 205474 800 205858 856
rect 206026 800 206410 856
rect 206578 800 206962 856
rect 207130 800 207514 856
rect 207682 800 208066 856
rect 208234 800 208618 856
rect 208786 800 209170 856
rect 209338 800 209722 856
rect 209890 800 210274 856
rect 210442 800 210826 856
rect 210994 800 211378 856
rect 211546 800 211930 856
rect 212098 800 212574 856
rect 212742 800 213126 856
rect 213294 800 213678 856
rect 213846 800 214230 856
rect 214398 800 214782 856
rect 214950 800 215334 856
rect 215502 800 215886 856
rect 216054 800 216438 856
rect 216606 800 216990 856
rect 217158 800 217542 856
rect 217710 800 218094 856
rect 218262 800 218646 856
rect 218814 800 219198 856
rect 219366 800 219842 856
rect 220010 800 220394 856
rect 220562 800 220946 856
rect 221114 800 221498 856
rect 221666 800 222050 856
rect 222218 800 222602 856
rect 222770 800 223154 856
rect 223322 800 223706 856
rect 223874 800 224258 856
rect 224426 800 224810 856
rect 224978 800 225362 856
rect 225530 800 225914 856
rect 226082 800 226466 856
rect 226634 800 227018 856
rect 227186 800 227662 856
rect 227830 800 228214 856
rect 228382 800 228766 856
rect 228934 800 229318 856
rect 229486 800 229870 856
rect 230038 800 230422 856
rect 230590 800 230974 856
rect 231142 800 231526 856
rect 231694 800 232078 856
rect 232246 800 232630 856
rect 232798 800 233182 856
rect 233350 800 233734 856
rect 233902 800 234286 856
rect 234454 800 234930 856
rect 235098 800 235482 856
rect 235650 800 236034 856
rect 236202 800 236586 856
rect 236754 800 237138 856
rect 237306 800 237690 856
rect 237858 800 238242 856
rect 238410 800 238794 856
rect 238962 800 239346 856
rect 239514 800 239898 856
rect 240066 800 240450 856
rect 240618 800 241002 856
rect 241170 800 241554 856
rect 241722 800 242106 856
rect 242274 800 242750 856
rect 242918 800 243302 856
rect 243470 800 243854 856
rect 244022 800 244406 856
rect 244574 800 244958 856
rect 245126 800 245510 856
rect 245678 800 246062 856
rect 246230 800 246614 856
rect 246782 800 247166 856
rect 247334 800 247718 856
rect 247886 800 248270 856
rect 248438 800 248822 856
rect 248990 800 249374 856
rect 249542 800 250018 856
rect 250186 800 250570 856
rect 250738 800 251122 856
rect 251290 800 251674 856
rect 251842 800 252226 856
rect 252394 800 252778 856
rect 252946 800 253330 856
rect 253498 800 253882 856
rect 254050 800 254434 856
rect 254602 800 254986 856
rect 255154 800 255538 856
rect 255706 800 256090 856
rect 256258 800 256642 856
rect 256810 800 257194 856
rect 257362 800 257838 856
rect 258006 800 258390 856
rect 258558 800 258942 856
rect 259110 800 259494 856
rect 259662 800 260046 856
rect 260214 800 260598 856
rect 260766 800 261150 856
rect 261318 800 261702 856
rect 261870 800 262254 856
rect 262422 800 262806 856
rect 262974 800 263358 856
rect 263526 800 263910 856
rect 264078 800 264462 856
rect 264630 800 265106 856
rect 265274 800 265658 856
rect 265826 800 266210 856
rect 266378 800 266762 856
rect 266930 800 267314 856
rect 267482 800 267866 856
rect 268034 800 268418 856
rect 268586 800 268970 856
rect 269138 800 269522 856
rect 269690 800 270074 856
rect 270242 800 270626 856
rect 270794 800 271178 856
rect 271346 800 271730 856
rect 271898 800 272282 856
rect 272450 800 272926 856
rect 273094 800 273478 856
rect 273646 800 274030 856
rect 274198 800 274582 856
rect 274750 800 275134 856
rect 275302 800 275686 856
rect 275854 800 276238 856
rect 276406 800 276790 856
rect 276958 800 277342 856
rect 277510 800 277894 856
rect 278062 800 278446 856
rect 278614 800 278740 856
<< metal3 >>
rect 279200 226584 280000 226704
rect 0 219920 800 220040
rect 279200 199928 280000 200048
rect 0 179936 800 180056
rect 279200 173272 280000 173392
rect 279200 146616 280000 146736
rect 0 139952 800 140072
rect 279200 119960 280000 120080
rect 0 99968 800 100088
rect 279200 93304 280000 93424
rect 279200 66648 280000 66768
rect 0 59984 800 60104
rect 279200 39992 280000 40112
rect 0 20000 800 20120
rect 279200 13336 280000 13456
<< obsm3 >>
rect 800 220120 265648 237761
rect 880 219840 265648 220120
rect 800 180136 265648 219840
rect 880 179856 265648 180136
rect 800 140152 265648 179856
rect 880 139872 265648 140152
rect 800 100168 265648 139872
rect 880 99888 265648 100168
rect 800 60184 265648 99888
rect 880 59904 265648 60184
rect 800 20200 265648 59904
rect 880 19920 265648 20200
rect 800 2143 265648 19920
<< metal4 >>
rect 4208 2128 4528 237776
rect 4868 2176 5188 237728
rect 5528 2176 5848 237728
rect 6188 2176 6508 237728
rect 19568 2128 19888 237776
rect 20228 2176 20548 237728
rect 20888 2176 21208 237728
rect 21548 2176 21868 237728
rect 34928 2128 35248 237776
rect 35588 2176 35908 237728
rect 36248 2176 36568 237728
rect 36908 2176 37228 237728
rect 50288 2128 50608 237776
rect 50948 2176 51268 237728
rect 51608 2176 51928 237728
rect 52268 2176 52588 237728
rect 65648 2128 65968 237776
rect 66308 2176 66628 237728
rect 66968 2176 67288 237728
rect 67628 2176 67948 237728
rect 81008 2128 81328 237776
rect 81668 2176 81988 237728
rect 82328 2176 82648 237728
rect 82988 2176 83308 237728
rect 96368 2128 96688 237776
rect 97028 2176 97348 237728
rect 97688 2176 98008 237728
rect 98348 2176 98668 237728
rect 111728 2128 112048 237776
rect 112388 2176 112708 237728
rect 113048 2176 113368 237728
rect 113708 2176 114028 237728
rect 127088 2128 127408 237776
rect 127748 2176 128068 237728
rect 128408 2176 128728 237728
rect 129068 2176 129388 237728
rect 142448 2128 142768 237776
rect 143108 2176 143428 237728
rect 143768 2176 144088 237728
rect 144428 2176 144748 237728
rect 157808 2128 158128 237776
rect 158468 2176 158788 237728
rect 159128 2176 159448 237728
rect 159788 2176 160108 237728
rect 173168 2128 173488 237776
rect 173828 2176 174148 237728
rect 174488 2176 174808 237728
rect 175148 2176 175468 237728
rect 188528 2128 188848 237776
rect 189188 2176 189508 237728
rect 189848 2176 190168 237728
rect 190508 2176 190828 237728
rect 203888 2128 204208 237776
rect 204548 2176 204868 237728
rect 205208 2176 205528 237728
rect 205868 2176 206188 237728
rect 219248 2128 219568 237776
rect 219908 2176 220228 237728
rect 220568 2176 220888 237728
rect 221228 2176 221548 237728
rect 234608 2128 234928 237776
rect 235268 2176 235588 237728
rect 235928 2176 236248 237728
rect 236588 2176 236908 237728
rect 249968 2128 250288 237776
rect 250628 2176 250948 237728
rect 251288 2176 251608 237728
rect 251948 2176 252268 237728
rect 265328 2128 265648 237776
rect 265988 2176 266308 237728
rect 266648 2176 266968 237728
rect 267308 2176 267628 237728
<< obsm4 >>
rect 69243 70211 80928 196621
rect 81408 70211 81588 196621
rect 82068 70211 82248 196621
rect 82728 70211 82908 196621
rect 83388 70211 96288 196621
rect 96768 70211 96948 196621
rect 97428 70211 97608 196621
rect 98088 70211 98268 196621
rect 98748 70211 111648 196621
rect 112128 70211 112308 196621
rect 112788 70211 112968 196621
rect 113448 70211 113628 196621
rect 114108 70211 127008 196621
rect 127488 70211 127668 196621
rect 128148 70211 128328 196621
rect 128808 70211 128988 196621
rect 129468 70211 142368 196621
rect 142848 70211 143028 196621
rect 143508 70211 143688 196621
rect 144168 70211 144348 196621
rect 144828 70211 157728 196621
rect 158208 70211 158388 196621
rect 158868 70211 159048 196621
rect 159528 70211 159708 196621
rect 160188 70211 173088 196621
rect 173568 70211 173748 196621
rect 174228 70211 174408 196621
rect 174888 70211 175068 196621
rect 175548 70211 188448 196621
rect 188928 70211 189108 196621
rect 189588 70211 189768 196621
rect 190248 70211 190428 196621
rect 190908 70211 203077 196621
<< labels >>
rlabel metal2 s 274086 0 274142 800 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 279200 93304 280000 93424 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 273994 239200 274050 240000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 276294 0 276350 800 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 279200 119960 280000 120080 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 276294 239200 276350 240000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 276846 0 276902 800 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 277398 0 277454 800 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 59984 800 60104 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 279200 146616 280000 146736 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 277950 0 278006 800 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 274638 0 274694 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 278502 0 278558 800 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 99968 800 100088 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 279200 173272 280000 173392 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 279054 0 279110 800 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 139952 800 140072 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 278686 239200 278742 240000 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 279200 199928 280000 200048 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 279200 226584 280000 226704 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 279606 0 279662 800 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 0 179936 800 180056 6 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal3 s 279200 13336 280000 13456 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s 0 219920 800 220040 6 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal2 s 275190 0 275246 800 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 0 20000 800 20120 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal3 s 279200 39992 280000 40112 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal3 s 279200 66648 280000 66768 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal2 s 269302 239200 269358 240000 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal2 s 275742 0 275798 800 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 271602 239200 271658 240000 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 1122 239200 1178 240000 6 io_in[0]
port 32 nsew signal input
rlabel metal2 s 71686 239200 71742 240000 6 io_in[10]
port 33 nsew signal input
rlabel metal2 s 78678 239200 78734 240000 6 io_in[11]
port 34 nsew signal input
rlabel metal2 s 85762 239200 85818 240000 6 io_in[12]
port 35 nsew signal input
rlabel metal2 s 92846 239200 92902 240000 6 io_in[13]
port 36 nsew signal input
rlabel metal2 s 99930 239200 99986 240000 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 106922 239200 106978 240000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 114006 239200 114062 240000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 121090 239200 121146 240000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 128082 239200 128138 240000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 135166 239200 135222 240000 6 io_in[19]
port 42 nsew signal input
rlabel metal2 s 8114 239200 8170 240000 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 142250 239200 142306 240000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 149334 239200 149390 240000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 156326 239200 156382 240000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 163410 239200 163466 240000 6 io_in[23]
port 47 nsew signal input
rlabel metal2 s 170494 239200 170550 240000 6 io_in[24]
port 48 nsew signal input
rlabel metal2 s 177486 239200 177542 240000 6 io_in[25]
port 49 nsew signal input
rlabel metal2 s 184570 239200 184626 240000 6 io_in[26]
port 50 nsew signal input
rlabel metal2 s 191654 239200 191710 240000 6 io_in[27]
port 51 nsew signal input
rlabel metal2 s 198738 239200 198794 240000 6 io_in[28]
port 52 nsew signal input
rlabel metal2 s 205730 239200 205786 240000 6 io_in[29]
port 53 nsew signal input
rlabel metal2 s 15198 239200 15254 240000 6 io_in[2]
port 54 nsew signal input
rlabel metal2 s 212814 239200 212870 240000 6 io_in[30]
port 55 nsew signal input
rlabel metal2 s 219898 239200 219954 240000 6 io_in[31]
port 56 nsew signal input
rlabel metal2 s 226890 239200 226946 240000 6 io_in[32]
port 57 nsew signal input
rlabel metal2 s 233974 239200 234030 240000 6 io_in[33]
port 58 nsew signal input
rlabel metal2 s 241058 239200 241114 240000 6 io_in[34]
port 59 nsew signal input
rlabel metal2 s 248142 239200 248198 240000 6 io_in[35]
port 60 nsew signal input
rlabel metal2 s 255134 239200 255190 240000 6 io_in[36]
port 61 nsew signal input
rlabel metal2 s 262218 239200 262274 240000 6 io_in[37]
port 62 nsew signal input
rlabel metal2 s 22282 239200 22338 240000 6 io_in[3]
port 63 nsew signal input
rlabel metal2 s 29274 239200 29330 240000 6 io_in[4]
port 64 nsew signal input
rlabel metal2 s 36358 239200 36414 240000 6 io_in[5]
port 65 nsew signal input
rlabel metal2 s 43442 239200 43498 240000 6 io_in[6]
port 66 nsew signal input
rlabel metal2 s 50526 239200 50582 240000 6 io_in[7]
port 67 nsew signal input
rlabel metal2 s 57518 239200 57574 240000 6 io_in[8]
port 68 nsew signal input
rlabel metal2 s 64602 239200 64658 240000 6 io_in[9]
port 69 nsew signal input
rlabel metal2 s 3422 239200 3478 240000 6 io_oeb[0]
port 70 nsew signal output
rlabel metal2 s 73986 239200 74042 240000 6 io_oeb[10]
port 71 nsew signal output
rlabel metal2 s 81070 239200 81126 240000 6 io_oeb[11]
port 72 nsew signal output
rlabel metal2 s 88154 239200 88210 240000 6 io_oeb[12]
port 73 nsew signal output
rlabel metal2 s 95146 239200 95202 240000 6 io_oeb[13]
port 74 nsew signal output
rlabel metal2 s 102230 239200 102286 240000 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 109314 239200 109370 240000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 116398 239200 116454 240000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 123390 239200 123446 240000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 130474 239200 130530 240000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 137558 239200 137614 240000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal2 s 10506 239200 10562 240000 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 144550 239200 144606 240000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 151634 239200 151690 240000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 158718 239200 158774 240000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 165802 239200 165858 240000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal2 s 172794 239200 172850 240000 6 io_oeb[24]
port 86 nsew signal output
rlabel metal2 s 179878 239200 179934 240000 6 io_oeb[25]
port 87 nsew signal output
rlabel metal2 s 186962 239200 187018 240000 6 io_oeb[26]
port 88 nsew signal output
rlabel metal2 s 193954 239200 194010 240000 6 io_oeb[27]
port 89 nsew signal output
rlabel metal2 s 201038 239200 201094 240000 6 io_oeb[28]
port 90 nsew signal output
rlabel metal2 s 208122 239200 208178 240000 6 io_oeb[29]
port 91 nsew signal output
rlabel metal2 s 17590 239200 17646 240000 6 io_oeb[2]
port 92 nsew signal output
rlabel metal2 s 215206 239200 215262 240000 6 io_oeb[30]
port 93 nsew signal output
rlabel metal2 s 222198 239200 222254 240000 6 io_oeb[31]
port 94 nsew signal output
rlabel metal2 s 229282 239200 229338 240000 6 io_oeb[32]
port 95 nsew signal output
rlabel metal2 s 236366 239200 236422 240000 6 io_oeb[33]
port 96 nsew signal output
rlabel metal2 s 243358 239200 243414 240000 6 io_oeb[34]
port 97 nsew signal output
rlabel metal2 s 250442 239200 250498 240000 6 io_oeb[35]
port 98 nsew signal output
rlabel metal2 s 257526 239200 257582 240000 6 io_oeb[36]
port 99 nsew signal output
rlabel metal2 s 264610 239200 264666 240000 6 io_oeb[37]
port 100 nsew signal output
rlabel metal2 s 24582 239200 24638 240000 6 io_oeb[3]
port 101 nsew signal output
rlabel metal2 s 31666 239200 31722 240000 6 io_oeb[4]
port 102 nsew signal output
rlabel metal2 s 38750 239200 38806 240000 6 io_oeb[5]
port 103 nsew signal output
rlabel metal2 s 45742 239200 45798 240000 6 io_oeb[6]
port 104 nsew signal output
rlabel metal2 s 52826 239200 52882 240000 6 io_oeb[7]
port 105 nsew signal output
rlabel metal2 s 59910 239200 59966 240000 6 io_oeb[8]
port 106 nsew signal output
rlabel metal2 s 66994 239200 67050 240000 6 io_oeb[9]
port 107 nsew signal output
rlabel metal2 s 5814 239200 5870 240000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 76378 239200 76434 240000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 83462 239200 83518 240000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 90454 239200 90510 240000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 97538 239200 97594 240000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 104622 239200 104678 240000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 111614 239200 111670 240000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 118698 239200 118754 240000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 125782 239200 125838 240000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 132866 239200 132922 240000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 139858 239200 139914 240000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 12806 239200 12862 240000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 146942 239200 146998 240000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 154026 239200 154082 240000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 161018 239200 161074 240000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 168102 239200 168158 240000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 175186 239200 175242 240000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 182270 239200 182326 240000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 189262 239200 189318 240000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 196346 239200 196402 240000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 203430 239200 203486 240000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 210422 239200 210478 240000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 19890 239200 19946 240000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 217506 239200 217562 240000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 224590 239200 224646 240000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 231674 239200 231730 240000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 238666 239200 238722 240000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 245750 239200 245806 240000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 252834 239200 252890 240000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 259826 239200 259882 240000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 266910 239200 266966 240000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 26974 239200 27030 240000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 34058 239200 34114 240000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 41050 239200 41106 240000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 48134 239200 48190 240000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 55218 239200 55274 240000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 62210 239200 62266 240000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 69294 239200 69350 240000 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 227074 0 227130 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 230478 0 230534 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 235538 0 235594 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 237194 0 237250 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 240506 0 240562 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 242162 0 242218 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 243910 0 243966 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 247222 0 247278 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 248878 0 248934 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 250626 0 250682 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 252282 0 252338 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 253938 0 253994 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 255594 0 255650 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 258998 0 259054 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 260654 0 260710 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 262310 0 262366 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 263966 0 264022 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 265714 0 265770 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 267370 0 267426 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 269026 0 269082 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 270682 0 270738 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 272338 0 272394 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 186870 0 186926 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 193586 0 193642 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 198646 0 198702 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 201958 0 202014 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 205362 0 205418 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 213734 0 213790 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 223762 0 223818 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 227718 0 227774 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 229374 0 229430 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 231030 0 231086 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 232686 0 232742 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 234342 0 234398 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 236090 0 236146 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 237746 0 237802 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 239402 0 239458 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 241058 0 241114 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 242806 0 242862 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 244462 0 244518 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 246118 0 246174 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 247774 0 247830 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 249430 0 249486 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 251178 0 251234 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 252834 0 252890 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 254490 0 254546 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 256146 0 256202 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 257894 0 257950 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 259550 0 259606 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 261206 0 261262 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 262862 0 262918 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 264518 0 264574 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 266266 0 266322 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 267922 0 267978 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 269578 0 269634 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 271234 0 271290 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 272982 0 273038 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 108670 0 108726 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 110326 0 110382 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 120354 0 120410 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 133786 0 133842 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 167366 0 167422 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 169022 0 169078 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 172334 0 172390 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 173990 0 174046 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 177394 0 177450 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 179050 0 179106 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 180706 0 180762 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 182454 0 182510 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 184110 0 184166 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 185766 0 185822 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 187422 0 187478 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 189078 0 189134 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 190826 0 190882 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 192482 0 192538 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 194138 0 194194 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 197542 0 197598 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 200854 0 200910 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 202510 0 202566 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 205914 0 205970 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 207570 0 207626 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 209226 0 209282 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 212630 0 212686 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 214286 0 214342 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 215942 0 215998 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 217598 0 217654 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 219254 0 219310 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 221002 0 221058 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 222658 0 222714 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 224314 0 224370 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 225970 0 226026 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 234986 0 235042 800 6 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 238298 0 238354 800 6 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 239954 0 240010 800 6 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 241610 0 241666 800 6 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 245014 0 245070 800 6 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 248326 0 248382 800 6 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 250074 0 250130 800 6 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 251730 0 251786 800 6 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 255042 0 255098 800 6 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 256698 0 256754 800 6 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 258446 0 258502 800 6 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 261758 0 261814 800 6 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 263414 0 263470 800 6 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 265162 0 265218 800 6 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 266818 0 266874 800 6 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 268474 0 268530 800 6 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 270130 0 270186 800 6 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 271786 0 271842 800 6 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 273534 0 273590 800 6 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 181258 0 181314 800 6 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 183006 0 183062 800 6 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 184662 0 184718 800 6 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 187974 0 188030 800 6 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 189722 0 189778 800 6 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 194690 0 194746 800 6 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 196346 0 196402 800 6 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 201406 0 201462 800 6 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 206466 0 206522 800 6 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 208122 0 208178 800 6 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 211434 0 211490 800 6 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 214838 0 214894 800 6 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 218150 0 218206 800 6 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 223210 0 223266 800 6 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 224866 0 224922 800 6 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 226522 0 226578 800 6 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 530 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 531 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 532 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 wbs_adr_i[0]
port 533 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[10]
port 534 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_adr_i[11]
port 535 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[12]
port 536 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_adr_i[13]
port 537 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[14]
port 538 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[15]
port 539 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_adr_i[16]
port 540 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_adr_i[17]
port 541 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_adr_i[18]
port 542 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[19]
port 543 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[1]
port 544 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_adr_i[20]
port 545 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_adr_i[21]
port 546 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 wbs_adr_i[22]
port 547 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 wbs_adr_i[23]
port 548 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wbs_adr_i[24]
port 549 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 wbs_adr_i[25]
port 550 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_adr_i[26]
port 551 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_adr_i[27]
port 552 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_adr_i[28]
port 553 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 wbs_adr_i[29]
port 554 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[2]
port 555 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 wbs_adr_i[30]
port 556 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 wbs_adr_i[31]
port 557 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[3]
port 558 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[4]
port 559 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[5]
port 560 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[6]
port 561 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[7]
port 562 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[8]
port 563 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[9]
port 564 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_cyc_i
port 565 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_i[0]
port 566 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[10]
port 567 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[11]
port 568 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_i[12]
port 569 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_i[13]
port 570 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_i[14]
port 571 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[15]
port 572 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[16]
port 573 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_i[17]
port 574 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_i[18]
port 575 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[19]
port 576 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_i[1]
port 577 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_i[20]
port 578 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_i[21]
port 579 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_dat_i[22]
port 580 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_i[23]
port 581 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_i[24]
port 582 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[25]
port 583 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wbs_dat_i[26]
port 584 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_i[27]
port 585 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_i[28]
port 586 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_i[29]
port 587 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_i[2]
port 588 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_i[30]
port 589 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_i[31]
port 590 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[3]
port 591 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[4]
port 592 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_i[5]
port 593 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[6]
port 594 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[7]
port 595 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[8]
port 596 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[9]
port 597 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_o[0]
port 598 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_o[10]
port 599 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[11]
port 600 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_o[12]
port 601 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[13]
port 602 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[14]
port 603 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[15]
port 604 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[16]
port 605 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_o[17]
port 606 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_o[18]
port 607 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_o[19]
port 608 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_o[1]
port 609 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_o[20]
port 610 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_o[21]
port 611 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 wbs_dat_o[22]
port 612 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_o[23]
port 613 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 wbs_dat_o[24]
port 614 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 wbs_dat_o[25]
port 615 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_o[26]
port 616 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_o[27]
port 617 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_o[28]
port 618 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 wbs_dat_o[29]
port 619 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[2]
port 620 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_o[30]
port 621 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_o[31]
port 622 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[3]
port 623 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_o[4]
port 624 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[5]
port 625 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[6]
port 626 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[7]
port 627 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[8]
port 628 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[9]
port 629 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 wbs_sel_i[0]
port 630 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_sel_i[1]
port 631 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_sel_i[2]
port 632 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_sel_i[3]
port 633 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_stb_i
port 634 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_we_i
port 635 nsew signal input
rlabel metal4 s 249968 2128 250288 237776 6 vccd1
port 636 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 237776 6 vccd1
port 637 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 237776 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 237776 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 237776 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 237776 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 237776 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 237776 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 237776 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 265328 2128 265648 237776 6 vssd1
port 645 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 237776 6 vssd1
port 646 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 237776 6 vssd1
port 647 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 237776 6 vssd1
port 648 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 237776 6 vssd1
port 649 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 237776 6 vssd1
port 650 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 237776 6 vssd1
port 651 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 237776 6 vssd1
port 652 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 237776 6 vssd1
port 653 nsew ground bidirectional
rlabel metal4 s 250628 2176 250948 237728 6 vccd2
port 654 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 237728 6 vccd2
port 655 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 237728 6 vccd2
port 656 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 237728 6 vccd2
port 657 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 237728 6 vccd2
port 658 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 237728 6 vccd2
port 659 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 237728 6 vccd2
port 660 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 237728 6 vccd2
port 661 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 237728 6 vccd2
port 662 nsew power bidirectional
rlabel metal4 s 265988 2176 266308 237728 6 vssd2
port 663 nsew ground bidirectional
rlabel metal4 s 235268 2176 235588 237728 6 vssd2
port 664 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 237728 6 vssd2
port 665 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 237728 6 vssd2
port 666 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 237728 6 vssd2
port 667 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 237728 6 vssd2
port 668 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 237728 6 vssd2
port 669 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 237728 6 vssd2
port 670 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 237728 6 vssd2
port 671 nsew ground bidirectional
rlabel metal4 s 251288 2176 251608 237728 6 vdda1
port 672 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 237728 6 vdda1
port 673 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 237728 6 vdda1
port 674 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 237728 6 vdda1
port 675 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 237728 6 vdda1
port 676 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 237728 6 vdda1
port 677 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 237728 6 vdda1
port 678 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 237728 6 vdda1
port 679 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 237728 6 vdda1
port 680 nsew power bidirectional
rlabel metal4 s 266648 2176 266968 237728 6 vssa1
port 681 nsew ground bidirectional
rlabel metal4 s 235928 2176 236248 237728 6 vssa1
port 682 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 237728 6 vssa1
port 683 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 237728 6 vssa1
port 684 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 237728 6 vssa1
port 685 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 237728 6 vssa1
port 686 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 237728 6 vssa1
port 687 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 237728 6 vssa1
port 688 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 237728 6 vssa1
port 689 nsew ground bidirectional
rlabel metal4 s 251948 2176 252268 237728 6 vdda2
port 690 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 237728 6 vdda2
port 691 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 237728 6 vdda2
port 692 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 237728 6 vdda2
port 693 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 237728 6 vdda2
port 694 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 237728 6 vdda2
port 695 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 237728 6 vdda2
port 696 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 237728 6 vdda2
port 697 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 237728 6 vdda2
port 698 nsew power bidirectional
rlabel metal4 s 267308 2176 267628 237728 6 vssa2
port 699 nsew ground bidirectional
rlabel metal4 s 236588 2176 236908 237728 6 vssa2
port 700 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 237728 6 vssa2
port 701 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 237728 6 vssa2
port 702 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 237728 6 vssa2
port 703 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 237728 6 vssa2
port 704 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 237728 6 vssa2
port 705 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 237728 6 vssa2
port 706 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 237728 6 vssa2
port 707 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 280000 240000
string LEFview TRUE
<< end >>
