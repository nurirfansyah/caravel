* NGSPICE file created from top_astria.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

.subckt top_astria analog_io[0] analog_io[10] analog_io[11] analog_io[12] analog_io[13]
+ analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18] analog_io[19]
+ analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23] analog_io[24]
+ analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[29] analog_io[2]
+ analog_io[30] analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8]
+ analog_io[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0]
+ la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i VPWR VGND
XFILLER_234_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_258_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0985_ _0987_/CLK _1161_/A VGND VGND VPWR VPWR io_out[28] sky130_fd_sc_hd__dfxtp_4
XFILLER_285_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_278_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_254_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_262_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0770_ VGND VGND VPWR VPWR _0770_/HI _1107_/A sky130_fd_sc_hd__conb_1
XFILLER_183_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_277_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0968_ io_out[18] VGND VGND VPWR VPWR la_data_out[18] sky130_fd_sc_hd__buf_2
XFILLER_105_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0899_ VGND VGND VPWR VPWR _0899_/HI _1158_/C sky130_fd_sc_hd__conb_1
XFILLER_88_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_284_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0822_ VGND VGND VPWR VPWR _0822_/HI _1127_/D sky130_fd_sc_hd__conb_1
XFILLER_102_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0753_ VGND VGND VPWR VPWR _0753_/HI _1100_/A sky130_fd_sc_hd__conb_1
XFILLER_196_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0684_ VGND VGND VPWR VPWR _0684_/HI _1072_/C sky130_fd_sc_hd__conb_1
XFILLER_48_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1167_ _1167_/A analog_io[24] _1167_/C _1167_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_65_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1098_ _1098_/A _1098_/B _1098_/C _1098_/Y VGND VGND VPWR VPWR _1098_/Y sky130_fd_sc_hd__nor4_1
XFILLER_80_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_276_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1021_ _1035_/CLK _1021_/D VGND VGND VPWR VPWR wbs_dat_o[7] sky130_fd_sc_hd__dfxtp_4
XFILLER_47_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0805_ VGND VGND VPWR VPWR _0805_/HI _1120_/D sky130_fd_sc_hd__conb_1
XFILLER_11_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0736_ VGND VGND VPWR VPWR _0736_/HI _1093_/B sky130_fd_sc_hd__conb_1
XFILLER_235_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0667_ VGND VGND VPWR VPWR _0667_/HI _1065_/C sky130_fd_sc_hd__conb_1
XFILLER_258_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0598_ VGND VGND VPWR VPWR _0598_/HI la_data_out[106] sky130_fd_sc_hd__conb_1
XFILLER_97_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_5 wb_rst_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0521_ VGND VGND VPWR VPWR _0521_/HI io_out[35] sky130_fd_sc_hd__conb_1
XFILLER_10_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0452_ _0459_/A VGND VGND VPWR VPWR _0452_/X sky130_fd_sc_hd__buf_2
XFILLER_234_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1004_ _1005_/CLK _1085_/A VGND VGND VPWR VPWR io_out[9] sky130_fd_sc_hd__dfxtp_4
XFILLER_63_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0719_ VGND VGND VPWR VPWR _0719_/HI _1086_/C sky130_fd_sc_hd__conb_1
XFILLER_239_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0504_ VGND VGND VPWR VPWR _0504_/HI _1169_/C sky130_fd_sc_hd__conb_1
XFILLER_67_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0984_ _0987_/CLK _1165_/A VGND VGND VPWR VPWR io_out[29] sky130_fd_sc_hd__dfxtp_4
XFILLER_125_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0967_ io_out[17] VGND VGND VPWR VPWR la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_277_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0898_ VGND VGND VPWR VPWR _0898_/HI _1158_/B sky130_fd_sc_hd__conb_1
XFILLER_238_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_262_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0821_ VGND VGND VPWR VPWR _0821_/HI _1127_/C sky130_fd_sc_hd__conb_1
XFILLER_187_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0752_ VGND VGND VPWR VPWR _0752_/HI _1099_/D sky130_fd_sc_hd__conb_1
XFILLER_196_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0683_ VGND VGND VPWR VPWR _0683_/HI _1072_/A sky130_fd_sc_hd__conb_1
XFILLER_192_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1166_ _1165_/Y _1166_/B _1166_/C _1165_/A VGND VGND VPWR VPWR _1165_/A sky130_fd_sc_hd__nor4_1
XFILLER_246_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1097_ _1098_/Y _1097_/B _1097_/C _1098_/A VGND VGND VPWR VPWR _1098_/A sky130_fd_sc_hd__nor4_1
XFILLER_209_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1020_ _1035_/CLK _0481_/X VGND VGND VPWR VPWR wbs_dat_o[6] sky130_fd_sc_hd__dfxtp_4
XFILLER_219_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0804_ VGND VGND VPWR VPWR _0804_/HI _1120_/C sky130_fd_sc_hd__conb_1
XFILLER_278_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0735_ VGND VGND VPWR VPWR _0735_/HI _1092_/D sky130_fd_sc_hd__conb_1
XFILLER_128_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0666_ VGND VGND VPWR VPWR _0666_/HI _1065_/B sky130_fd_sc_hd__conb_1
XFILLER_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0597_ VGND VGND VPWR VPWR _0597_/HI la_data_out[105] sky130_fd_sc_hd__conb_1
XFILLER_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1149_ _1149_/A _1149_/B _1149_/C _1149_/D VGND VGND VPWR VPWR _1149_/D sky130_fd_sc_hd__nor4_1
XFILLER_38_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_267_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0520_ VGND VGND VPWR VPWR _0520_/HI io_out[34] sky130_fd_sc_hd__conb_1
XFILLER_4_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0451_ wbs_dat_o[27] _0450_/X io_out[27] _0444_/X VGND VGND VPWR VPWR _1041_/D sky130_fd_sc_hd__o22a_4
XFILLER_45_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1003_ _1003_/CLK _1089_/A VGND VGND VPWR VPWR io_out[10] sky130_fd_sc_hd__dfxtp_4
XFILLER_267_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0718_ VGND VGND VPWR VPWR _0718_/HI _1086_/B sky130_fd_sc_hd__conb_1
XFILLER_104_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0649_ VGND VGND VPWR VPWR _0649_/HI _1058_/C sky130_fd_sc_hd__conb_1
XFILLER_83_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0503_ VGND VGND VPWR VPWR _0503_/HI _1169_/B sky130_fd_sc_hd__conb_1
XFILLER_99_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0983_ _0987_/CLK _1169_/A VGND VGND VPWR VPWR io_out[30] sky130_fd_sc_hd__dfxtp_4
XFILLER_242_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_270_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0966_ io_out[16] VGND VGND VPWR VPWR la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_118_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0897_ VGND VGND VPWR VPWR _0897_/HI _1157_/C sky130_fd_sc_hd__conb_1
XFILLER_127_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_254_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0820_ VGND VGND VPWR VPWR _0820_/HI _1127_/A sky130_fd_sc_hd__conb_1
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0751_ VGND VGND VPWR VPWR _0751_/HI _1099_/C sky130_fd_sc_hd__conb_1
XFILLER_7_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0682_ VGND VGND VPWR VPWR _0682_/HI _1071_/D sky130_fd_sc_hd__conb_1
XFILLER_183_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1165_ _1165_/A _1165_/B _1165_/C _1165_/Y VGND VGND VPWR VPWR _1165_/Y sky130_fd_sc_hd__nor4_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1096_ _1096_/A analog_io[25] _1096_/C _1096_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_225_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0949_ _0949_/A VGND VGND VPWR VPWR io_oeb[36] sky130_fd_sc_hd__buf_2
XFILLER_107_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0803_ VGND VGND VPWR VPWR _0803_/HI _1120_/A sky130_fd_sc_hd__conb_1
XFILLER_198_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0734_ VGND VGND VPWR VPWR _0734_/HI _1092_/C sky130_fd_sc_hd__conb_1
XFILLER_171_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0665_ VGND VGND VPWR VPWR _0665_/HI _1064_/D sky130_fd_sc_hd__conb_1
XFILLER_217_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0596_ VGND VGND VPWR VPWR _0596_/HI la_data_out[104] sky130_fd_sc_hd__conb_1
XFILLER_48_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1148_ _1148_/A analog_io[25] _1148_/C _1148_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1079_ _1079_/A analog_io[24] _1079_/C _1079_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_94_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0450_ _0449_/X VGND VGND VPWR VPWR _0450_/X sky130_fd_sc_hd__buf_2
XFILLER_49_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1002_ _1005_/CLK _1093_/A VGND VGND VPWR VPWR io_out[11] sky130_fd_sc_hd__dfxtp_4
XFILLER_35_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0717_ VGND VGND VPWR VPWR _0717_/HI _1085_/C sky130_fd_sc_hd__conb_1
XFILLER_102_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0648_ VGND VGND VPWR VPWR _0648_/HI _1058_/B sky130_fd_sc_hd__conb_1
XFILLER_217_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0579_ VGND VGND VPWR VPWR _0579_/HI la_data_out[87] sky130_fd_sc_hd__conb_1
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0502_ VGND VGND VPWR VPWR _0502_/HI _1168_/D sky130_fd_sc_hd__conb_1
XFILLER_141_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_270_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0982_ _0987_/CLK _1173_/A VGND VGND VPWR VPWR io_out[31] sky130_fd_sc_hd__dfxtp_4
XFILLER_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_275_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0965_ io_out[15] VGND VGND VPWR VPWR la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_140_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0896_ VGND VGND VPWR VPWR _0896_/HI _1157_/B sky130_fd_sc_hd__conb_1
XFILLER_105_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_274_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0750_ VGND VGND VPWR VPWR _0750_/HI _1099_/A sky130_fd_sc_hd__conb_1
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0681_ VGND VGND VPWR VPWR _0681_/HI _1071_/C sky130_fd_sc_hd__conb_1
XFILLER_87_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1164_ _1164_/A analog_io[25] _1164_/C _1164_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_226_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1095_ _1095_/A analog_io[24] _1095_/C _1095_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_92_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0948_ _0949_/A VGND VGND VPWR VPWR io_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_174_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0879_ VGND VGND VPWR VPWR _0879_/HI _1150_/C sky130_fd_sc_hd__conb_1
XFILLER_109_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_255_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0802_ VGND VGND VPWR VPWR _0802_/HI _1119_/D sky130_fd_sc_hd__conb_1
XFILLER_50_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0733_ VGND VGND VPWR VPWR _0733_/HI _1092_/A sky130_fd_sc_hd__conb_1
XFILLER_102_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0664_ VGND VGND VPWR VPWR _0664_/HI _1064_/C sky130_fd_sc_hd__conb_1
XFILLER_115_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0595_ VGND VGND VPWR VPWR _0595_/HI la_data_out[103] sky130_fd_sc_hd__conb_1
XFILLER_258_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1147_ _1147_/A analog_io[24] _1147_/C _1147_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1078_ _1077_/Y _1078_/B _1078_/C _1077_/A VGND VGND VPWR VPWR _1077_/A sky130_fd_sc_hd__nor4_1
XFILLER_0_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1001_ _1005_/CLK _1098_/Y VGND VGND VPWR VPWR io_out[12] sky130_fd_sc_hd__dfxtp_4
XFILLER_130_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0716_ VGND VGND VPWR VPWR _0716_/HI _1085_/B sky130_fd_sc_hd__conb_1
XFILLER_237_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0647_ VGND VGND VPWR VPWR _0647_/HI _1057_/C sky130_fd_sc_hd__conb_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0578_ VGND VGND VPWR VPWR _0578_/HI la_data_out[86] sky130_fd_sc_hd__conb_1
XFILLER_140_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0501_ VGND VGND VPWR VPWR _0501_/HI _1168_/C sky130_fd_sc_hd__conb_1
XFILLER_113_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_278_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0981_ io_out[31] VGND VGND VPWR VPWR la_data_out[31] sky130_fd_sc_hd__buf_2
XFILLER_73_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0964_ io_out[14] VGND VGND VPWR VPWR la_data_out[14] sky130_fd_sc_hd__buf_2
XFILLER_203_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0895_ VGND VGND VPWR VPWR _0895_/HI _1156_/D sky130_fd_sc_hd__conb_1
XFILLER_145_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0680_ VGND VGND VPWR VPWR _0680_/HI _1071_/A sky130_fd_sc_hd__conb_1
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1163_ _1163_/A analog_io[24] _1163_/C _1163_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_225_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1094_ _1093_/D _1094_/B _1094_/C _1093_/A VGND VGND VPWR VPWR _1093_/A sky130_fd_sc_hd__nor4_1
XFILLER_98_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0947_ _0949_/A VGND VGND VPWR VPWR io_oeb[34] sky130_fd_sc_hd__buf_2
XFILLER_147_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0878_ VGND VGND VPWR VPWR _0878_/HI _1150_/B sky130_fd_sc_hd__conb_1
XFILLER_118_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0801_ VGND VGND VPWR VPWR _0801_/HI _1119_/C sky130_fd_sc_hd__conb_1
XFILLER_200_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0732_ VGND VGND VPWR VPWR _0732_/HI _1091_/D sky130_fd_sc_hd__conb_1
XFILLER_176_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0663_ VGND VGND VPWR VPWR _0663_/HI _1064_/A sky130_fd_sc_hd__conb_1
XFILLER_115_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0594_ VGND VGND VPWR VPWR _0594_/HI la_data_out[102] sky130_fd_sc_hd__conb_1
XFILLER_83_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1146_ _1145_/D _1146_/B _1146_/C _1145_/A VGND VGND VPWR VPWR _1145_/A sky130_fd_sc_hd__nor4_1
XFILLER_77_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1077_ _1077_/A _1077_/B _1077_/C _1077_/Y VGND VGND VPWR VPWR _1077_/Y sky130_fd_sc_hd__nor4_1
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1000_ _1006_/CLK _1101_/A VGND VGND VPWR VPWR io_out[13] sky130_fd_sc_hd__dfxtp_4
XFILLER_47_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0715_ VGND VGND VPWR VPWR _0715_/HI _1084_/D sky130_fd_sc_hd__conb_1
XFILLER_176_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0646_ VGND VGND VPWR VPWR _0646_/HI _1057_/B sky130_fd_sc_hd__conb_1
XFILLER_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0577_ VGND VGND VPWR VPWR _0577_/HI la_data_out[85] sky130_fd_sc_hd__conb_1
XFILLER_213_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1129_ _1129_/A _1129_/B _1129_/C _1129_/Y VGND VGND VPWR VPWR _1129_/Y sky130_fd_sc_hd__nor4_1
XFILLER_183_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0500_ VGND VGND VPWR VPWR _0500_/HI _1168_/A sky130_fd_sc_hd__conb_1
XFILLER_207_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0629_ VGND VGND VPWR VPWR _0629_/HI _1050_/C sky130_fd_sc_hd__conb_1
XFILLER_252_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0980_ io_out[30] VGND VGND VPWR VPWR la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_203_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_253_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_269_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0963_ io_out[13] VGND VGND VPWR VPWR la_data_out[13] sky130_fd_sc_hd__buf_2
XFILLER_119_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0894_ VGND VGND VPWR VPWR _0894_/HI _1156_/C sky130_fd_sc_hd__conb_1
XFILLER_199_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_252_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_285_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1162_ _1161_/Y _1162_/B _1162_/C _1161_/A VGND VGND VPWR VPWR _1161_/A sky130_fd_sc_hd__nor4_1
XFILLER_49_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1093_ _1093_/A _1093_/B _1093_/C _1093_/D VGND VGND VPWR VPWR _1093_/D sky130_fd_sc_hd__nor4_1
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0946_ _0949_/A VGND VGND VPWR VPWR io_oeb[33] sky130_fd_sc_hd__buf_2
XFILLER_277_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0877_ VGND VGND VPWR VPWR _0877_/HI _1149_/C sky130_fd_sc_hd__conb_1
XFILLER_88_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0800_ VGND VGND VPWR VPWR _0800_/HI _1119_/A sky130_fd_sc_hd__conb_1
XFILLER_180_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0731_ VGND VGND VPWR VPWR _0731_/HI _1091_/C sky130_fd_sc_hd__conb_1
XFILLER_183_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0662_ VGND VGND VPWR VPWR _0662_/HI _1063_/D sky130_fd_sc_hd__conb_1
XFILLER_171_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0593_ VGND VGND VPWR VPWR _0593_/HI la_data_out[101] sky130_fd_sc_hd__conb_1
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1145_ _1145_/A _1145_/B _1145_/C _1145_/D VGND VGND VPWR VPWR _1145_/D sky130_fd_sc_hd__nor4_1
XFILLER_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1076_ _1076_/A analog_io[25] _1076_/C _1076_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_168_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0929_ _0949_/A VGND VGND VPWR VPWR io_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_105_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_262_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_250_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0714_ VGND VGND VPWR VPWR _0714_/HI _1084_/C sky130_fd_sc_hd__conb_1
XFILLER_219_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0645_ VGND VGND VPWR VPWR _0645_/HI _1056_/D sky130_fd_sc_hd__conb_1
XFILLER_48_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0576_ VGND VGND VPWR VPWR _0576_/HI la_data_out[84] sky130_fd_sc_hd__conb_1
XFILLER_217_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1128_ _1128_/A analog_io[25] _1128_/C _1128_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_241_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1059_ _1059_/A analog_io[24] _1059_/C _1059_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_53_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_270_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_268_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0628_ VGND VGND VPWR VPWR _0628_/HI _1050_/B sky130_fd_sc_hd__conb_1
XFILLER_113_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0559_ VGND VGND VPWR VPWR _0559_/HI la_data_out[67] sky130_fd_sc_hd__conb_1
XFILLER_115_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0962_ io_out[12] VGND VGND VPWR VPWR la_data_out[12] sky130_fd_sc_hd__buf_2
XFILLER_229_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0893_ VGND VGND VPWR VPWR _0893_/HI _1156_/A sky130_fd_sc_hd__conb_1
XFILLER_199_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1161_ _1161_/A _1161_/B _1161_/C _1161_/Y VGND VGND VPWR VPWR _1161_/Y sky130_fd_sc_hd__nor4_1
XFILLER_92_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1092_ _1092_/A analog_io[25] _1092_/C _1092_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_59_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0945_ _0949_/A VGND VGND VPWR VPWR io_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_222_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0876_ VGND VGND VPWR VPWR _0876_/HI _1149_/B sky130_fd_sc_hd__conb_1
XFILLER_174_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0730_ VGND VGND VPWR VPWR _0730_/HI _1091_/A sky130_fd_sc_hd__conb_1
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0661_ VGND VGND VPWR VPWR _0661_/HI _1063_/C sky130_fd_sc_hd__conb_1
XFILLER_13_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0592_ VGND VGND VPWR VPWR _0592_/HI la_data_out[100] sky130_fd_sc_hd__conb_1
XFILLER_152_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1144_ _1144_/A analog_io[25] _1144_/C _1144_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1075_ _1075_/A analog_io[24] _1075_/C _1075_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_46_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0928_ _0949_/A VGND VGND VPWR VPWR io_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_222_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0859_ VGND VGND VPWR VPWR _0859_/HI _1142_/C sky130_fd_sc_hd__conb_1
XFILLER_106_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0713_ VGND VGND VPWR VPWR _0713_/HI _1084_/A sky130_fd_sc_hd__conb_1
XFILLER_32_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0644_ VGND VGND VPWR VPWR _0644_/HI _1056_/C sky130_fd_sc_hd__conb_1
XFILLER_176_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0575_ VGND VGND VPWR VPWR _0575_/HI la_data_out[83] sky130_fd_sc_hd__conb_1
XFILLER_135_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1127_ _1127_/A analog_io[24] _1127_/C _1127_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_54_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1058_ _1057_/Y _1058_/B _1058_/C _1057_/A VGND VGND VPWR VPWR _1057_/A sky130_fd_sc_hd__nor4_1
XFILLER_22_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_281_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0627_ VGND VGND VPWR VPWR _0627_/HI _1049_/C sky130_fd_sc_hd__conb_1
XFILLER_63_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0558_ VGND VGND VPWR VPWR _0558_/HI la_data_out[66] sky130_fd_sc_hd__conb_1
XFILLER_285_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0489_ la_data_in[66] la_oen[66] wb_clk_i _0488_/Y VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__o22a_4
XFILLER_280_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0961_ io_out[11] VGND VGND VPWR VPWR la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_92_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0892_ VGND VGND VPWR VPWR _0892_/HI _1155_/D sky130_fd_sc_hd__conb_1
XFILLER_9_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_stoch_adc_comp.clk _1164_/Y VGND VGND VPWR VPWR clkbuf_0_stoch_adc_comp.clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_259_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1160_ _1160_/A analog_io[25] _1160_/C _1160_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_92_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1091_ _1091_/A analog_io[24] _1091_/C _1091_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_225_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0944_ _0949_/A VGND VGND VPWR VPWR io_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_18_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0875_ VGND VGND VPWR VPWR _0875_/HI _1148_/D sky130_fd_sc_hd__conb_1
XFILLER_173_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_259_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0660_ VGND VGND VPWR VPWR _0660_/HI _1063_/A sky130_fd_sc_hd__conb_1
XFILLER_196_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0591_ VGND VGND VPWR VPWR _0591_/HI la_data_out[99] sky130_fd_sc_hd__conb_1
XFILLER_100_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1143_ _1143_/A analog_io[24] _1143_/C _1143_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1074_ _1073_/Y _1074_/B _1074_/C _1073_/A VGND VGND VPWR VPWR _1073_/A sky130_fd_sc_hd__nor4_1
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0927_ _0949_/A VGND VGND VPWR VPWR io_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_179_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0858_ VGND VGND VPWR VPWR _0858_/HI _1142_/B sky130_fd_sc_hd__conb_1
XFILLER_106_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0789_ VGND VGND VPWR VPWR _0789_/HI _1114_/C sky130_fd_sc_hd__conb_1
XFILLER_66_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0712_ VGND VGND VPWR VPWR _0712_/HI _1083_/D sky130_fd_sc_hd__conb_1
XFILLER_7_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0643_ VGND VGND VPWR VPWR _0643_/HI _1056_/A sky130_fd_sc_hd__conb_1
XFILLER_143_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0574_ VGND VGND VPWR VPWR _0574_/HI la_data_out[82] sky130_fd_sc_hd__conb_1
XFILLER_139_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1126_ _1125_/Y _1126_/B _1126_/C _1125_/A VGND VGND VPWR VPWR _1125_/A sky130_fd_sc_hd__nor4_1
XFILLER_54_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1057_ _1057_/A _1057_/B _1057_/C _1057_/Y VGND VGND VPWR VPWR _1057_/Y sky130_fd_sc_hd__nor4_1
XFILLER_181_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_276_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_281_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_251_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0626_ VGND VGND VPWR VPWR _0626_/HI _1049_/B sky130_fd_sc_hd__conb_1
XFILLER_132_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0557_ VGND VGND VPWR VPWR _0557_/HI la_data_out[65] sky130_fd_sc_hd__conb_1
XFILLER_28_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0488_ la_oen[66] VGND VGND VPWR VPWR _0488_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1109_ _1110_/Y _1109_/B _1109_/C _1110_/A VGND VGND VPWR VPWR _1110_/A sky130_fd_sc_hd__nor4_1
XPHY_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_282_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0609_ VGND VGND VPWR VPWR _0609_/HI la_data_out[117] sky130_fd_sc_hd__conb_1
XFILLER_217_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_261_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0960_ io_out[10] VGND VGND VPWR VPWR la_data_out[10] sky130_fd_sc_hd__buf_2
XPHY_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0891_ VGND VGND VPWR VPWR _0891_/HI _1155_/C sky130_fd_sc_hd__conb_1
XFILLER_173_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_stoch_adc_comp.clk clkbuf_2_0_0_stoch_adc_comp.clk/X VGND VGND VPWR
+ VPWR _1035_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1090_ _1089_/D _1090_/B _1090_/C _1089_/A VGND VGND VPWR VPWR _1089_/A sky130_fd_sc_hd__nor4_1
XFILLER_65_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_stoch_adc_comp.clk clkbuf_3_2_0_stoch_adc_comp.clk/A VGND VGND VPWR
+ VPWR _1006_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0943_ _0949_/A VGND VGND VPWR VPWR io_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_220_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0874_ VGND VGND VPWR VPWR _0874_/HI _1148_/C sky130_fd_sc_hd__conb_1
XFILLER_70_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_251_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5_0_stoch_adc_comp.clk clkbuf_3_5_0_stoch_adc_comp.clk/A VGND VGND VPWR
+ VPWR _0989_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_74_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_249_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0590_ VGND VGND VPWR VPWR _0590_/HI la_data_out[98] sky130_fd_sc_hd__conb_1
XFILLER_48_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1142_ _1141_/D _1142_/B _1142_/C _1141_/A VGND VGND VPWR VPWR _1141_/A sky130_fd_sc_hd__nor4_1
XFILLER_253_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1073_ _1073_/A _1073_/B _1073_/C _1073_/Y VGND VGND VPWR VPWR _1073_/Y sky130_fd_sc_hd__nor4_1
XFILLER_65_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0926_ _0949_/A VGND VGND VPWR VPWR io_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_174_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0857_ VGND VGND VPWR VPWR _0857_/HI _1141_/C sky130_fd_sc_hd__conb_1
XFILLER_274_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0788_ VGND VGND VPWR VPWR _0788_/HI _1114_/B sky130_fd_sc_hd__conb_1
Xclkbuf_3_7_0_stoch_adc_comp.clk clkbuf_2_3_0_stoch_adc_comp.clk/X VGND VGND VPWR
+ VPWR _0987_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0711_ VGND VGND VPWR VPWR _0711_/HI _1083_/C sky130_fd_sc_hd__conb_1
XFILLER_184_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0642_ VGND VGND VPWR VPWR _0642_/HI _1055_/D sky130_fd_sc_hd__conb_1
XFILLER_125_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0573_ VGND VGND VPWR VPWR _0573_/HI la_data_out[81] sky130_fd_sc_hd__conb_1
XFILLER_258_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1125_ _1125_/A _1125_/B _1125_/C _1125_/Y VGND VGND VPWR VPWR _1125_/Y sky130_fd_sc_hd__nor4_1
XFILLER_113_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1056_ _1056_/A analog_io[25] _1056_/C _1056_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_228_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0909_ VGND VGND VPWR VPWR _0909_/HI _1162_/C sky130_fd_sc_hd__conb_1
XFILLER_147_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_stoch_adc_comp.clk clkbuf_2_1_0_stoch_adc_comp.clk/A VGND VGND VPWR
+ VPWR clkbuf_2_0_0_stoch_adc_comp.clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0625_ VGND VGND VPWR VPWR _0625_/HI _1048_/D sky130_fd_sc_hd__conb_1
XFILLER_172_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0556_ VGND VGND VPWR VPWR _0556_/HI la_data_out[64] sky130_fd_sc_hd__conb_1
XFILLER_63_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0487_ wbs_dat_o[0] _0449_/X io_out[0] _0459_/A VGND VGND VPWR VPWR _1014_/D sky130_fd_sc_hd__o22a_4
XFILLER_86_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1108_ _1108_/A analog_io[25] _1108_/C _1108_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XPHY_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1039_ _1003_/CLK _1039_/D VGND VGND VPWR VPWR wbs_dat_o[25] sky130_fd_sc_hd__dfxtp_4
XFILLER_81_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_stoch_adc_comp.clk clkbuf_2_3_0_stoch_adc_comp.clk/A VGND VGND VPWR
+ VPWR clkbuf_3_5_0_stoch_adc_comp.clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_194_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_260_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0608_ VGND VGND VPWR VPWR _0608_/HI la_data_out[116] sky130_fd_sc_hd__conb_1
XFILLER_259_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0539_ VGND VGND VPWR VPWR _0539_/HI la_data_out[47] sky130_fd_sc_hd__conb_1
XFILLER_274_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_277_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0890_ VGND VGND VPWR VPWR _0890_/HI _1155_/A sky130_fd_sc_hd__conb_1
XFILLER_220_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_258_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0942_ _0949_/A VGND VGND VPWR VPWR io_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_261_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0873_ VGND VGND VPWR VPWR _0873_/HI _1148_/A sky130_fd_sc_hd__conb_1
XFILLER_277_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0_stoch_adc_comp.clk clkbuf_0_stoch_adc_comp.clk/X VGND VGND VPWR VPWR
+ clkbuf_2_3_0_stoch_adc_comp.clk/A sky130_fd_sc_hd__clkbuf_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1141_ _1141_/A _1141_/B _1141_/C _1141_/D VGND VGND VPWR VPWR _1141_/D sky130_fd_sc_hd__nor4_1
XFILLER_66_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1072_ _1072_/A analog_io[25] _1072_/C _1072_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0925_ _0949_/A VGND VGND VPWR VPWR io_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_267_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0856_ VGND VGND VPWR VPWR _0856_/HI _1141_/B sky130_fd_sc_hd__conb_1
XFILLER_220_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0787_ VGND VGND VPWR VPWR _0787_/HI _1113_/C sky130_fd_sc_hd__conb_1
XFILLER_143_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0710_ VGND VGND VPWR VPWR _0710_/HI _1083_/A sky130_fd_sc_hd__conb_1
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0641_ VGND VGND VPWR VPWR _0641_/HI _1055_/C sky130_fd_sc_hd__conb_1
XFILLER_125_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0572_ VGND VGND VPWR VPWR _0572_/HI la_data_out[80] sky130_fd_sc_hd__conb_1
XFILLER_174_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1124_ _1124_/A analog_io[25] _1124_/C _1124_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_20_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1055_ _1055_/A analog_io[24] _1055_/C _1055_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_213_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0908_ VGND VGND VPWR VPWR _0908_/HI _1162_/B sky130_fd_sc_hd__conb_1
XFILLER_174_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0839_ VGND VGND VPWR VPWR _0839_/HI _1134_/C sky130_fd_sc_hd__conb_1
XFILLER_200_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0624_ VGND VGND VPWR VPWR _0624_/HI _1048_/C sky130_fd_sc_hd__conb_1
XFILLER_119_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0555_ VGND VGND VPWR VPWR _0555_/HI la_data_out[63] sky130_fd_sc_hd__conb_1
XFILLER_285_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0486_ wbs_dat_o[1] _0449_/X io_out[1] _0459_/A VGND VGND VPWR VPWR _0486_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1107_ _1107_/A analog_io[24] _1107_/C _1107_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_242_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1038_ _1003_/CLK _0455_/X VGND VGND VPWR VPWR wbs_dat_o[24] sky130_fd_sc_hd__dfxtp_4
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_268_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0607_ VGND VGND VPWR VPWR _0607_/HI la_data_out[115] sky130_fd_sc_hd__conb_1
XFILLER_99_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0538_ VGND VGND VPWR VPWR _0538_/HI la_data_out[46] sky130_fd_sc_hd__conb_1
XFILLER_274_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0469_ wbs_dat_o[14] _0464_/X io_out[14] _0466_/X VGND VGND VPWR VPWR _1028_/D sky130_fd_sc_hd__o22a_4
XFILLER_255_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_256_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_269_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_265_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ _0949_/A VGND VGND VPWR VPWR io_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_207_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0872_ VGND VGND VPWR VPWR _0872_/HI _1147_/D sky130_fd_sc_hd__conb_1
XFILLER_179_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1140_ _1140_/A analog_io[25] _1140_/C _1140_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_172_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1071_ _1071_/A analog_io[24] _1071_/C _1071_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_248_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0924_ _0949_/A VGND VGND VPWR VPWR io_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_146_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0855_ VGND VGND VPWR VPWR _0855_/HI _1140_/D sky130_fd_sc_hd__conb_1
XFILLER_140_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0786_ VGND VGND VPWR VPWR _0786_/HI _1113_/B sky130_fd_sc_hd__conb_1
XFILLER_255_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0640_ VGND VGND VPWR VPWR _0640_/HI _1055_/A sky130_fd_sc_hd__conb_1
XFILLER_171_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0571_ VGND VGND VPWR VPWR _0571_/HI la_data_out[79] sky130_fd_sc_hd__conb_1
XFILLER_87_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1123_ _1123_/A analog_io[24] _1123_/C _1123_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_187_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1054_ _1053_/Y _1054_/B _1054_/C _1053_/A VGND VGND VPWR VPWR _1053_/A sky130_fd_sc_hd__nor4_1
XFILLER_0_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0907_ VGND VGND VPWR VPWR _0907_/HI _1161_/C sky130_fd_sc_hd__conb_1
XFILLER_119_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0838_ VGND VGND VPWR VPWR _0838_/HI _1134_/B sky130_fd_sc_hd__conb_1
XFILLER_134_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0769_ VGND VGND VPWR VPWR _0769_/HI _1106_/C sky130_fd_sc_hd__conb_1
XFILLER_1_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0623_ VGND VGND VPWR VPWR _0623_/HI _1048_/A sky130_fd_sc_hd__conb_1
XFILLER_194_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0554_ VGND VGND VPWR VPWR _0554_/HI la_data_out[62] sky130_fd_sc_hd__conb_1
XFILLER_112_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0485_ wbs_dat_o[2] _0449_/X io_out[2] _0480_/X VGND VGND VPWR VPWR _1016_/D sky130_fd_sc_hd__o22a_4
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1106_ _1105_/Y _1106_/B _1106_/C _1105_/A VGND VGND VPWR VPWR _1105_/A sky130_fd_sc_hd__nor4_1
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1037_ _1003_/CLK _1037_/D VGND VGND VPWR VPWR wbs_dat_o[23] sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0606_ VGND VGND VPWR VPWR _0606_/HI la_data_out[114] sky130_fd_sc_hd__conb_1
XFILLER_113_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0537_ VGND VGND VPWR VPWR _0537_/HI la_data_out[45] sky130_fd_sc_hd__conb_1
XFILLER_115_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0468_ wbs_dat_o[15] _0464_/X io_out[15] _0466_/X VGND VGND VPWR VPWR _1029_/D sky130_fd_sc_hd__o22a_4
XFILLER_85_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ _0949_/A VGND VGND VPWR VPWR io_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_186_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0871_ VGND VGND VPWR VPWR _0871_/HI _1147_/C sky130_fd_sc_hd__conb_1
XFILLER_174_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1070_ _1069_/Y _1070_/B _1070_/C _1069_/A VGND VGND VPWR VPWR _1069_/A sky130_fd_sc_hd__nor4_1
XFILLER_280_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0923_ _0949_/A VGND VGND VPWR VPWR io_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_186_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0854_ VGND VGND VPWR VPWR _0854_/HI _1140_/C sky130_fd_sc_hd__conb_1
XFILLER_174_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0785_ VGND VGND VPWR VPWR _0785_/HI _1112_/D sky130_fd_sc_hd__conb_1
XFILLER_128_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0570_ VGND VGND VPWR VPWR _0570_/HI la_data_out[78] sky130_fd_sc_hd__conb_1
XFILLER_152_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1122_ _1122_/A _1122_/B _1122_/C _1122_/Y VGND VGND VPWR VPWR _1122_/Y sky130_fd_sc_hd__nor4_1
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1053_ _1053_/A _1053_/B _1053_/C _1053_/Y VGND VGND VPWR VPWR _1053_/Y sky130_fd_sc_hd__nor4_1
XFILLER_59_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0906_ VGND VGND VPWR VPWR _0906_/HI _1161_/B sky130_fd_sc_hd__conb_1
XFILLER_200_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0837_ VGND VGND VPWR VPWR _0837_/HI _1133_/C sky130_fd_sc_hd__conb_1
XFILLER_278_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0768_ VGND VGND VPWR VPWR _0768_/HI _1106_/B sky130_fd_sc_hd__conb_1
XFILLER_115_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0699_ VGND VGND VPWR VPWR _0699_/HI _1078_/C sky130_fd_sc_hd__conb_1
XFILLER_118_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0622_ VGND VGND VPWR VPWR _0622_/HI _1047_/D sky130_fd_sc_hd__conb_1
XFILLER_256_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0553_ VGND VGND VPWR VPWR _0553_/HI la_data_out[61] sky130_fd_sc_hd__conb_1
XFILLER_119_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0484_ wbs_dat_o[3] _0478_/X io_out[3] _0480_/X VGND VGND VPWR VPWR _0484_/X sky130_fd_sc_hd__o22a_4
XFILLER_140_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1105_ _1105_/A _1105_/B _1105_/C _1105_/Y VGND VGND VPWR VPWR _1105_/Y sky130_fd_sc_hd__nor4_1
XFILLER_54_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1036_ _1035_/CLK _1036_/D VGND VGND VPWR VPWR wbs_dat_o[22] sky130_fd_sc_hd__dfxtp_4
XFILLER_35_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_285_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0605_ VGND VGND VPWR VPWR _0605_/HI la_data_out[113] sky130_fd_sc_hd__conb_1
XFILLER_160_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0536_ VGND VGND VPWR VPWR _0536_/HI la_data_out[44] sky130_fd_sc_hd__conb_1
XFILLER_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0467_ wbs_dat_o[16] _0464_/X io_out[16] _0466_/X VGND VGND VPWR VPWR _0467_/X sky130_fd_sc_hd__o22a_4
XFILLER_45_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1019_ _1035_/CLK _1019_/D VGND VGND VPWR VPWR wbs_dat_o[5] sky130_fd_sc_hd__dfxtp_4
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_260_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_260_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0519_ VGND VGND VPWR VPWR _0519_/HI io_out[33] sky130_fd_sc_hd__conb_1
XFILLER_86_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0870_ VGND VGND VPWR VPWR _0870_/HI _1147_/A sky130_fd_sc_hd__conb_1
XFILLER_35_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0999_ _1006_/CLK _1105_/A VGND VGND VPWR VPWR io_out[14] sky130_fd_sc_hd__dfxtp_4
XFILLER_192_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0922_ _0949_/A VGND VGND VPWR VPWR io_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_226_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0853_ VGND VGND VPWR VPWR _0853_/HI _1140_/A sky130_fd_sc_hd__conb_1
XFILLER_174_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0784_ VGND VGND VPWR VPWR _0784_/HI _1112_/C sky130_fd_sc_hd__conb_1
XFILLER_157_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_262_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1121_ _1122_/Y _1121_/B _1121_/C _1122_/A VGND VGND VPWR VPWR _1122_/A sky130_fd_sc_hd__nor4_1
XFILLER_254_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1052_ _1052_/A analog_io[25] _1052_/C _1052_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_20_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0905_ VGND VGND VPWR VPWR _0905_/HI _1160_/D sky130_fd_sc_hd__conb_1
XFILLER_179_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0836_ VGND VGND VPWR VPWR _0836_/HI _1133_/B sky130_fd_sc_hd__conb_1
XFILLER_190_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0767_ VGND VGND VPWR VPWR _0767_/HI _1105_/C sky130_fd_sc_hd__conb_1
XFILLER_66_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0698_ VGND VGND VPWR VPWR _0698_/HI _1078_/B sky130_fd_sc_hd__conb_1
XFILLER_170_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_263_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_251_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0621_ VGND VGND VPWR VPWR _0621_/HI _1047_/C sky130_fd_sc_hd__conb_1
XFILLER_67_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0552_ VGND VGND VPWR VPWR _0552_/HI la_data_out[60] sky130_fd_sc_hd__conb_1
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0483_ wbs_dat_o[4] _0478_/X io_out[4] _0480_/X VGND VGND VPWR VPWR _1018_/D sky130_fd_sc_hd__o22a_4
XFILLER_267_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1104_ _1104_/A analog_io[25] _1104_/C _1104_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_94_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1035_ _1035_/CLK _1035_/D VGND VGND VPWR VPWR wbs_dat_o[21] sky130_fd_sc_hd__dfxtp_4
XFILLER_165_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0819_ VGND VGND VPWR VPWR _0819_/HI _1126_/C sky130_fd_sc_hd__conb_1
XFILLER_190_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0604_ VGND VGND VPWR VPWR _0604_/HI la_data_out[112] sky130_fd_sc_hd__conb_1
XFILLER_67_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0535_ VGND VGND VPWR VPWR _0535_/HI la_data_out[43] sky130_fd_sc_hd__conb_1
XFILLER_236_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0466_ _0466_/A VGND VGND VPWR VPWR _0466_/X sky130_fd_sc_hd__buf_2
XFILLER_112_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1018_ _1030_/CLK _1018_/D VGND VGND VPWR VPWR wbs_dat_o[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_74_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_277_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_264_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0518_ VGND VGND VPWR VPWR _0518_/HI io_out[32] sky130_fd_sc_hd__conb_1
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0449_ _0464_/A VGND VGND VPWR VPWR _0449_/X sky130_fd_sc_hd__buf_2
XFILLER_67_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0998_ _1006_/CLK _1110_/Y VGND VGND VPWR VPWR io_out[15] sky130_fd_sc_hd__dfxtp_4
XFILLER_160_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ _0949_/A VGND VGND VPWR VPWR io_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_198_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0852_ VGND VGND VPWR VPWR _0852_/HI _1139_/D sky130_fd_sc_hd__conb_1
XFILLER_186_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0783_ VGND VGND VPWR VPWR _0783_/HI _1112_/A sky130_fd_sc_hd__conb_1
XFILLER_31_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1120_ _1120_/A analog_io[25] _1120_/C _1120_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_226_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1051_ _1051_/A analog_io[24] _1051_/C _1051_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0904_ VGND VGND VPWR VPWR _0904_/HI _1160_/C sky130_fd_sc_hd__conb_1
XFILLER_147_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0835_ VGND VGND VPWR VPWR _0835_/HI _1132_/D sky130_fd_sc_hd__conb_1
XFILLER_70_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0766_ VGND VGND VPWR VPWR _0766_/HI _1105_/B sky130_fd_sc_hd__conb_1
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0697_ VGND VGND VPWR VPWR _0697_/HI _1077_/C sky130_fd_sc_hd__conb_1
XFILLER_153_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0620_ VGND VGND VPWR VPWR _0620_/HI _1047_/A sky130_fd_sc_hd__conb_1
XFILLER_125_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0551_ VGND VGND VPWR VPWR _0551_/HI la_data_out[59] sky130_fd_sc_hd__conb_1
XFILLER_256_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0482_ wbs_dat_o[5] _0478_/X io_out[5] _0480_/X VGND VGND VPWR VPWR _1019_/D sky130_fd_sc_hd__o22a_4
XFILLER_80_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1103_ _1103_/A analog_io[24] _1103_/C _1103_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_113_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1034_ _1035_/CLK _1034_/D VGND VGND VPWR VPWR wbs_dat_o[20] sky130_fd_sc_hd__dfxtp_4
XFILLER_78_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0818_ VGND VGND VPWR VPWR _0818_/HI _1126_/B sky130_fd_sc_hd__conb_1
XFILLER_239_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0749_ VGND VGND VPWR VPWR _0749_/HI _1098_/C sky130_fd_sc_hd__conb_1
XFILLER_103_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_283_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_264_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0603_ VGND VGND VPWR VPWR _0603_/HI la_data_out[111] sky130_fd_sc_hd__conb_1
XFILLER_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0534_ VGND VGND VPWR VPWR _0534_/HI la_data_out[42] sky130_fd_sc_hd__conb_1
XFILLER_63_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0465_ wbs_dat_o[17] _0464_/X io_out[17] _0459_/X VGND VGND VPWR VPWR _1031_/D sky130_fd_sc_hd__o22a_4
XFILLER_86_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1017_ _1030_/CLK _0484_/X VGND VGND VPWR VPWR wbs_dat_o[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_240_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_252_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0517_ VGND VGND VPWR VPWR _0517_/HI io_oeb[37] sky130_fd_sc_hd__conb_1
XFILLER_271_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0448_ wbs_dat_o[28] _0442_/X io_out[28] _0444_/X VGND VGND VPWR VPWR _0448_/X sky130_fd_sc_hd__o22a_4
XFILLER_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0997_ _1006_/CLK _1114_/Y VGND VGND VPWR VPWR io_out[16] sky130_fd_sc_hd__dfxtp_4
XFILLER_164_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_254_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ _0949_/A VGND VGND VPWR VPWR io_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_261_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0851_ VGND VGND VPWR VPWR _0851_/HI _1139_/C sky130_fd_sc_hd__conb_1
XFILLER_220_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0782_ VGND VGND VPWR VPWR _0782_/HI _1111_/D sky130_fd_sc_hd__conb_1
XFILLER_31_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_284_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1050_ _1050_/A _1050_/B _1050_/C _1013_/D VGND VGND VPWR VPWR _1013_/D sky130_fd_sc_hd__nor4_1
XFILLER_47_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0903_ VGND VGND VPWR VPWR _0903_/HI _1160_/A sky130_fd_sc_hd__conb_1
XFILLER_187_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0834_ VGND VGND VPWR VPWR _0834_/HI _1132_/C sky130_fd_sc_hd__conb_1
XFILLER_175_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0765_ VGND VGND VPWR VPWR _0765_/HI _1104_/D sky130_fd_sc_hd__conb_1
XFILLER_196_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0696_ VGND VGND VPWR VPWR _0696_/HI _1077_/B sky130_fd_sc_hd__conb_1
XFILLER_131_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_256_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0550_ VGND VGND VPWR VPWR _0550_/HI la_data_out[58] sky130_fd_sc_hd__conb_1
XFILLER_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0481_ wbs_dat_o[6] _0478_/X io_out[6] _0480_/X VGND VGND VPWR VPWR _0481_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1102_ _1101_/Y _1102_/B _1102_/C _1101_/A VGND VGND VPWR VPWR _1101_/A sky130_fd_sc_hd__nor4_1
XFILLER_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1033_ _1035_/CLK _0462_/X VGND VGND VPWR VPWR wbs_dat_o[19] sky130_fd_sc_hd__dfxtp_4
XFILLER_34_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0817_ VGND VGND VPWR VPWR _0817_/HI _1125_/C sky130_fd_sc_hd__conb_1
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0748_ VGND VGND VPWR VPWR _0748_/HI _1098_/B sky130_fd_sc_hd__conb_1
XFILLER_85_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0679_ VGND VGND VPWR VPWR _0679_/HI _1070_/C sky130_fd_sc_hd__conb_1
XFILLER_107_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_252_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_272_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_273_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_279_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_264_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0602_ VGND VGND VPWR VPWR _0602_/HI la_data_out[110] sky130_fd_sc_hd__conb_1
XFILLER_99_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0533_ VGND VGND VPWR VPWR _0533_/HI la_data_out[41] sky130_fd_sc_hd__conb_1
XFILLER_180_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0464_ _0464_/A VGND VGND VPWR VPWR _0464_/X sky130_fd_sc_hd__buf_2
XFILLER_230_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_255_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1016_ _1030_/CLK _1016_/D VGND VGND VPWR VPWR wbs_dat_o[2] sky130_fd_sc_hd__dfxtp_4
XFILLER_223_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0516_ VGND VGND VPWR VPWR _0516_/HI _1174_/C sky130_fd_sc_hd__conb_1
XFILLER_87_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0447_ wbs_dat_o[29] _0442_/X io_out[29] _0444_/X VGND VGND VPWR VPWR _0447_/X sky130_fd_sc_hd__o22a_4
XFILLER_255_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0996_ _1006_/CLK _1117_/A VGND VGND VPWR VPWR io_out[17] sky130_fd_sc_hd__dfxtp_4
XFILLER_146_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0850_ VGND VGND VPWR VPWR _0850_/HI _1139_/A sky130_fd_sc_hd__conb_1
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0781_ VGND VGND VPWR VPWR _0781_/HI _1111_/C sky130_fd_sc_hd__conb_1
XFILLER_196_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0979_ io_out[29] VGND VGND VPWR VPWR la_data_out[29] sky130_fd_sc_hd__buf_2
XFILLER_69_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0902_ VGND VGND VPWR VPWR _0902_/HI _1159_/D sky130_fd_sc_hd__conb_1
XFILLER_202_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0833_ VGND VGND VPWR VPWR _0833_/HI _1132_/A sky130_fd_sc_hd__conb_1
XFILLER_259_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0764_ VGND VGND VPWR VPWR _0764_/HI _1104_/C sky130_fd_sc_hd__conb_1
XFILLER_239_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0695_ VGND VGND VPWR VPWR _0695_/HI _1076_/D sky130_fd_sc_hd__conb_1
XFILLER_48_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_271_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0480_ _0466_/A VGND VGND VPWR VPWR _0480_/X sky130_fd_sc_hd__buf_2
XFILLER_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1101_ _1101_/A _1101_/B _1101_/C _1101_/Y VGND VGND VPWR VPWR _1101_/Y sky130_fd_sc_hd__nor4_1
XFILLER_4_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1032_ _1013_/CLK _1032_/D VGND VGND VPWR VPWR wbs_dat_o[18] sky130_fd_sc_hd__dfxtp_4
XFILLER_47_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0816_ VGND VGND VPWR VPWR _0816_/HI _1125_/B sky130_fd_sc_hd__conb_1
XFILLER_11_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0747_ VGND VGND VPWR VPWR _0747_/HI _1097_/C sky130_fd_sc_hd__conb_1
XFILLER_115_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0678_ VGND VGND VPWR VPWR _0678_/HI _1070_/B sky130_fd_sc_hd__conb_1
XFILLER_258_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_272_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0601_ VGND VGND VPWR VPWR _0601_/HI la_data_out[109] sky130_fd_sc_hd__conb_1
XFILLER_256_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0532_ VGND VGND VPWR VPWR _0532_/HI la_data_out[40] sky130_fd_sc_hd__conb_1
XFILLER_125_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0463_ wbs_dat_o[18] _0457_/X io_out[18] _0459_/X VGND VGND VPWR VPWR _1032_/D sky130_fd_sc_hd__o22a_4
XFILLER_258_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1015_ _1035_/CLK _0486_/X VGND VGND VPWR VPWR wbs_dat_o[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_263_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_260_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0515_ VGND VGND VPWR VPWR _0515_/HI _1174_/B sky130_fd_sc_hd__conb_1
XFILLER_214_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0446_ wbs_dat_o[30] _0442_/X io_out[30] _0444_/X VGND VGND VPWR VPWR _1044_/D sky130_fd_sc_hd__o22a_4
XFILLER_100_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_282_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0995_ _1005_/CLK _1122_/Y VGND VGND VPWR VPWR io_out[18] sky130_fd_sc_hd__dfxtp_4
XFILLER_277_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0780_ VGND VGND VPWR VPWR _0780_/HI _1111_/A sky130_fd_sc_hd__conb_1
XFILLER_220_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0978_ io_out[28] VGND VGND VPWR VPWR la_data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_277_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0901_ VGND VGND VPWR VPWR _0901_/HI _1159_/C sky130_fd_sc_hd__conb_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0832_ VGND VGND VPWR VPWR _0832_/HI _1131_/D sky130_fd_sc_hd__conb_1
XFILLER_31_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0763_ VGND VGND VPWR VPWR _0763_/HI _1104_/A sky130_fd_sc_hd__conb_1
XFILLER_200_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0694_ VGND VGND VPWR VPWR _0694_/HI _1076_/C sky130_fd_sc_hd__conb_1
XFILLER_6_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1100_ _1100_/A analog_io[25] _1100_/C _1100_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_152_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1031_ _1035_/CLK _1031_/D VGND VGND VPWR VPWR wbs_dat_o[17] sky130_fd_sc_hd__dfxtp_4
XFILLER_59_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0815_ VGND VGND VPWR VPWR _0815_/HI _1124_/D sky130_fd_sc_hd__conb_1
XFILLER_174_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0746_ VGND VGND VPWR VPWR _0746_/HI _1097_/B sky130_fd_sc_hd__conb_1
XFILLER_239_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0677_ VGND VGND VPWR VPWR _0677_/HI _1069_/C sky130_fd_sc_hd__conb_1
XFILLER_83_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_272_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0600_ VGND VGND VPWR VPWR _0600_/HI la_data_out[108] sky130_fd_sc_hd__conb_1
XFILLER_201_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0531_ VGND VGND VPWR VPWR _0531_/HI la_data_out[39] sky130_fd_sc_hd__conb_1
XFILLER_259_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0462_ wbs_dat_o[19] _0457_/X io_out[19] _0459_/X VGND VGND VPWR VPWR _0462_/X sky130_fd_sc_hd__o22a_4
XFILLER_45_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1014_ _1035_/CLK _1014_/D VGND VGND VPWR VPWR wbs_dat_o[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_267_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0729_ VGND VGND VPWR VPWR _0729_/HI _1090_/C sky130_fd_sc_hd__conb_1
XFILLER_89_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0514_ VGND VGND VPWR VPWR _0514_/HI _1173_/C sky130_fd_sc_hd__conb_1
XFILLER_80_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0445_ wbs_dat_o[31] _0442_/X io_out[31] _0444_/X VGND VGND VPWR VPWR _0445_/X sky130_fd_sc_hd__o22a_4
XFILLER_41_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_276_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_276_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_261_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0994_ _1005_/CLK _1125_/A VGND VGND VPWR VPWR io_out[19] sky130_fd_sc_hd__dfxtp_4
XFILLER_34_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0977_ io_out[27] VGND VGND VPWR VPWR la_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0900_ VGND VGND VPWR VPWR _0900_/HI _1159_/A sky130_fd_sc_hd__conb_1
XFILLER_226_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0831_ VGND VGND VPWR VPWR _0831_/HI _1131_/C sky130_fd_sc_hd__conb_1
XFILLER_35_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_278_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0762_ VGND VGND VPWR VPWR _0762_/HI _1103_/D sky130_fd_sc_hd__conb_1
XFILLER_227_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0693_ VGND VGND VPWR VPWR _0693_/HI _1076_/A sky130_fd_sc_hd__conb_1
XFILLER_196_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_284_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_277_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1030_ _1030_/CLK _0467_/X VGND VGND VPWR VPWR wbs_dat_o[16] sky130_fd_sc_hd__dfxtp_4
XFILLER_35_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0814_ VGND VGND VPWR VPWR _0814_/HI _1124_/C sky130_fd_sc_hd__conb_1
XFILLER_141_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0745_ VGND VGND VPWR VPWR _0745_/HI _1096_/D sky130_fd_sc_hd__conb_1
XFILLER_171_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0676_ VGND VGND VPWR VPWR _0676_/HI _1069_/B sky130_fd_sc_hd__conb_1
XFILLER_170_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1159_ _1159_/A analog_io[24] _1159_/C _1159_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_240_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0530_ VGND VGND VPWR VPWR _0530_/HI la_data_out[38] sky130_fd_sc_hd__conb_1
XFILLER_99_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0461_ wbs_dat_o[20] _0457_/X io_out[20] _0459_/X VGND VGND VPWR VPWR _1034_/D sky130_fd_sc_hd__o22a_4
XFILLER_65_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1013_ _1013_/CLK _1013_/D VGND VGND VPWR VPWR io_out[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_35_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0728_ VGND VGND VPWR VPWR _0728_/HI _1090_/B sky130_fd_sc_hd__conb_1
XFILLER_274_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0659_ VGND VGND VPWR VPWR _0659_/HI _1062_/C sky130_fd_sc_hd__conb_1
XFILLER_217_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0513_ VGND VGND VPWR VPWR _0513_/HI _1173_/B sky130_fd_sc_hd__conb_1
XFILLER_236_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0444_ _0459_/A VGND VGND VPWR VPWR _0444_/X sky130_fd_sc_hd__buf_2
XFILLER_45_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_269_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0993_ _0987_/CLK _1129_/A VGND VGND VPWR VPWR io_out[20] sky130_fd_sc_hd__dfxtp_4
XFILLER_242_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0976_ io_out[26] VGND VGND VPWR VPWR la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_158_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_254_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_265_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0830_ VGND VGND VPWR VPWR _0830_/HI _1131_/A sky130_fd_sc_hd__conb_1
XFILLER_159_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0761_ VGND VGND VPWR VPWR _0761_/HI _1103_/C sky130_fd_sc_hd__conb_1
XFILLER_31_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0692_ VGND VGND VPWR VPWR _0692_/HI _1075_/D sky130_fd_sc_hd__conb_1
XFILLER_142_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0959_ io_out[9] VGND VGND VPWR VPWR la_data_out[9] sky130_fd_sc_hd__buf_2
XFILLER_88_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0813_ VGND VGND VPWR VPWR _0813_/HI _1124_/A sky130_fd_sc_hd__conb_1
XFILLER_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0744_ VGND VGND VPWR VPWR _0744_/HI _1096_/C sky130_fd_sc_hd__conb_1
XFILLER_102_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0675_ VGND VGND VPWR VPWR _0675_/HI _1068_/D sky130_fd_sc_hd__conb_1
XFILLER_115_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1158_ _1157_/Y _1158_/B _1158_/C _1157_/A VGND VGND VPWR VPWR _1157_/A sky130_fd_sc_hd__nor4_1
XFILLER_168_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1089_ _1089_/A _1089_/B _1089_/C _1089_/D VGND VGND VPWR VPWR _1089_/D sky130_fd_sc_hd__nor4_1
XFILLER_244_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0460_ wbs_dat_o[21] _0457_/X io_out[21] _0459_/X VGND VGND VPWR VPWR _1035_/D sky130_fd_sc_hd__o22a_4
XFILLER_171_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1012_ _1013_/CLK _1053_/A VGND VGND VPWR VPWR io_out[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_130_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0727_ VGND VGND VPWR VPWR _0727_/HI _1089_/C sky130_fd_sc_hd__conb_1
XFILLER_171_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0658_ VGND VGND VPWR VPWR _0658_/HI _1062_/B sky130_fd_sc_hd__conb_1
XFILLER_217_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0589_ VGND VGND VPWR VPWR _0589_/HI la_data_out[97] sky130_fd_sc_hd__conb_1
XFILLER_83_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_285_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0512_ VGND VGND VPWR VPWR _0512_/HI _1172_/D sky130_fd_sc_hd__conb_1
XFILLER_113_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0443_ _0466_/A VGND VGND VPWR VPWR _0459_/A sky130_fd_sc_hd__buf_2
XFILLER_80_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0992_ _1005_/CLK _1133_/A VGND VGND VPWR VPWR io_out[21] sky130_fd_sc_hd__dfxtp_4
XFILLER_13_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_260_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_250_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_284_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0975_ io_out[25] VGND VGND VPWR VPWR la_data_out[25] sky130_fd_sc_hd__buf_2
XFILLER_53_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0760_ VGND VGND VPWR VPWR _0760_/HI _1103_/A sky130_fd_sc_hd__conb_1
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0691_ VGND VGND VPWR VPWR _0691_/HI _1075_/C sky130_fd_sc_hd__conb_1
XFILLER_155_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1174_ _1173_/Y _1174_/B _1174_/C _1173_/A VGND VGND VPWR VPWR _1173_/A sky130_fd_sc_hd__nor4_1
XFILLER_168_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0958_ io_out[8] VGND VGND VPWR VPWR la_data_out[8] sky130_fd_sc_hd__buf_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0889_ VGND VGND VPWR VPWR _0889_/HI _1154_/C sky130_fd_sc_hd__conb_1
XFILLER_284_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0812_ VGND VGND VPWR VPWR _0812_/HI _1123_/D sky130_fd_sc_hd__conb_1
XFILLER_175_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0743_ VGND VGND VPWR VPWR _0743_/HI _1096_/A sky130_fd_sc_hd__conb_1
XFILLER_143_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_254_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0674_ VGND VGND VPWR VPWR _0674_/HI _1068_/C sky130_fd_sc_hd__conb_1
XFILLER_157_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1157_ _1157_/A _1157_/B _1157_/C _1157_/Y VGND VGND VPWR VPWR _1157_/Y sky130_fd_sc_hd__nor4_1
XFILLER_225_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1088_ _1088_/A analog_io[25] _1088_/C _1088_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_34_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1011_ _1013_/CLK _1057_/A VGND VGND VPWR VPWR io_out[2] sky130_fd_sc_hd__dfxtp_4
XFILLER_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0726_ VGND VGND VPWR VPWR _0726_/HI _1089_/B sky130_fd_sc_hd__conb_1
XFILLER_85_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0657_ VGND VGND VPWR VPWR _0657_/HI _1061_/C sky130_fd_sc_hd__conb_1
XFILLER_252_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0588_ VGND VGND VPWR VPWR _0588_/HI la_data_out[96] sky130_fd_sc_hd__conb_1
XFILLER_213_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_257_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_281_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0511_ VGND VGND VPWR VPWR _0511_/HI _1172_/C sky130_fd_sc_hd__conb_1
XFILLER_158_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0442_ _0464_/A VGND VGND VPWR VPWR _0442_/X sky130_fd_sc_hd__buf_2
XFILLER_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_255_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0709_ VGND VGND VPWR VPWR _0709_/HI _1082_/C sky130_fd_sc_hd__conb_1
XFILLER_145_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0991_ _0989_/CLK _1137_/A VGND VGND VPWR VPWR io_out[22] sky130_fd_sc_hd__dfxtp_4
XFILLER_207_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0974_ io_out[24] VGND VGND VPWR VPWR la_data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_119_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0690_ VGND VGND VPWR VPWR _0690_/HI _1075_/A sky130_fd_sc_hd__conb_1
XFILLER_100_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1173_ _1173_/A _1173_/B _1173_/C _1173_/Y VGND VGND VPWR VPWR _1173_/Y sky130_fd_sc_hd__nor4_1
XFILLER_252_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0957_ io_out[7] VGND VGND VPWR VPWR la_data_out[7] sky130_fd_sc_hd__buf_2
XFILLER_146_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0888_ VGND VGND VPWR VPWR _0888_/HI _1154_/B sky130_fd_sc_hd__conb_1
XFILLER_88_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0811_ VGND VGND VPWR VPWR _0811_/HI _1123_/C sky130_fd_sc_hd__conb_1
XFILLER_180_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0742_ VGND VGND VPWR VPWR _0742_/HI _1095_/D sky130_fd_sc_hd__conb_1
XFILLER_196_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0673_ VGND VGND VPWR VPWR _0673_/HI _1068_/A sky130_fd_sc_hd__conb_1
XFILLER_171_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1156_ _1156_/A analog_io[25] _1156_/C _1156_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_38_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1087_ _1087_/A analog_io[24] _1087_/C _1087_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_168_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1010_ _1013_/CLK _1061_/A VGND VGND VPWR VPWR io_out[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_47_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0725_ VGND VGND VPWR VPWR _0725_/HI _1088_/D sky130_fd_sc_hd__conb_1
XFILLER_239_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0656_ VGND VGND VPWR VPWR _0656_/HI _1061_/B sky130_fd_sc_hd__conb_1
XFILLER_256_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0587_ VGND VGND VPWR VPWR _0587_/HI la_data_out[95] sky130_fd_sc_hd__conb_1
XFILLER_217_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1139_ _1139_/A analog_io[24] _1139_/C _1139_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_214_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_281_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0510_ VGND VGND VPWR VPWR _0510_/HI _1172_/A sky130_fd_sc_hd__conb_1
XFILLER_125_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0441_ _0466_/A VGND VGND VPWR VPWR _0464_/A sky130_fd_sc_hd__inv_2
XFILLER_234_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0708_ VGND VGND VPWR VPWR _0708_/HI _1082_/B sky130_fd_sc_hd__conb_1
XFILLER_132_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0639_ VGND VGND VPWR VPWR _0639_/HI _1054_/C sky130_fd_sc_hd__conb_1
XFILLER_258_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0990_ _1005_/CLK _1141_/A VGND VGND VPWR VPWR io_out[23] sky130_fd_sc_hd__dfxtp_4
XFILLER_203_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_253_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0973_ io_out[23] VGND VGND VPWR VPWR la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_146_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_278_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1172_ _1172_/A analog_io[25] _1172_/C _1172_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_38_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0956_ io_out[6] VGND VGND VPWR VPWR la_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_105_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0887_ VGND VGND VPWR VPWR _0887_/HI _1153_/C sky130_fd_sc_hd__conb_1
XFILLER_31_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0810_ VGND VGND VPWR VPWR _0810_/HI _1123_/A sky130_fd_sc_hd__conb_1
XFILLER_30_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0741_ VGND VGND VPWR VPWR _0741_/HI _1095_/C sky130_fd_sc_hd__conb_1
XFILLER_239_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0672_ VGND VGND VPWR VPWR _0672_/HI _1067_/D sky130_fd_sc_hd__conb_1
XFILLER_171_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1155_ _1155_/A analog_io[24] _1155_/C _1155_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_285_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1086_ _1085_/Y _1086_/B _1086_/C _1085_/A VGND VGND VPWR VPWR _1085_/A sky130_fd_sc_hd__nor4_1
XFILLER_283_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0939_ _0949_/A VGND VGND VPWR VPWR io_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_228_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_263_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0724_ VGND VGND VPWR VPWR _0724_/HI _1088_/C sky130_fd_sc_hd__conb_1
XFILLER_155_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0655_ VGND VGND VPWR VPWR _0655_/HI _1060_/D sky130_fd_sc_hd__conb_1
XFILLER_98_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0586_ VGND VGND VPWR VPWR _0586_/HI la_data_out[94] sky130_fd_sc_hd__conb_1
XFILLER_135_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1138_ _1137_/Y _1138_/B _1138_/C _1137_/A VGND VGND VPWR VPWR _1137_/A sky130_fd_sc_hd__nor4_1
XPHY_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1069_ _1069_/A _1069_/B _1069_/C _1069_/Y VGND VGND VPWR VPWR _1069_/Y sky130_fd_sc_hd__nor4_1
XFILLER_230_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_260_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0440_ _0436_/Y _0437_/Y wbs_ack_o _0949_/A VGND VGND VPWR VPWR _0466_/A sky130_fd_sc_hd__or4_4
XFILLER_98_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0707_ VGND VGND VPWR VPWR _0707_/HI _1081_/C sky130_fd_sc_hd__conb_1
XFILLER_137_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0638_ VGND VGND VPWR VPWR _0638_/HI _1054_/B sky130_fd_sc_hd__conb_1
XFILLER_154_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0569_ VGND VGND VPWR VPWR _0569_/HI la_data_out[77] sky130_fd_sc_hd__conb_1
XFILLER_115_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_261_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0972_ io_out[22] VGND VGND VPWR VPWR la_data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_242_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1171_ _1171_/A analog_io[24] _1171_/C _1171_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0955_ io_out[5] VGND VGND VPWR VPWR la_data_out[5] sky130_fd_sc_hd__buf_2
XFILLER_222_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_284_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0886_ VGND VGND VPWR VPWR _0886_/HI _1153_/B sky130_fd_sc_hd__conb_1
XFILLER_174_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0740_ VGND VGND VPWR VPWR _0740_/HI _1095_/A sky130_fd_sc_hd__conb_1
XFILLER_7_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0671_ VGND VGND VPWR VPWR _0671_/HI _1067_/C sky130_fd_sc_hd__conb_1
XFILLER_196_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1154_ _1153_/Y _1154_/B _1154_/C _1153_/A VGND VGND VPWR VPWR _1153_/A sky130_fd_sc_hd__nor4_1
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1085_ _1085_/A _1085_/B _1085_/C _1085_/Y VGND VGND VPWR VPWR _1085_/Y sky130_fd_sc_hd__nor4_1
XFILLER_279_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0938_ _0949_/A VGND VGND VPWR VPWR io_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_140_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0869_ VGND VGND VPWR VPWR _0869_/HI _1146_/C sky130_fd_sc_hd__conb_1
XFILLER_106_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0723_ VGND VGND VPWR VPWR _0723_/HI _1088_/A sky130_fd_sc_hd__conb_1
XFILLER_265_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0654_ VGND VGND VPWR VPWR _0654_/HI _1060_/C sky130_fd_sc_hd__conb_1
XFILLER_217_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0585_ VGND VGND VPWR VPWR _0585_/HI la_data_out[93] sky130_fd_sc_hd__conb_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1137_ _1137_/A _1137_/B _1137_/C _1137_/Y VGND VGND VPWR VPWR _1137_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1068_ _1068_/A analog_io[25] _1068_/C _1068_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_181_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0706_ VGND VGND VPWR VPWR _0706_/HI _1081_/B sky130_fd_sc_hd__conb_1
XFILLER_171_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0637_ VGND VGND VPWR VPWR _0637_/HI _1053_/C sky130_fd_sc_hd__conb_1
XFILLER_132_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0568_ VGND VGND VPWR VPWR _0568_/HI la_data_out[76] sky130_fd_sc_hd__conb_1
XFILLER_58_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0499_ VGND VGND VPWR VPWR _0499_/HI _1167_/D sky130_fd_sc_hd__conb_1
XFILLER_285_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_259_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0971_ io_out[21] VGND VGND VPWR VPWR la_data_out[21] sky130_fd_sc_hd__buf_2
XFILLER_158_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1170_ _1169_/Y _1170_/B _1170_/C _1169_/A VGND VGND VPWR VPWR _1169_/A sky130_fd_sc_hd__nor4_1
XFILLER_77_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0954_ io_out[4] VGND VGND VPWR VPWR la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_192_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0885_ VGND VGND VPWR VPWR _0885_/HI _1152_/D sky130_fd_sc_hd__conb_1
XFILLER_284_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0670_ VGND VGND VPWR VPWR _0670_/HI _1067_/A sky130_fd_sc_hd__conb_1
XFILLER_183_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1153_ _1153_/A _1153_/B _1153_/C _1153_/Y VGND VGND VPWR VPWR _1153_/Y sky130_fd_sc_hd__nor4_1
XFILLER_285_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1084_ _1084_/A analog_io[25] _1084_/C _1084_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_241_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0937_ _0949_/A VGND VGND VPWR VPWR io_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_147_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0868_ VGND VGND VPWR VPWR _0868_/HI _1146_/B sky130_fd_sc_hd__conb_1
XFILLER_173_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0799_ VGND VGND VPWR VPWR _0799_/HI _1118_/C sky130_fd_sc_hd__conb_1
XPHY_8108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0722_ VGND VGND VPWR VPWR _0722_/HI _1087_/D sky130_fd_sc_hd__conb_1
XFILLER_184_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0653_ VGND VGND VPWR VPWR _0653_/HI _1060_/A sky130_fd_sc_hd__conb_1
XFILLER_217_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0584_ VGND VGND VPWR VPWR _0584_/HI la_data_out[92] sky130_fd_sc_hd__conb_1
XFILLER_98_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1136_ _1136_/A analog_io[25] _1136_/C _1136_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_26_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1067_ _1067_/A analog_io[24] _1067_/C _1067_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_230_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_255_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_280_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0705_ VGND VGND VPWR VPWR _0705_/HI _1080_/D sky130_fd_sc_hd__conb_1
XFILLER_258_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0636_ VGND VGND VPWR VPWR _0636_/HI _1053_/B sky130_fd_sc_hd__conb_1
XFILLER_125_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0567_ VGND VGND VPWR VPWR _0567_/HI la_data_out[75] sky130_fd_sc_hd__conb_1
XFILLER_225_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0498_ VGND VGND VPWR VPWR _0498_/HI _1167_/C sky130_fd_sc_hd__conb_1
XFILLER_230_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_273_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ _1119_/A analog_io[24] _1119_/C _1119_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XPHY_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0619_ VGND VGND VPWR VPWR _0619_/HI la_data_out[127] sky130_fd_sc_hd__conb_1
XFILLER_217_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0970_ io_out[20] VGND VGND VPWR VPWR la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_220_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_250_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0953_ io_out[3] VGND VGND VPWR VPWR la_data_out[3] sky130_fd_sc_hd__buf_2
XFILLER_53_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0884_ VGND VGND VPWR VPWR _0884_/HI _1152_/C sky130_fd_sc_hd__conb_1
XFILLER_12_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1152_ _1152_/A analog_io[25] _1152_/C _1152_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_20_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1083_ _1083_/A analog_io[24] _1083_/C _1083_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_34_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0936_ _0949_/A VGND VGND VPWR VPWR io_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_174_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0867_ VGND VGND VPWR VPWR _0867_/HI _1145_/C sky130_fd_sc_hd__conb_1
XFILLER_175_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0798_ VGND VGND VPWR VPWR _0798_/HI _1118_/B sky130_fd_sc_hd__conb_1
XPHY_8109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0721_ VGND VGND VPWR VPWR _0721_/HI _1087_/C sky130_fd_sc_hd__conb_1
XFILLER_184_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0652_ VGND VGND VPWR VPWR _0652_/HI _1059_/D sky130_fd_sc_hd__conb_1
XFILLER_155_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0583_ VGND VGND VPWR VPWR _0583_/HI la_data_out[91] sky130_fd_sc_hd__conb_1
XFILLER_63_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1135_ _1135_/A analog_io[24] _1135_/C _1135_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_20_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1066_ _1065_/Y _1066_/B _1066_/C _1065_/A VGND VGND VPWR VPWR _1065_/A sky130_fd_sc_hd__nor4_1
XFILLER_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0919_ _0949_/A VGND VGND VPWR VPWR io_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_266_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0704_ VGND VGND VPWR VPWR _0704_/HI _1080_/C sky130_fd_sc_hd__conb_1
XFILLER_190_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0635_ VGND VGND VPWR VPWR _0635_/HI _1052_/D sky130_fd_sc_hd__conb_1
XFILLER_131_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0566_ VGND VGND VPWR VPWR _0566_/HI la_data_out[74] sky130_fd_sc_hd__conb_1
XFILLER_213_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0497_ VGND VGND VPWR VPWR _0497_/HI _1167_/A sky130_fd_sc_hd__conb_1
XFILLER_6_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1118_ _1117_/Y _1118_/B _1118_/C _1117_/A VGND VGND VPWR VPWR _1117_/A sky130_fd_sc_hd__nor4_1
XPHY_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1049_ _1013_/D _1049_/B _1049_/C _1050_/A VGND VGND VPWR VPWR _1050_/A sky130_fd_sc_hd__nor4_1
XFILLER_126_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0618_ VGND VGND VPWR VPWR _0618_/HI la_data_out[126] sky130_fd_sc_hd__conb_1
XFILLER_252_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0549_ VGND VGND VPWR VPWR _0549_/HI la_data_out[57] sky130_fd_sc_hd__conb_1
XFILLER_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0952_ io_out[2] VGND VGND VPWR VPWR la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_207_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0883_ VGND VGND VPWR VPWR _0883_/HI _1152_/A sky130_fd_sc_hd__conb_1
XFILLER_140_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1151_ _1151_/A analog_io[24] _1151_/C _1151_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_4_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1082_ _1081_/Y _1082_/B _1082_/C _1081_/A VGND VGND VPWR VPWR _1081_/A sky130_fd_sc_hd__nor4_1
XFILLER_281_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0935_ _0949_/A VGND VGND VPWR VPWR io_oeb[22] sky130_fd_sc_hd__buf_2
XFILLER_146_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0866_ VGND VGND VPWR VPWR _0866_/HI _1145_/B sky130_fd_sc_hd__conb_1
XFILLER_88_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0797_ VGND VGND VPWR VPWR _0797_/HI _1117_/C sky130_fd_sc_hd__conb_1
XFILLER_255_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_280_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0720_ VGND VGND VPWR VPWR _0720_/HI _1087_/A sky130_fd_sc_hd__conb_1
XFILLER_156_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0651_ VGND VGND VPWR VPWR _0651_/HI _1059_/C sky130_fd_sc_hd__conb_1
XFILLER_144_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0582_ VGND VGND VPWR VPWR _0582_/HI la_data_out[90] sky130_fd_sc_hd__conb_1
XFILLER_217_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1134_ _1133_/Y _1134_/B _1134_/C _1133_/A VGND VGND VPWR VPWR _1133_/A sky130_fd_sc_hd__nor4_1
XFILLER_38_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1065_ _1065_/A _1065_/B _1065_/C _1065_/Y VGND VGND VPWR VPWR _1065_/Y sky130_fd_sc_hd__nor4_1
XFILLER_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0918_ _0949_/A VGND VGND VPWR VPWR io_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_105_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0849_ VGND VGND VPWR VPWR _0849_/HI _1138_/C sky130_fd_sc_hd__conb_1
XFILLER_88_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_0_0_stoch_adc_comp.clk clkbuf_2_0_0_stoch_adc_comp.clk/X VGND VGND VPWR
+ VPWR _1030_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0703_ VGND VGND VPWR VPWR _0703_/HI _1080_/A sky130_fd_sc_hd__conb_1
XFILLER_8_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0634_ VGND VGND VPWR VPWR _0634_/HI _1052_/C sky130_fd_sc_hd__conb_1
XFILLER_48_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0565_ VGND VGND VPWR VPWR _0565_/HI la_data_out[73] sky130_fd_sc_hd__conb_1
XFILLER_112_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0496_ VGND VGND VPWR VPWR _0496_/HI _1166_/C sky130_fd_sc_hd__conb_1
XFILLER_100_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_285_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_stoch_adc_comp.clk clkbuf_3_2_0_stoch_adc_comp.clk/A VGND VGND VPWR
+ VPWR _1013_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_226_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1117_ _1117_/A _1117_/B _1117_/C _1117_/Y VGND VGND VPWR VPWR _1117_/Y sky130_fd_sc_hd__nor4_1
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1048_ _1048_/A analog_io[25] _1048_/C _1048_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_277_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_stoch_adc_comp.clk clkbuf_3_5_0_stoch_adc_comp.clk/A VGND VGND VPWR
+ VPWR _1003_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_153_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0617_ VGND VGND VPWR VPWR _0617_/HI la_data_out[125] sky130_fd_sc_hd__conb_1
XFILLER_113_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0548_ VGND VGND VPWR VPWR _0548_/HI la_data_out[56] sky130_fd_sc_hd__conb_1
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0479_ wbs_dat_o[7] _0478_/X io_out[7] _0473_/X VGND VGND VPWR VPWR _1021_/D sky130_fd_sc_hd__o22a_4
XFILLER_41_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_stoch_adc_comp.clk clkbuf_2_3_0_stoch_adc_comp.clk/X VGND VGND VPWR
+ VPWR _1005_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_283_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0951_ io_out[1] VGND VGND VPWR VPWR la_data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_105_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0882_ VGND VGND VPWR VPWR _0882_/HI _1151_/D sky130_fd_sc_hd__conb_1
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_stoch_adc_comp.clk clkbuf_2_1_0_stoch_adc_comp.clk/A VGND VGND VPWR
+ VPWR clkbuf_3_2_0_stoch_adc_comp.clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_266_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1150_ _1149_/D _1150_/B _1150_/C _1149_/A VGND VGND VPWR VPWR _1149_/A sky130_fd_sc_hd__nor4_1
XFILLER_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1081_ _1081_/A _1081_/B _1081_/C _1081_/Y VGND VGND VPWR VPWR _1081_/Y sky130_fd_sc_hd__nor4_1
XFILLER_59_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0934_ _0949_/A VGND VGND VPWR VPWR io_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_14_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0865_ VGND VGND VPWR VPWR _0865_/HI _1144_/D sky130_fd_sc_hd__conb_1
XFILLER_228_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0796_ VGND VGND VPWR VPWR _0796_/HI _1117_/B sky130_fd_sc_hd__conb_1
XFILLER_115_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_stoch_adc_comp.clk clkbuf_2_3_0_stoch_adc_comp.clk/A VGND VGND VPWR
+ VPWR clkbuf_2_3_0_stoch_adc_comp.clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_279_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0650_ VGND VGND VPWR VPWR _0650_/HI _1059_/A sky130_fd_sc_hd__conb_1
XFILLER_13_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0581_ VGND VGND VPWR VPWR _0581_/HI la_data_out[89] sky130_fd_sc_hd__conb_1
XFILLER_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1133_ _1133_/A _1133_/B _1133_/C _1133_/Y VGND VGND VPWR VPWR _1133_/Y sky130_fd_sc_hd__nor4_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1064_ _1064_/A analog_io[25] _1064_/C _1064_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_19_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0917_ _0949_/A VGND VGND VPWR VPWR io_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_175_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0848_ VGND VGND VPWR VPWR _0848_/HI _1138_/B sky130_fd_sc_hd__conb_1
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0779_ VGND VGND VPWR VPWR _0779_/HI _1110_/C sky130_fd_sc_hd__conb_1
XFILLER_115_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0702_ VGND VGND VPWR VPWR _0702_/HI _1079_/D sky130_fd_sc_hd__conb_1
XFILLER_239_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0633_ VGND VGND VPWR VPWR _0633_/HI _1052_/A sky130_fd_sc_hd__conb_1
XFILLER_48_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0564_ VGND VGND VPWR VPWR _0564_/HI la_data_out[72] sky130_fd_sc_hd__conb_1
XFILLER_135_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0495_ VGND VGND VPWR VPWR _0495_/HI _1166_/B sky130_fd_sc_hd__conb_1
XFILLER_61_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1116_ _1116_/A analog_io[25] _1116_/C _1116_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_81_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1047_ _1047_/A analog_io[24] _1047_/C _1047_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_250_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_253_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_stoch_adc_comp.clk clkbuf_0_stoch_adc_comp.clk/X VGND VGND VPWR VPWR
+ clkbuf_2_1_0_stoch_adc_comp.clk/A sky130_fd_sc_hd__clkbuf_1
XPHY_6870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0616_ VGND VGND VPWR VPWR _0616_/HI la_data_out[124] sky130_fd_sc_hd__conb_1
XFILLER_160_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0547_ VGND VGND VPWR VPWR _0547_/HI la_data_out[55] sky130_fd_sc_hd__conb_1
XFILLER_86_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0478_ _0464_/A VGND VGND VPWR VPWR _0478_/X sky130_fd_sc_hd__buf_2
XFILLER_67_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_260_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0950_ io_out[0] VGND VGND VPWR VPWR la_data_out[0] sky130_fd_sc_hd__buf_2
XPHY_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0881_ VGND VGND VPWR VPWR _0881_/HI _1151_/C sky130_fd_sc_hd__conb_1
XFILLER_174_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1080_ _1080_/A analog_io[25] _1080_/C _1080_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_225_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0933_ _0949_/A VGND VGND VPWR VPWR io_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0864_ VGND VGND VPWR VPWR _0864_/HI _1144_/C sky130_fd_sc_hd__conb_1
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0795_ VGND VGND VPWR VPWR _0795_/HI _1116_/D sky130_fd_sc_hd__conb_1
XFILLER_157_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0580_ VGND VGND VPWR VPWR _0580_/HI la_data_out[88] sky130_fd_sc_hd__conb_1
XFILLER_152_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1132_ _1132_/A analog_io[25] _1132_/C _1132_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_281_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1063_ _1063_/A analog_io[24] _1063_/C _1063_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0916_ _0949_/A VGND VGND VPWR VPWR io_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_179_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0847_ VGND VGND VPWR VPWR _0847_/HI _1137_/C sky130_fd_sc_hd__conb_1
XFILLER_192_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0778_ VGND VGND VPWR VPWR _0778_/HI _1110_/B sky130_fd_sc_hd__conb_1
XFILLER_66_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_281_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0701_ VGND VGND VPWR VPWR _0701_/HI _1079_/C sky130_fd_sc_hd__conb_1
XFILLER_117_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0632_ VGND VGND VPWR VPWR _0632_/HI _1051_/D sky130_fd_sc_hd__conb_1
XFILLER_67_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0563_ VGND VGND VPWR VPWR _0563_/HI la_data_out[71] sky130_fd_sc_hd__conb_1
XFILLER_48_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0494_ VGND VGND VPWR VPWR _0494_/HI _1165_/C sky130_fd_sc_hd__conb_1
XFILLER_112_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1115_ _1115_/A analog_io[24] _1115_/C _1115_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_54_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1046_ _1030_/CLK _0442_/X VGND VGND VPWR VPWR wbs_ack_o sky130_fd_sc_hd__dfxtp_4
XFILLER_74_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0615_ VGND VGND VPWR VPWR _0615_/HI la_data_out[123] sky130_fd_sc_hd__conb_1
XFILLER_158_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0546_ VGND VGND VPWR VPWR _0546_/HI la_data_out[54] sky130_fd_sc_hd__conb_1
XFILLER_258_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0477_ wbs_dat_o[8] _0471_/X io_out[8] _0473_/X VGND VGND VPWR VPWR _0477_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1029_ _1030_/CLK _1029_/D VGND VGND VPWR VPWR wbs_dat_o[15] sky130_fd_sc_hd__dfxtp_4
XFILLER_74_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_253_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0529_ VGND VGND VPWR VPWR _0529_/HI la_data_out[37] sky130_fd_sc_hd__conb_1
XFILLER_100_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_254_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0880_ VGND VGND VPWR VPWR _0880_/HI _1151_/A sky130_fd_sc_hd__conb_1
XFILLER_146_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0932_ _0949_/A VGND VGND VPWR VPWR io_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_140_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0863_ VGND VGND VPWR VPWR _0863_/HI _1144_/A sky130_fd_sc_hd__conb_1
XFILLER_146_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0794_ VGND VGND VPWR VPWR _0794_/HI _1116_/C sky130_fd_sc_hd__conb_1
XFILLER_127_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_266_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_249_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1131_ _1131_/A analog_io[24] _1131_/C _1131_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_226_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1062_ _1061_/Y _1062_/B _1062_/C _1061_/A VGND VGND VPWR VPWR _1061_/A sky130_fd_sc_hd__nor4_1
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0915_ _0949_/A VGND VGND VPWR VPWR io_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_147_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0846_ VGND VGND VPWR VPWR _0846_/HI _1137_/B sky130_fd_sc_hd__conb_1
XFILLER_105_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0777_ VGND VGND VPWR VPWR _0777_/HI _1109_/C sky130_fd_sc_hd__conb_1
XFILLER_161_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_279_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0700_ VGND VGND VPWR VPWR _0700_/HI _1079_/A sky130_fd_sc_hd__conb_1
XFILLER_209_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0631_ VGND VGND VPWR VPWR _0631_/HI _1051_/C sky130_fd_sc_hd__conb_1
XFILLER_125_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0562_ VGND VGND VPWR VPWR _0562_/HI la_data_out[70] sky130_fd_sc_hd__conb_1
XFILLER_256_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0493_ VGND VGND VPWR VPWR _0493_/HI _1165_/B sky130_fd_sc_hd__conb_1
XFILLER_239_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1114_ _1113_/Y _1114_/B _1114_/C _1114_/Y VGND VGND VPWR VPWR _1114_/Y sky130_fd_sc_hd__nor4_1
XFILLER_285_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1045_ _0989_/CLK _0445_/X VGND VGND VPWR VPWR wbs_dat_o[31] sky130_fd_sc_hd__dfxtp_4
XFILLER_94_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0829_ VGND VGND VPWR VPWR _0829_/HI _1130_/C sky130_fd_sc_hd__conb_1
XFILLER_128_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0614_ VGND VGND VPWR VPWR _0614_/HI la_data_out[122] sky130_fd_sc_hd__conb_1
XFILLER_217_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0545_ VGND VGND VPWR VPWR _0545_/HI la_data_out[53] sky130_fd_sc_hd__conb_1
XFILLER_98_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0476_ wbs_dat_o[9] _0471_/X io_out[9] _0473_/X VGND VGND VPWR VPWR _1023_/D sky130_fd_sc_hd__o22a_4
XFILLER_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1028_ _1030_/CLK _1028_/D VGND VGND VPWR VPWR wbs_dat_o[14] sky130_fd_sc_hd__dfxtp_4
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_283_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_282_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0528_ VGND VGND VPWR VPWR _0528_/HI la_data_out[36] sky130_fd_sc_hd__conb_1
XFILLER_247_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0459_ _0459_/A VGND VGND VPWR VPWR _0459_/X sky130_fd_sc_hd__buf_2
XFILLER_39_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_273_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_254_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_270_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_274_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_278_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ _0949_/A VGND VGND VPWR VPWR io_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_187_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0862_ VGND VGND VPWR VPWR _0862_/HI _1143_/D sky130_fd_sc_hd__conb_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0793_ VGND VGND VPWR VPWR _0793_/HI _1116_/A sky130_fd_sc_hd__conb_1
XFILLER_31_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1130_ _1129_/Y _1130_/B _1130_/C _1129_/A VGND VGND VPWR VPWR _1129_/A sky130_fd_sc_hd__nor4_1
XFILLER_66_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1061_ _1061_/A _1061_/B _1061_/C _1061_/Y VGND VGND VPWR VPWR _1061_/Y sky130_fd_sc_hd__nor4_1
XFILLER_81_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0914_ _0949_/A VGND VGND VPWR VPWR io_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_239_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0845_ VGND VGND VPWR VPWR _0845_/HI _1136_/D sky130_fd_sc_hd__conb_1
XFILLER_175_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0776_ VGND VGND VPWR VPWR _0776_/HI _1109_/B sky130_fd_sc_hd__conb_1
XFILLER_196_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0630_ VGND VGND VPWR VPWR _0630_/HI _1051_/A sky130_fd_sc_hd__conb_1
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0561_ VGND VGND VPWR VPWR _0561_/HI la_data_out[69] sky130_fd_sc_hd__conb_1
XFILLER_174_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0492_ VGND VGND VPWR VPWR _0492_/HI _1164_/D sky130_fd_sc_hd__conb_1
XFILLER_139_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1113_ _1114_/Y _1113_/B _1113_/C _1113_/Y VGND VGND VPWR VPWR _1113_/Y sky130_fd_sc_hd__nor4_1
XFILLER_66_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1044_ _0989_/CLK _1044_/D VGND VGND VPWR VPWR wbs_dat_o[30] sky130_fd_sc_hd__dfxtp_4
XFILLER_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0828_ VGND VGND VPWR VPWR _0828_/HI _1130_/B sky130_fd_sc_hd__conb_1
XFILLER_200_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0759_ VGND VGND VPWR VPWR _0759_/HI _1102_/C sky130_fd_sc_hd__conb_1
XFILLER_116_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0613_ VGND VGND VPWR VPWR _0613_/HI la_data_out[121] sky130_fd_sc_hd__conb_1
XFILLER_119_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0544_ VGND VGND VPWR VPWR _0544_/HI la_data_out[52] sky130_fd_sc_hd__conb_1
XFILLER_67_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0475_ wbs_dat_o[10] _0471_/X io_out[10] _0473_/X VGND VGND VPWR VPWR _0475_/X sky130_fd_sc_hd__o22a_4
XFILLER_234_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1027_ _1035_/CLK _1027_/D VGND VGND VPWR VPWR wbs_dat_o[13] sky130_fd_sc_hd__dfxtp_4
XFILLER_223_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0527_ VGND VGND VPWR VPWR _0527_/HI la_data_out[35] sky130_fd_sc_hd__conb_1
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0458_ wbs_dat_o[22] _0457_/X io_out[22] _0452_/X VGND VGND VPWR VPWR _1036_/D sky130_fd_sc_hd__o22a_4
XFILLER_255_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0930_ _0949_/A VGND VGND VPWR VPWR io_oeb[17] sky130_fd_sc_hd__buf_2
XPHY_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0861_ VGND VGND VPWR VPWR _0861_/HI _1143_/C sky130_fd_sc_hd__conb_1
XFILLER_158_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0792_ VGND VGND VPWR VPWR _0792_/HI _1115_/D sky130_fd_sc_hd__conb_1
XFILLER_173_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1060_ _1060_/A analog_io[25] _1060_/C _1060_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_248_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0913_ _0949_/A VGND VGND VPWR VPWR io_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_163_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0844_ VGND VGND VPWR VPWR _0844_/HI _1136_/C sky130_fd_sc_hd__conb_1
XFILLER_179_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0775_ VGND VGND VPWR VPWR _0775_/HI _1108_/D sky130_fd_sc_hd__conb_1
XFILLER_255_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0560_ VGND VGND VPWR VPWR _0560_/HI la_data_out[68] sky130_fd_sc_hd__conb_1
XFILLER_217_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0491_ VGND VGND VPWR VPWR _0491_/HI _1164_/C sky130_fd_sc_hd__conb_1
XFILLER_225_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1112_ _1112_/A analog_io[25] _1112_/C _1112_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_238_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1043_ _0989_/CLK _0447_/X VGND VGND VPWR VPWR wbs_dat_o[29] sky130_fd_sc_hd__dfxtp_4
XFILLER_235_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0827_ VGND VGND VPWR VPWR _0827_/HI _1129_/C sky130_fd_sc_hd__conb_1
XFILLER_134_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0758_ VGND VGND VPWR VPWR _0758_/HI _1102_/B sky130_fd_sc_hd__conb_1
XFILLER_115_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0689_ VGND VGND VPWR VPWR _0689_/HI _1074_/C sky130_fd_sc_hd__conb_1
XFILLER_103_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0612_ VGND VGND VPWR VPWR _0612_/HI la_data_out[120] sky130_fd_sc_hd__conb_1
XFILLER_119_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0543_ VGND VGND VPWR VPWR _0543_/HI la_data_out[51] sky130_fd_sc_hd__conb_1
XFILLER_112_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0474_ wbs_dat_o[11] _0471_/X io_out[11] _0473_/X VGND VGND VPWR VPWR _1025_/D sky130_fd_sc_hd__o22a_4
XFILLER_100_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1026_ _1030_/CLK _1026_/D VGND VGND VPWR VPWR wbs_dat_o[12] sky130_fd_sc_hd__dfxtp_4
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_0 io_out[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_275_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0526_ VGND VGND VPWR VPWR _0526_/HI la_data_out[34] sky130_fd_sc_hd__conb_1
XFILLER_45_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0457_ _0449_/X VGND VGND VPWR VPWR _0457_/X sky130_fd_sc_hd__buf_2
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1009_ _1013_/CLK _1065_/A VGND VGND VPWR VPWR io_out[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_274_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_284_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0509_ VGND VGND VPWR VPWR _0509_/HI _1171_/D sky130_fd_sc_hd__conb_1
XFILLER_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0860_ VGND VGND VPWR VPWR _0860_/HI _1143_/A sky130_fd_sc_hd__conb_1
XFILLER_144_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0791_ VGND VGND VPWR VPWR _0791_/HI _1115_/C sky130_fd_sc_hd__conb_1
XFILLER_70_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_272_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0989_ _0989_/CLK _1145_/A VGND VGND VPWR VPWR io_out[24] sky130_fd_sc_hd__dfxtp_4
XFILLER_285_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0912_ VGND VGND VPWR VPWR _0912_/HI _1163_/D sky130_fd_sc_hd__conb_1
XFILLER_222_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0843_ VGND VGND VPWR VPWR _0843_/HI _1136_/A sky130_fd_sc_hd__conb_1
XFILLER_35_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0774_ VGND VGND VPWR VPWR _0774_/HI _1108_/C sky130_fd_sc_hd__conb_1
XFILLER_259_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0490_ VGND VGND VPWR VPWR _0490_/HI _1164_/A sky130_fd_sc_hd__conb_1
XFILLER_140_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1111_ _1111_/A analog_io[24] _1111_/C _1111_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_152_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1042_ _0989_/CLK _0448_/X VGND VGND VPWR VPWR wbs_dat_o[28] sky130_fd_sc_hd__dfxtp_4
XFILLER_59_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0826_ VGND VGND VPWR VPWR _0826_/HI _1129_/B sky130_fd_sc_hd__conb_1
XFILLER_116_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0757_ VGND VGND VPWR VPWR _0757_/HI _1101_/C sky130_fd_sc_hd__conb_1
XFILLER_239_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0688_ VGND VGND VPWR VPWR _0688_/HI _1074_/B sky130_fd_sc_hd__conb_1
XFILLER_83_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0611_ VGND VGND VPWR VPWR _0611_/HI la_data_out[119] sky130_fd_sc_hd__conb_1
XFILLER_256_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0542_ VGND VGND VPWR VPWR _0542_/HI la_data_out[50] sky130_fd_sc_hd__conb_1
XFILLER_4_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0473_ _0466_/A VGND VGND VPWR VPWR _0473_/X sky130_fd_sc_hd__buf_2
XFILLER_61_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_252_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1025_ _1030_/CLK _1025_/D VGND VGND VPWR VPWR wbs_dat_o[11] sky130_fd_sc_hd__dfxtp_4
XFILLER_267_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0809_ VGND VGND VPWR VPWR _0809_/HI _1122_/C sky130_fd_sc_hd__conb_1
XFILLER_176_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_1 io_out[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0525_ VGND VGND VPWR VPWR _0525_/HI la_data_out[33] sky130_fd_sc_hd__conb_1
XFILLER_99_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0456_ wbs_dat_o[23] _0450_/X io_out[23] _0452_/X VGND VGND VPWR VPWR _1037_/D sky130_fd_sc_hd__o22a_4
XFILLER_67_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1008_ _1013_/CLK _1069_/A VGND VGND VPWR VPWR io_out[5] sky130_fd_sc_hd__dfxtp_4
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0508_ VGND VGND VPWR VPWR _0508_/HI _1171_/C sky130_fd_sc_hd__conb_1
XFILLER_236_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0439_ la_data_in[67] la_oen[67] wb_rst_i _0438_/Y VGND VGND VPWR VPWR _0949_/A sky130_fd_sc_hd__o22a_4
XFILLER_67_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0790_ VGND VGND VPWR VPWR _0790_/HI _1115_/A sky130_fd_sc_hd__conb_1
XFILLER_220_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0988_ _0987_/CLK _1149_/A VGND VGND VPWR VPWR io_out[25] sky130_fd_sc_hd__dfxtp_4
XFILLER_14_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_249_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0911_ VGND VGND VPWR VPWR _0911_/HI _1163_/C sky130_fd_sc_hd__conb_1
XFILLER_239_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0842_ VGND VGND VPWR VPWR _0842_/HI _1135_/D sky130_fd_sc_hd__conb_1
XFILLER_31_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0773_ VGND VGND VPWR VPWR _0773_/HI _1108_/A sky130_fd_sc_hd__conb_1
XFILLER_128_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_252_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_284_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_273_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1110_ _1110_/A _1110_/B _1110_/C _1110_/Y VGND VGND VPWR VPWR _1110_/Y sky130_fd_sc_hd__nor4_1
XFILLER_43_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1041_ _1003_/CLK _1041_/D VGND VGND VPWR VPWR wbs_dat_o[27] sky130_fd_sc_hd__dfxtp_4
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0825_ VGND VGND VPWR VPWR _0825_/HI _1128_/D sky130_fd_sc_hd__conb_1
XFILLER_198_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0756_ VGND VGND VPWR VPWR _0756_/HI _1101_/B sky130_fd_sc_hd__conb_1
XFILLER_66_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0687_ VGND VGND VPWR VPWR _0687_/HI _1073_/C sky130_fd_sc_hd__conb_1
XFILLER_170_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_281_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_279_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0610_ VGND VGND VPWR VPWR _0610_/HI la_data_out[118] sky130_fd_sc_hd__conb_1
XFILLER_109_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0541_ VGND VGND VPWR VPWR _0541_/HI la_data_out[49] sky130_fd_sc_hd__conb_1
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0472_ wbs_dat_o[12] _0471_/X io_out[12] _0466_/X VGND VGND VPWR VPWR _1026_/D sky130_fd_sc_hd__o22a_4
XFILLER_65_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1024_ _1030_/CLK _0475_/X VGND VGND VPWR VPWR wbs_dat_o[10] sky130_fd_sc_hd__dfxtp_4
XFILLER_19_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0808_ VGND VGND VPWR VPWR _0808_/HI _1122_/B sky130_fd_sc_hd__conb_1
XFILLER_89_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0739_ VGND VGND VPWR VPWR _0739_/HI _1094_/C sky130_fd_sc_hd__conb_1
XFILLER_274_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_2 io_out[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0524_ VGND VGND VPWR VPWR _0524_/HI la_data_out[32] sky130_fd_sc_hd__conb_1
XFILLER_99_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0455_ wbs_dat_o[24] _0450_/X io_out[24] _0452_/X VGND VGND VPWR VPWR _0455_/X sky130_fd_sc_hd__o22a_4
XFILLER_112_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1007_ _1013_/CLK _1073_/A VGND VGND VPWR VPWR io_out[6] sky130_fd_sc_hd__dfxtp_4
XFILLER_165_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0507_ VGND VGND VPWR VPWR _0507_/HI _1171_/A sky130_fd_sc_hd__conb_1
XFILLER_28_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0438_ la_oen[67] VGND VGND VPWR VPWR _0438_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0987_ _0987_/CLK _1153_/A VGND VGND VPWR VPWR io_out[26] sky130_fd_sc_hd__dfxtp_4
XFILLER_160_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0910_ VGND VGND VPWR VPWR _0910_/HI _1163_/A sky130_fd_sc_hd__conb_1
XPHY_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0841_ VGND VGND VPWR VPWR _0841_/HI _1135_/C sky130_fd_sc_hd__conb_1
XFILLER_146_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0772_ VGND VGND VPWR VPWR _0772_/HI _1107_/D sky130_fd_sc_hd__conb_1
XFILLER_31_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1040_ _1003_/CLK _1040_/D VGND VGND VPWR VPWR wbs_dat_o[26] sky130_fd_sc_hd__dfxtp_4
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0824_ VGND VGND VPWR VPWR _0824_/HI _1128_/C sky130_fd_sc_hd__conb_1
XFILLER_70_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0755_ VGND VGND VPWR VPWR _0755_/HI _1100_/D sky130_fd_sc_hd__conb_1
XFILLER_274_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0686_ VGND VGND VPWR VPWR _0686_/HI _1073_/B sky130_fd_sc_hd__conb_1
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1169_ _1169_/A _1169_/B _1169_/C _1169_/Y VGND VGND VPWR VPWR _1169_/Y sky130_fd_sc_hd__nor4_1
XFILLER_168_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0540_ VGND VGND VPWR VPWR _0540_/HI la_data_out[48] sky130_fd_sc_hd__conb_1
XFILLER_256_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0471_ _0464_/A VGND VGND VPWR VPWR _0471_/X sky130_fd_sc_hd__buf_2
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_278_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1023_ _1035_/CLK _1023_/D VGND VGND VPWR VPWR wbs_dat_o[9] sky130_fd_sc_hd__dfxtp_4
XFILLER_78_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0807_ VGND VGND VPWR VPWR _0807_/HI _1121_/C sky130_fd_sc_hd__conb_1
XFILLER_200_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0738_ VGND VGND VPWR VPWR _0738_/HI _1094_/B sky130_fd_sc_hd__conb_1
XFILLER_226_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_274_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0669_ VGND VGND VPWR VPWR _0669_/HI _1066_/C sky130_fd_sc_hd__conb_1
XFILLER_226_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_3 io_out[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0523_ VGND VGND VPWR VPWR _0523_/HI io_out[37] sky130_fd_sc_hd__conb_1
XFILLER_140_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0454_ wbs_dat_o[25] _0450_/X io_out[25] _0452_/X VGND VGND VPWR VPWR _1039_/D sky130_fd_sc_hd__o22a_4
XFILLER_239_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1006_ _1006_/CLK _1077_/A VGND VGND VPWR VPWR io_out[7] sky130_fd_sc_hd__dfxtp_4
XFILLER_78_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0506_ VGND VGND VPWR VPWR _0506_/HI _1170_/C sky130_fd_sc_hd__conb_1
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0437_ wbs_cyc_i VGND VGND VPWR VPWR _0437_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0986_ _0987_/CLK _1157_/A VGND VGND VPWR VPWR io_out[27] sky130_fd_sc_hd__dfxtp_4
XFILLER_203_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0840_ VGND VGND VPWR VPWR _0840_/HI _1135_/A sky130_fd_sc_hd__conb_1
XFILLER_204_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0771_ VGND VGND VPWR VPWR _0771_/HI _1107_/C sky130_fd_sc_hd__conb_1
XFILLER_31_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0969_ io_out[19] VGND VGND VPWR VPWR la_data_out[19] sky130_fd_sc_hd__buf_2
XFILLER_203_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_267_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0823_ VGND VGND VPWR VPWR _0823_/HI _1128_/A sky130_fd_sc_hd__conb_1
XFILLER_204_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0754_ VGND VGND VPWR VPWR _0754_/HI _1100_/C sky130_fd_sc_hd__conb_1
XFILLER_190_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0685_ VGND VGND VPWR VPWR _0685_/HI _1072_/D sky130_fd_sc_hd__conb_1
XFILLER_131_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1168_ _1168_/A analog_io[25] _1168_/C _1168_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1099_ _1099_/A analog_io[24] _1099_/C _1099_/D VGND VGND VPWR VPWR _1164_/Y sky130_fd_sc_hd__nor4_1
XFILLER_164_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0470_ wbs_dat_o[13] _0464_/X io_out[13] _0466_/X VGND VGND VPWR VPWR _1027_/D sky130_fd_sc_hd__o22a_4
XFILLER_79_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1022_ _1035_/CLK _0477_/X VGND VGND VPWR VPWR wbs_dat_o[8] sky130_fd_sc_hd__dfxtp_4
XFILLER_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0806_ VGND VGND VPWR VPWR _0806_/HI _1121_/B sky130_fd_sc_hd__conb_1
XFILLER_162_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0737_ VGND VGND VPWR VPWR _0737_/HI _1093_/C sky130_fd_sc_hd__conb_1
XFILLER_85_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0668_ VGND VGND VPWR VPWR _0668_/HI _1066_/B sky130_fd_sc_hd__conb_1
XFILLER_252_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0599_ VGND VGND VPWR VPWR _0599_/HI la_data_out[107] sky130_fd_sc_hd__conb_1
XFILLER_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_282_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_4 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0522_ VGND VGND VPWR VPWR _0522_/HI io_out[36] sky130_fd_sc_hd__conb_1
XFILLER_275_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0453_ wbs_dat_o[26] _0450_/X io_out[26] _0452_/X VGND VGND VPWR VPWR _1040_/D sky130_fd_sc_hd__o22a_4
XFILLER_141_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1005_ _1005_/CLK _1081_/A VGND VGND VPWR VPWR io_out[8] sky130_fd_sc_hd__dfxtp_4
XFILLER_228_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0505_ VGND VGND VPWR VPWR _0505_/HI _1170_/B sky130_fd_sc_hd__conb_1
XFILLER_87_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0436_ wbs_stb_i VGND VGND VPWR VPWR _0436_/Y sky130_fd_sc_hd__inv_2
.ends

