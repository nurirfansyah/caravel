magic
tech sky130A
magscale 1 2
timestamp 1608062367
<< obsli1 >>
rect 1104 2159 278852 237745
<< obsm1 >>
rect 1104 1368 278852 237776
<< metal2 >>
rect 1122 239200 1178 240000
rect 3422 239200 3478 240000
rect 5722 239200 5778 240000
rect 8022 239200 8078 240000
rect 10322 239200 10378 240000
rect 12622 239200 12678 240000
rect 14922 239200 14978 240000
rect 17314 239200 17370 240000
rect 19614 239200 19670 240000
rect 21914 239200 21970 240000
rect 24214 239200 24270 240000
rect 26514 239200 26570 240000
rect 28814 239200 28870 240000
rect 31114 239200 31170 240000
rect 33506 239200 33562 240000
rect 35806 239200 35862 240000
rect 38106 239200 38162 240000
rect 40406 239200 40462 240000
rect 42706 239200 42762 240000
rect 45006 239200 45062 240000
rect 47306 239200 47362 240000
rect 49698 239200 49754 240000
rect 51998 239200 52054 240000
rect 54298 239200 54354 240000
rect 56598 239200 56654 240000
rect 58898 239200 58954 240000
rect 61198 239200 61254 240000
rect 63590 239200 63646 240000
rect 65890 239200 65946 240000
rect 68190 239200 68246 240000
rect 70490 239200 70546 240000
rect 72790 239200 72846 240000
rect 75090 239200 75146 240000
rect 77390 239200 77446 240000
rect 79782 239200 79838 240000
rect 82082 239200 82138 240000
rect 84382 239200 84438 240000
rect 86682 239200 86738 240000
rect 88982 239200 89038 240000
rect 91282 239200 91338 240000
rect 93582 239200 93638 240000
rect 95974 239200 96030 240000
rect 98274 239200 98330 240000
rect 100574 239200 100630 240000
rect 102874 239200 102930 240000
rect 105174 239200 105230 240000
rect 107474 239200 107530 240000
rect 109774 239200 109830 240000
rect 112166 239200 112222 240000
rect 114466 239200 114522 240000
rect 116766 239200 116822 240000
rect 119066 239200 119122 240000
rect 121366 239200 121422 240000
rect 123666 239200 123722 240000
rect 126058 239200 126114 240000
rect 128358 239200 128414 240000
rect 130658 239200 130714 240000
rect 132958 239200 133014 240000
rect 135258 239200 135314 240000
rect 137558 239200 137614 240000
rect 139858 239200 139914 240000
rect 142250 239200 142306 240000
rect 144550 239200 144606 240000
rect 146850 239200 146906 240000
rect 149150 239200 149206 240000
rect 151450 239200 151506 240000
rect 153750 239200 153806 240000
rect 156050 239200 156106 240000
rect 158442 239200 158498 240000
rect 160742 239200 160798 240000
rect 163042 239200 163098 240000
rect 165342 239200 165398 240000
rect 167642 239200 167698 240000
rect 169942 239200 169998 240000
rect 172334 239200 172390 240000
rect 174634 239200 174690 240000
rect 176934 239200 176990 240000
rect 179234 239200 179290 240000
rect 181534 239200 181590 240000
rect 183834 239200 183890 240000
rect 186134 239200 186190 240000
rect 188526 239200 188582 240000
rect 190826 239200 190882 240000
rect 193126 239200 193182 240000
rect 195426 239200 195482 240000
rect 197726 239200 197782 240000
rect 200026 239200 200082 240000
rect 202326 239200 202382 240000
rect 204718 239200 204774 240000
rect 207018 239200 207074 240000
rect 209318 239200 209374 240000
rect 211618 239200 211674 240000
rect 213918 239200 213974 240000
rect 216218 239200 216274 240000
rect 218518 239200 218574 240000
rect 220910 239200 220966 240000
rect 223210 239200 223266 240000
rect 225510 239200 225566 240000
rect 227810 239200 227866 240000
rect 230110 239200 230166 240000
rect 232410 239200 232466 240000
rect 234802 239200 234858 240000
rect 237102 239200 237158 240000
rect 239402 239200 239458 240000
rect 241702 239200 241758 240000
rect 244002 239200 244058 240000
rect 246302 239200 246358 240000
rect 248602 239200 248658 240000
rect 250994 239200 251050 240000
rect 253294 239200 253350 240000
rect 255594 239200 255650 240000
rect 257894 239200 257950 240000
rect 260194 239200 260250 240000
rect 262494 239200 262550 240000
rect 264794 239200 264850 240000
rect 267186 239200 267242 240000
rect 269486 239200 269542 240000
rect 271786 239200 271842 240000
rect 274086 239200 274142 240000
rect 276386 239200 276442 240000
rect 278686 239200 278742 240000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8758 0 8814 800
rect 9310 0 9366 800
rect 9862 0 9918 800
rect 10414 0 10470 800
rect 10966 0 11022 800
rect 11518 0 11574 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13266 0 13322 800
rect 13818 0 13874 800
rect 14370 0 14426 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 16026 0 16082 800
rect 16578 0 16634 800
rect 17222 0 17278 800
rect 17774 0 17830 800
rect 18326 0 18382 800
rect 18878 0 18934 800
rect 19430 0 19486 800
rect 19982 0 20038 800
rect 20534 0 20590 800
rect 21086 0 21142 800
rect 21730 0 21786 800
rect 22282 0 22338 800
rect 22834 0 22890 800
rect 23386 0 23442 800
rect 23938 0 23994 800
rect 24490 0 24546 800
rect 25042 0 25098 800
rect 25686 0 25742 800
rect 26238 0 26294 800
rect 26790 0 26846 800
rect 27342 0 27398 800
rect 27894 0 27950 800
rect 28446 0 28502 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30194 0 30250 800
rect 30746 0 30802 800
rect 31298 0 31354 800
rect 31850 0 31906 800
rect 32402 0 32458 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36358 0 36414 800
rect 36910 0 36966 800
rect 37462 0 37518 800
rect 38106 0 38162 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39762 0 39818 800
rect 40314 0 40370 800
rect 40866 0 40922 800
rect 41418 0 41474 800
rect 41970 0 42026 800
rect 42614 0 42670 800
rect 43166 0 43222 800
rect 43718 0 43774 800
rect 44270 0 44326 800
rect 44822 0 44878 800
rect 45374 0 45430 800
rect 45926 0 45982 800
rect 46570 0 46626 800
rect 47122 0 47178 800
rect 47674 0 47730 800
rect 48226 0 48282 800
rect 48778 0 48834 800
rect 49330 0 49386 800
rect 49882 0 49938 800
rect 50526 0 50582 800
rect 51078 0 51134 800
rect 51630 0 51686 800
rect 52182 0 52238 800
rect 52734 0 52790 800
rect 53286 0 53342 800
rect 53838 0 53894 800
rect 54390 0 54446 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58990 0 59046 800
rect 59542 0 59598 800
rect 60094 0 60150 800
rect 60646 0 60702 800
rect 61198 0 61254 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62854 0 62910 800
rect 63498 0 63554 800
rect 64050 0 64106 800
rect 64602 0 64658 800
rect 65154 0 65210 800
rect 65706 0 65762 800
rect 66258 0 66314 800
rect 66810 0 66866 800
rect 67454 0 67510 800
rect 68006 0 68062 800
rect 68558 0 68614 800
rect 69110 0 69166 800
rect 69662 0 69718 800
rect 70214 0 70270 800
rect 70766 0 70822 800
rect 71410 0 71466 800
rect 71962 0 72018 800
rect 72514 0 72570 800
rect 73066 0 73122 800
rect 73618 0 73674 800
rect 74170 0 74226 800
rect 74722 0 74778 800
rect 75274 0 75330 800
rect 75918 0 75974 800
rect 76470 0 76526 800
rect 77022 0 77078 800
rect 77574 0 77630 800
rect 78126 0 78182 800
rect 78678 0 78734 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 80426 0 80482 800
rect 80978 0 81034 800
rect 81530 0 81586 800
rect 82082 0 82138 800
rect 82634 0 82690 800
rect 83186 0 83242 800
rect 83738 0 83794 800
rect 84382 0 84438 800
rect 84934 0 84990 800
rect 85486 0 85542 800
rect 86038 0 86094 800
rect 86590 0 86646 800
rect 87142 0 87198 800
rect 87694 0 87750 800
rect 88338 0 88394 800
rect 88890 0 88946 800
rect 89442 0 89498 800
rect 89994 0 90050 800
rect 90546 0 90602 800
rect 91098 0 91154 800
rect 91650 0 91706 800
rect 92294 0 92350 800
rect 92846 0 92902 800
rect 93398 0 93454 800
rect 93950 0 94006 800
rect 94502 0 94558 800
rect 95054 0 95110 800
rect 95606 0 95662 800
rect 96158 0 96214 800
rect 96802 0 96858 800
rect 97354 0 97410 800
rect 97906 0 97962 800
rect 98458 0 98514 800
rect 99010 0 99066 800
rect 99562 0 99618 800
rect 100114 0 100170 800
rect 100758 0 100814 800
rect 101310 0 101366 800
rect 101862 0 101918 800
rect 102414 0 102470 800
rect 102966 0 103022 800
rect 103518 0 103574 800
rect 104070 0 104126 800
rect 104622 0 104678 800
rect 105266 0 105322 800
rect 105818 0 105874 800
rect 106370 0 106426 800
rect 106922 0 106978 800
rect 107474 0 107530 800
rect 108026 0 108082 800
rect 108578 0 108634 800
rect 109222 0 109278 800
rect 109774 0 109830 800
rect 110326 0 110382 800
rect 110878 0 110934 800
rect 111430 0 111486 800
rect 111982 0 112038 800
rect 112534 0 112590 800
rect 113178 0 113234 800
rect 113730 0 113786 800
rect 114282 0 114338 800
rect 114834 0 114890 800
rect 115386 0 115442 800
rect 115938 0 115994 800
rect 116490 0 116546 800
rect 117042 0 117098 800
rect 117686 0 117742 800
rect 118238 0 118294 800
rect 118790 0 118846 800
rect 119342 0 119398 800
rect 119894 0 119950 800
rect 120446 0 120502 800
rect 120998 0 121054 800
rect 121642 0 121698 800
rect 122194 0 122250 800
rect 122746 0 122802 800
rect 123298 0 123354 800
rect 123850 0 123906 800
rect 124402 0 124458 800
rect 124954 0 125010 800
rect 125506 0 125562 800
rect 126150 0 126206 800
rect 126702 0 126758 800
rect 127254 0 127310 800
rect 127806 0 127862 800
rect 128358 0 128414 800
rect 128910 0 128966 800
rect 129462 0 129518 800
rect 130106 0 130162 800
rect 130658 0 130714 800
rect 131210 0 131266 800
rect 131762 0 131818 800
rect 132314 0 132370 800
rect 132866 0 132922 800
rect 133418 0 133474 800
rect 134062 0 134118 800
rect 134614 0 134670 800
rect 135166 0 135222 800
rect 135718 0 135774 800
rect 136270 0 136326 800
rect 136822 0 136878 800
rect 137374 0 137430 800
rect 137926 0 137982 800
rect 138570 0 138626 800
rect 139122 0 139178 800
rect 139674 0 139730 800
rect 140226 0 140282 800
rect 140778 0 140834 800
rect 141330 0 141386 800
rect 141882 0 141938 800
rect 142526 0 142582 800
rect 143078 0 143134 800
rect 143630 0 143686 800
rect 144182 0 144238 800
rect 144734 0 144790 800
rect 145286 0 145342 800
rect 145838 0 145894 800
rect 146390 0 146446 800
rect 147034 0 147090 800
rect 147586 0 147642 800
rect 148138 0 148194 800
rect 148690 0 148746 800
rect 149242 0 149298 800
rect 149794 0 149850 800
rect 150346 0 150402 800
rect 150990 0 151046 800
rect 151542 0 151598 800
rect 152094 0 152150 800
rect 152646 0 152702 800
rect 153198 0 153254 800
rect 153750 0 153806 800
rect 154302 0 154358 800
rect 154946 0 155002 800
rect 155498 0 155554 800
rect 156050 0 156106 800
rect 156602 0 156658 800
rect 157154 0 157210 800
rect 157706 0 157762 800
rect 158258 0 158314 800
rect 158810 0 158866 800
rect 159454 0 159510 800
rect 160006 0 160062 800
rect 160558 0 160614 800
rect 161110 0 161166 800
rect 161662 0 161718 800
rect 162214 0 162270 800
rect 162766 0 162822 800
rect 163410 0 163466 800
rect 163962 0 164018 800
rect 164514 0 164570 800
rect 165066 0 165122 800
rect 165618 0 165674 800
rect 166170 0 166226 800
rect 166722 0 166778 800
rect 167274 0 167330 800
rect 167918 0 167974 800
rect 168470 0 168526 800
rect 169022 0 169078 800
rect 169574 0 169630 800
rect 170126 0 170182 800
rect 170678 0 170734 800
rect 171230 0 171286 800
rect 171874 0 171930 800
rect 172426 0 172482 800
rect 172978 0 173034 800
rect 173530 0 173586 800
rect 174082 0 174138 800
rect 174634 0 174690 800
rect 175186 0 175242 800
rect 175830 0 175886 800
rect 176382 0 176438 800
rect 176934 0 176990 800
rect 177486 0 177542 800
rect 178038 0 178094 800
rect 178590 0 178646 800
rect 179142 0 179198 800
rect 179694 0 179750 800
rect 180338 0 180394 800
rect 180890 0 180946 800
rect 181442 0 181498 800
rect 181994 0 182050 800
rect 182546 0 182602 800
rect 183098 0 183154 800
rect 183650 0 183706 800
rect 184294 0 184350 800
rect 184846 0 184902 800
rect 185398 0 185454 800
rect 185950 0 186006 800
rect 186502 0 186558 800
rect 187054 0 187110 800
rect 187606 0 187662 800
rect 188158 0 188214 800
rect 188802 0 188858 800
rect 189354 0 189410 800
rect 189906 0 189962 800
rect 190458 0 190514 800
rect 191010 0 191066 800
rect 191562 0 191618 800
rect 192114 0 192170 800
rect 192758 0 192814 800
rect 193310 0 193366 800
rect 193862 0 193918 800
rect 194414 0 194470 800
rect 194966 0 195022 800
rect 195518 0 195574 800
rect 196070 0 196126 800
rect 196714 0 196770 800
rect 197266 0 197322 800
rect 197818 0 197874 800
rect 198370 0 198426 800
rect 198922 0 198978 800
rect 199474 0 199530 800
rect 200026 0 200082 800
rect 200578 0 200634 800
rect 201222 0 201278 800
rect 201774 0 201830 800
rect 202326 0 202382 800
rect 202878 0 202934 800
rect 203430 0 203486 800
rect 203982 0 204038 800
rect 204534 0 204590 800
rect 205178 0 205234 800
rect 205730 0 205786 800
rect 206282 0 206338 800
rect 206834 0 206890 800
rect 207386 0 207442 800
rect 207938 0 207994 800
rect 208490 0 208546 800
rect 209042 0 209098 800
rect 209686 0 209742 800
rect 210238 0 210294 800
rect 210790 0 210846 800
rect 211342 0 211398 800
rect 211894 0 211950 800
rect 212446 0 212502 800
rect 212998 0 213054 800
rect 213642 0 213698 800
rect 214194 0 214250 800
rect 214746 0 214802 800
rect 215298 0 215354 800
rect 215850 0 215906 800
rect 216402 0 216458 800
rect 216954 0 217010 800
rect 217598 0 217654 800
rect 218150 0 218206 800
rect 218702 0 218758 800
rect 219254 0 219310 800
rect 219806 0 219862 800
rect 220358 0 220414 800
rect 220910 0 220966 800
rect 221462 0 221518 800
rect 222106 0 222162 800
rect 222658 0 222714 800
rect 223210 0 223266 800
rect 223762 0 223818 800
rect 224314 0 224370 800
rect 224866 0 224922 800
rect 225418 0 225474 800
rect 226062 0 226118 800
rect 226614 0 226670 800
rect 227166 0 227222 800
rect 227718 0 227774 800
rect 228270 0 228326 800
rect 228822 0 228878 800
rect 229374 0 229430 800
rect 229926 0 229982 800
rect 230570 0 230626 800
rect 231122 0 231178 800
rect 231674 0 231730 800
rect 232226 0 232282 800
rect 232778 0 232834 800
rect 233330 0 233386 800
rect 233882 0 233938 800
rect 234526 0 234582 800
rect 235078 0 235134 800
rect 235630 0 235686 800
rect 236182 0 236238 800
rect 236734 0 236790 800
rect 237286 0 237342 800
rect 237838 0 237894 800
rect 238482 0 238538 800
rect 239034 0 239090 800
rect 239586 0 239642 800
rect 240138 0 240194 800
rect 240690 0 240746 800
rect 241242 0 241298 800
rect 241794 0 241850 800
rect 242346 0 242402 800
rect 242990 0 243046 800
rect 243542 0 243598 800
rect 244094 0 244150 800
rect 244646 0 244702 800
rect 245198 0 245254 800
rect 245750 0 245806 800
rect 246302 0 246358 800
rect 246946 0 247002 800
rect 247498 0 247554 800
rect 248050 0 248106 800
rect 248602 0 248658 800
rect 249154 0 249210 800
rect 249706 0 249762 800
rect 250258 0 250314 800
rect 250810 0 250866 800
rect 251454 0 251510 800
rect 252006 0 252062 800
rect 252558 0 252614 800
rect 253110 0 253166 800
rect 253662 0 253718 800
rect 254214 0 254270 800
rect 254766 0 254822 800
rect 255410 0 255466 800
rect 255962 0 256018 800
rect 256514 0 256570 800
rect 257066 0 257122 800
rect 257618 0 257674 800
rect 258170 0 258226 800
rect 258722 0 258778 800
rect 259366 0 259422 800
rect 259918 0 259974 800
rect 260470 0 260526 800
rect 261022 0 261078 800
rect 261574 0 261630 800
rect 262126 0 262182 800
rect 262678 0 262734 800
rect 263230 0 263286 800
rect 263874 0 263930 800
rect 264426 0 264482 800
rect 264978 0 265034 800
rect 265530 0 265586 800
rect 266082 0 266138 800
rect 266634 0 266690 800
rect 267186 0 267242 800
rect 267830 0 267886 800
rect 268382 0 268438 800
rect 268934 0 268990 800
rect 269486 0 269542 800
rect 270038 0 270094 800
rect 270590 0 270646 800
rect 271142 0 271198 800
rect 271694 0 271750 800
rect 272338 0 272394 800
rect 272890 0 272946 800
rect 273442 0 273498 800
rect 273994 0 274050 800
rect 274546 0 274602 800
rect 275098 0 275154 800
rect 275650 0 275706 800
rect 276294 0 276350 800
rect 276846 0 276902 800
rect 277398 0 277454 800
rect 277950 0 278006 800
rect 278502 0 278558 800
rect 279054 0 279110 800
rect 279606 0 279662 800
<< obsm2 >>
rect 294 239144 1066 239200
rect 1234 239144 3366 239200
rect 3534 239144 5666 239200
rect 5834 239144 7966 239200
rect 8134 239144 10266 239200
rect 10434 239144 12566 239200
rect 12734 239144 14866 239200
rect 15034 239144 17258 239200
rect 17426 239144 19558 239200
rect 19726 239144 21858 239200
rect 22026 239144 24158 239200
rect 24326 239144 26458 239200
rect 26626 239144 28758 239200
rect 28926 239144 31058 239200
rect 31226 239144 33450 239200
rect 33618 239144 35750 239200
rect 35918 239144 38050 239200
rect 38218 239144 40350 239200
rect 40518 239144 42650 239200
rect 42818 239144 44950 239200
rect 45118 239144 47250 239200
rect 47418 239144 49642 239200
rect 49810 239144 51942 239200
rect 52110 239144 54242 239200
rect 54410 239144 56542 239200
rect 56710 239144 58842 239200
rect 59010 239144 61142 239200
rect 61310 239144 63534 239200
rect 63702 239144 65834 239200
rect 66002 239144 68134 239200
rect 68302 239144 70434 239200
rect 70602 239144 72734 239200
rect 72902 239144 75034 239200
rect 75202 239144 77334 239200
rect 77502 239144 79726 239200
rect 79894 239144 82026 239200
rect 82194 239144 84326 239200
rect 84494 239144 86626 239200
rect 86794 239144 88926 239200
rect 89094 239144 91226 239200
rect 91394 239144 93526 239200
rect 93694 239144 95918 239200
rect 96086 239144 98218 239200
rect 98386 239144 100518 239200
rect 100686 239144 102818 239200
rect 102986 239144 105118 239200
rect 105286 239144 107418 239200
rect 107586 239144 109718 239200
rect 109886 239144 112110 239200
rect 112278 239144 114410 239200
rect 114578 239144 116710 239200
rect 116878 239144 119010 239200
rect 119178 239144 121310 239200
rect 121478 239144 123610 239200
rect 123778 239144 126002 239200
rect 126170 239144 128302 239200
rect 128470 239144 130602 239200
rect 130770 239144 132902 239200
rect 133070 239144 135202 239200
rect 135370 239144 137502 239200
rect 137670 239144 139802 239200
rect 139970 239144 142194 239200
rect 142362 239144 144494 239200
rect 144662 239144 146794 239200
rect 146962 239144 149094 239200
rect 149262 239144 151394 239200
rect 151562 239144 153694 239200
rect 153862 239144 155994 239200
rect 156162 239144 158386 239200
rect 158554 239144 160686 239200
rect 160854 239144 162986 239200
rect 163154 239144 165286 239200
rect 165454 239144 167586 239200
rect 167754 239144 169886 239200
rect 170054 239144 172278 239200
rect 172446 239144 174578 239200
rect 174746 239144 176878 239200
rect 177046 239144 179178 239200
rect 179346 239144 181478 239200
rect 181646 239144 183778 239200
rect 183946 239144 186078 239200
rect 186246 239144 188470 239200
rect 188638 239144 190770 239200
rect 190938 239144 193070 239200
rect 193238 239144 195370 239200
rect 195538 239144 197670 239200
rect 197838 239144 199970 239200
rect 200138 239144 202270 239200
rect 202438 239144 204662 239200
rect 204830 239144 206962 239200
rect 207130 239144 209262 239200
rect 209430 239144 211562 239200
rect 211730 239144 213862 239200
rect 214030 239144 216162 239200
rect 216330 239144 218462 239200
rect 218630 239144 220854 239200
rect 221022 239144 223154 239200
rect 223322 239144 225454 239200
rect 225622 239144 227754 239200
rect 227922 239144 230054 239200
rect 230222 239144 232354 239200
rect 232522 239144 234746 239200
rect 234914 239144 237046 239200
rect 237214 239144 239346 239200
rect 239514 239144 241646 239200
rect 241814 239144 243946 239200
rect 244114 239144 246246 239200
rect 246414 239144 248546 239200
rect 248714 239144 250938 239200
rect 251106 239144 253238 239200
rect 253406 239144 255538 239200
rect 255706 239144 257838 239200
rect 258006 239144 260138 239200
rect 260306 239144 262438 239200
rect 262606 239144 264738 239200
rect 264906 239144 267130 239200
rect 267298 239144 269430 239200
rect 269598 239144 271730 239200
rect 271898 239144 274030 239200
rect 274198 239144 276330 239200
rect 276498 239144 276626 239200
rect 294 856 276626 239144
rect 406 800 790 856
rect 958 800 1342 856
rect 1510 800 1894 856
rect 2062 800 2446 856
rect 2614 800 2998 856
rect 3166 800 3550 856
rect 3718 800 4102 856
rect 4270 800 4746 856
rect 4914 800 5298 856
rect 5466 800 5850 856
rect 6018 800 6402 856
rect 6570 800 6954 856
rect 7122 800 7506 856
rect 7674 800 8058 856
rect 8226 800 8702 856
rect 8870 800 9254 856
rect 9422 800 9806 856
rect 9974 800 10358 856
rect 10526 800 10910 856
rect 11078 800 11462 856
rect 11630 800 12014 856
rect 12182 800 12566 856
rect 12734 800 13210 856
rect 13378 800 13762 856
rect 13930 800 14314 856
rect 14482 800 14866 856
rect 15034 800 15418 856
rect 15586 800 15970 856
rect 16138 800 16522 856
rect 16690 800 17166 856
rect 17334 800 17718 856
rect 17886 800 18270 856
rect 18438 800 18822 856
rect 18990 800 19374 856
rect 19542 800 19926 856
rect 20094 800 20478 856
rect 20646 800 21030 856
rect 21198 800 21674 856
rect 21842 800 22226 856
rect 22394 800 22778 856
rect 22946 800 23330 856
rect 23498 800 23882 856
rect 24050 800 24434 856
rect 24602 800 24986 856
rect 25154 800 25630 856
rect 25798 800 26182 856
rect 26350 800 26734 856
rect 26902 800 27286 856
rect 27454 800 27838 856
rect 28006 800 28390 856
rect 28558 800 28942 856
rect 29110 800 29586 856
rect 29754 800 30138 856
rect 30306 800 30690 856
rect 30858 800 31242 856
rect 31410 800 31794 856
rect 31962 800 32346 856
rect 32514 800 32898 856
rect 33066 800 33450 856
rect 33618 800 34094 856
rect 34262 800 34646 856
rect 34814 800 35198 856
rect 35366 800 35750 856
rect 35918 800 36302 856
rect 36470 800 36854 856
rect 37022 800 37406 856
rect 37574 800 38050 856
rect 38218 800 38602 856
rect 38770 800 39154 856
rect 39322 800 39706 856
rect 39874 800 40258 856
rect 40426 800 40810 856
rect 40978 800 41362 856
rect 41530 800 41914 856
rect 42082 800 42558 856
rect 42726 800 43110 856
rect 43278 800 43662 856
rect 43830 800 44214 856
rect 44382 800 44766 856
rect 44934 800 45318 856
rect 45486 800 45870 856
rect 46038 800 46514 856
rect 46682 800 47066 856
rect 47234 800 47618 856
rect 47786 800 48170 856
rect 48338 800 48722 856
rect 48890 800 49274 856
rect 49442 800 49826 856
rect 49994 800 50470 856
rect 50638 800 51022 856
rect 51190 800 51574 856
rect 51742 800 52126 856
rect 52294 800 52678 856
rect 52846 800 53230 856
rect 53398 800 53782 856
rect 53950 800 54334 856
rect 54502 800 54978 856
rect 55146 800 55530 856
rect 55698 800 56082 856
rect 56250 800 56634 856
rect 56802 800 57186 856
rect 57354 800 57738 856
rect 57906 800 58290 856
rect 58458 800 58934 856
rect 59102 800 59486 856
rect 59654 800 60038 856
rect 60206 800 60590 856
rect 60758 800 61142 856
rect 61310 800 61694 856
rect 61862 800 62246 856
rect 62414 800 62798 856
rect 62966 800 63442 856
rect 63610 800 63994 856
rect 64162 800 64546 856
rect 64714 800 65098 856
rect 65266 800 65650 856
rect 65818 800 66202 856
rect 66370 800 66754 856
rect 66922 800 67398 856
rect 67566 800 67950 856
rect 68118 800 68502 856
rect 68670 800 69054 856
rect 69222 800 69606 856
rect 69774 800 70158 856
rect 70326 800 70710 856
rect 70878 800 71354 856
rect 71522 800 71906 856
rect 72074 800 72458 856
rect 72626 800 73010 856
rect 73178 800 73562 856
rect 73730 800 74114 856
rect 74282 800 74666 856
rect 74834 800 75218 856
rect 75386 800 75862 856
rect 76030 800 76414 856
rect 76582 800 76966 856
rect 77134 800 77518 856
rect 77686 800 78070 856
rect 78238 800 78622 856
rect 78790 800 79174 856
rect 79342 800 79818 856
rect 79986 800 80370 856
rect 80538 800 80922 856
rect 81090 800 81474 856
rect 81642 800 82026 856
rect 82194 800 82578 856
rect 82746 800 83130 856
rect 83298 800 83682 856
rect 83850 800 84326 856
rect 84494 800 84878 856
rect 85046 800 85430 856
rect 85598 800 85982 856
rect 86150 800 86534 856
rect 86702 800 87086 856
rect 87254 800 87638 856
rect 87806 800 88282 856
rect 88450 800 88834 856
rect 89002 800 89386 856
rect 89554 800 89938 856
rect 90106 800 90490 856
rect 90658 800 91042 856
rect 91210 800 91594 856
rect 91762 800 92238 856
rect 92406 800 92790 856
rect 92958 800 93342 856
rect 93510 800 93894 856
rect 94062 800 94446 856
rect 94614 800 94998 856
rect 95166 800 95550 856
rect 95718 800 96102 856
rect 96270 800 96746 856
rect 96914 800 97298 856
rect 97466 800 97850 856
rect 98018 800 98402 856
rect 98570 800 98954 856
rect 99122 800 99506 856
rect 99674 800 100058 856
rect 100226 800 100702 856
rect 100870 800 101254 856
rect 101422 800 101806 856
rect 101974 800 102358 856
rect 102526 800 102910 856
rect 103078 800 103462 856
rect 103630 800 104014 856
rect 104182 800 104566 856
rect 104734 800 105210 856
rect 105378 800 105762 856
rect 105930 800 106314 856
rect 106482 800 106866 856
rect 107034 800 107418 856
rect 107586 800 107970 856
rect 108138 800 108522 856
rect 108690 800 109166 856
rect 109334 800 109718 856
rect 109886 800 110270 856
rect 110438 800 110822 856
rect 110990 800 111374 856
rect 111542 800 111926 856
rect 112094 800 112478 856
rect 112646 800 113122 856
rect 113290 800 113674 856
rect 113842 800 114226 856
rect 114394 800 114778 856
rect 114946 800 115330 856
rect 115498 800 115882 856
rect 116050 800 116434 856
rect 116602 800 116986 856
rect 117154 800 117630 856
rect 117798 800 118182 856
rect 118350 800 118734 856
rect 118902 800 119286 856
rect 119454 800 119838 856
rect 120006 800 120390 856
rect 120558 800 120942 856
rect 121110 800 121586 856
rect 121754 800 122138 856
rect 122306 800 122690 856
rect 122858 800 123242 856
rect 123410 800 123794 856
rect 123962 800 124346 856
rect 124514 800 124898 856
rect 125066 800 125450 856
rect 125618 800 126094 856
rect 126262 800 126646 856
rect 126814 800 127198 856
rect 127366 800 127750 856
rect 127918 800 128302 856
rect 128470 800 128854 856
rect 129022 800 129406 856
rect 129574 800 130050 856
rect 130218 800 130602 856
rect 130770 800 131154 856
rect 131322 800 131706 856
rect 131874 800 132258 856
rect 132426 800 132810 856
rect 132978 800 133362 856
rect 133530 800 134006 856
rect 134174 800 134558 856
rect 134726 800 135110 856
rect 135278 800 135662 856
rect 135830 800 136214 856
rect 136382 800 136766 856
rect 136934 800 137318 856
rect 137486 800 137870 856
rect 138038 800 138514 856
rect 138682 800 139066 856
rect 139234 800 139618 856
rect 139786 800 140170 856
rect 140338 800 140722 856
rect 140890 800 141274 856
rect 141442 800 141826 856
rect 141994 800 142470 856
rect 142638 800 143022 856
rect 143190 800 143574 856
rect 143742 800 144126 856
rect 144294 800 144678 856
rect 144846 800 145230 856
rect 145398 800 145782 856
rect 145950 800 146334 856
rect 146502 800 146978 856
rect 147146 800 147530 856
rect 147698 800 148082 856
rect 148250 800 148634 856
rect 148802 800 149186 856
rect 149354 800 149738 856
rect 149906 800 150290 856
rect 150458 800 150934 856
rect 151102 800 151486 856
rect 151654 800 152038 856
rect 152206 800 152590 856
rect 152758 800 153142 856
rect 153310 800 153694 856
rect 153862 800 154246 856
rect 154414 800 154890 856
rect 155058 800 155442 856
rect 155610 800 155994 856
rect 156162 800 156546 856
rect 156714 800 157098 856
rect 157266 800 157650 856
rect 157818 800 158202 856
rect 158370 800 158754 856
rect 158922 800 159398 856
rect 159566 800 159950 856
rect 160118 800 160502 856
rect 160670 800 161054 856
rect 161222 800 161606 856
rect 161774 800 162158 856
rect 162326 800 162710 856
rect 162878 800 163354 856
rect 163522 800 163906 856
rect 164074 800 164458 856
rect 164626 800 165010 856
rect 165178 800 165562 856
rect 165730 800 166114 856
rect 166282 800 166666 856
rect 166834 800 167218 856
rect 167386 800 167862 856
rect 168030 800 168414 856
rect 168582 800 168966 856
rect 169134 800 169518 856
rect 169686 800 170070 856
rect 170238 800 170622 856
rect 170790 800 171174 856
rect 171342 800 171818 856
rect 171986 800 172370 856
rect 172538 800 172922 856
rect 173090 800 173474 856
rect 173642 800 174026 856
rect 174194 800 174578 856
rect 174746 800 175130 856
rect 175298 800 175774 856
rect 175942 800 176326 856
rect 176494 800 176878 856
rect 177046 800 177430 856
rect 177598 800 177982 856
rect 178150 800 178534 856
rect 178702 800 179086 856
rect 179254 800 179638 856
rect 179806 800 180282 856
rect 180450 800 180834 856
rect 181002 800 181386 856
rect 181554 800 181938 856
rect 182106 800 182490 856
rect 182658 800 183042 856
rect 183210 800 183594 856
rect 183762 800 184238 856
rect 184406 800 184790 856
rect 184958 800 185342 856
rect 185510 800 185894 856
rect 186062 800 186446 856
rect 186614 800 186998 856
rect 187166 800 187550 856
rect 187718 800 188102 856
rect 188270 800 188746 856
rect 188914 800 189298 856
rect 189466 800 189850 856
rect 190018 800 190402 856
rect 190570 800 190954 856
rect 191122 800 191506 856
rect 191674 800 192058 856
rect 192226 800 192702 856
rect 192870 800 193254 856
rect 193422 800 193806 856
rect 193974 800 194358 856
rect 194526 800 194910 856
rect 195078 800 195462 856
rect 195630 800 196014 856
rect 196182 800 196658 856
rect 196826 800 197210 856
rect 197378 800 197762 856
rect 197930 800 198314 856
rect 198482 800 198866 856
rect 199034 800 199418 856
rect 199586 800 199970 856
rect 200138 800 200522 856
rect 200690 800 201166 856
rect 201334 800 201718 856
rect 201886 800 202270 856
rect 202438 800 202822 856
rect 202990 800 203374 856
rect 203542 800 203926 856
rect 204094 800 204478 856
rect 204646 800 205122 856
rect 205290 800 205674 856
rect 205842 800 206226 856
rect 206394 800 206778 856
rect 206946 800 207330 856
rect 207498 800 207882 856
rect 208050 800 208434 856
rect 208602 800 208986 856
rect 209154 800 209630 856
rect 209798 800 210182 856
rect 210350 800 210734 856
rect 210902 800 211286 856
rect 211454 800 211838 856
rect 212006 800 212390 856
rect 212558 800 212942 856
rect 213110 800 213586 856
rect 213754 800 214138 856
rect 214306 800 214690 856
rect 214858 800 215242 856
rect 215410 800 215794 856
rect 215962 800 216346 856
rect 216514 800 216898 856
rect 217066 800 217542 856
rect 217710 800 218094 856
rect 218262 800 218646 856
rect 218814 800 219198 856
rect 219366 800 219750 856
rect 219918 800 220302 856
rect 220470 800 220854 856
rect 221022 800 221406 856
rect 221574 800 222050 856
rect 222218 800 222602 856
rect 222770 800 223154 856
rect 223322 800 223706 856
rect 223874 800 224258 856
rect 224426 800 224810 856
rect 224978 800 225362 856
rect 225530 800 226006 856
rect 226174 800 226558 856
rect 226726 800 227110 856
rect 227278 800 227662 856
rect 227830 800 228214 856
rect 228382 800 228766 856
rect 228934 800 229318 856
rect 229486 800 229870 856
rect 230038 800 230514 856
rect 230682 800 231066 856
rect 231234 800 231618 856
rect 231786 800 232170 856
rect 232338 800 232722 856
rect 232890 800 233274 856
rect 233442 800 233826 856
rect 233994 800 234470 856
rect 234638 800 235022 856
rect 235190 800 235574 856
rect 235742 800 236126 856
rect 236294 800 236678 856
rect 236846 800 237230 856
rect 237398 800 237782 856
rect 237950 800 238426 856
rect 238594 800 238978 856
rect 239146 800 239530 856
rect 239698 800 240082 856
rect 240250 800 240634 856
rect 240802 800 241186 856
rect 241354 800 241738 856
rect 241906 800 242290 856
rect 242458 800 242934 856
rect 243102 800 243486 856
rect 243654 800 244038 856
rect 244206 800 244590 856
rect 244758 800 245142 856
rect 245310 800 245694 856
rect 245862 800 246246 856
rect 246414 800 246890 856
rect 247058 800 247442 856
rect 247610 800 247994 856
rect 248162 800 248546 856
rect 248714 800 249098 856
rect 249266 800 249650 856
rect 249818 800 250202 856
rect 250370 800 250754 856
rect 250922 800 251398 856
rect 251566 800 251950 856
rect 252118 800 252502 856
rect 252670 800 253054 856
rect 253222 800 253606 856
rect 253774 800 254158 856
rect 254326 800 254710 856
rect 254878 800 255354 856
rect 255522 800 255906 856
rect 256074 800 256458 856
rect 256626 800 257010 856
rect 257178 800 257562 856
rect 257730 800 258114 856
rect 258282 800 258666 856
rect 258834 800 259310 856
rect 259478 800 259862 856
rect 260030 800 260414 856
rect 260582 800 260966 856
rect 261134 800 261518 856
rect 261686 800 262070 856
rect 262238 800 262622 856
rect 262790 800 263174 856
rect 263342 800 263818 856
rect 263986 800 264370 856
rect 264538 800 264922 856
rect 265090 800 265474 856
rect 265642 800 266026 856
rect 266194 800 266578 856
rect 266746 800 267130 856
rect 267298 800 267774 856
rect 267942 800 268326 856
rect 268494 800 268878 856
rect 269046 800 269430 856
rect 269598 800 269982 856
rect 270150 800 270534 856
rect 270702 800 271086 856
rect 271254 800 271638 856
rect 271806 800 272282 856
rect 272450 800 272834 856
rect 273002 800 273386 856
rect 273554 800 273938 856
rect 274106 800 274490 856
rect 274658 800 275042 856
rect 275210 800 275594 856
rect 275762 800 276238 856
rect 276406 800 276626 856
<< metal3 >>
rect 279200 229032 280000 229152
rect 0 222776 800 222896
rect 279200 207272 280000 207392
rect 0 188504 800 188624
rect 279200 185376 280000 185496
rect 279200 163616 280000 163736
rect 0 154232 800 154352
rect 279200 141720 280000 141840
rect 0 119960 800 120080
rect 279200 119960 280000 120080
rect 279200 98064 280000 98184
rect 0 85688 800 85808
rect 279200 76304 280000 76424
rect 279200 54408 280000 54528
rect 0 51416 800 51536
rect 279200 32648 280000 32768
rect 0 17144 800 17264
rect 279200 10888 280000 11008
<< obsm3 >>
rect 289 229232 279200 237761
rect 289 228952 279120 229232
rect 289 222976 279200 228952
rect 880 222696 279200 222976
rect 289 207472 279200 222696
rect 289 207192 279120 207472
rect 289 188704 279200 207192
rect 880 188424 279200 188704
rect 289 185576 279200 188424
rect 289 185296 279120 185576
rect 289 163816 279200 185296
rect 289 163536 279120 163816
rect 289 154432 279200 163536
rect 880 154152 279200 154432
rect 289 141920 279200 154152
rect 289 141640 279120 141920
rect 289 120160 279200 141640
rect 880 119880 279120 120160
rect 289 98264 279200 119880
rect 289 97984 279120 98264
rect 289 85888 279200 97984
rect 880 85608 279200 85888
rect 289 76504 279200 85608
rect 289 76224 279120 76504
rect 289 54608 279200 76224
rect 289 54328 279120 54608
rect 289 51616 279200 54328
rect 880 51336 279200 51616
rect 289 32848 279200 51336
rect 289 32568 279120 32848
rect 289 17344 279200 32568
rect 880 17064 279200 17344
rect 289 11088 279200 17064
rect 289 10808 279120 11088
rect 289 851 279200 10808
<< metal4 >>
rect 4208 2128 4528 237776
rect 19568 2128 19888 237776
<< obsm4 >>
rect 34928 2128 265648 237776
<< labels >>
rlabel metal3 s 0 17144 800 17264 6 analog_io[0]
port 1 nsew default bidirectional
rlabel metal3 s 0 154232 800 154352 6 analog_io[10]
port 2 nsew default bidirectional
rlabel metal2 s 267186 239200 267242 240000 6 analog_io[11]
port 3 nsew default bidirectional
rlabel metal3 s 0 188504 800 188624 6 analog_io[12]
port 4 nsew default bidirectional
rlabel metal3 s 279200 54408 280000 54528 6 analog_io[13]
port 5 nsew default bidirectional
rlabel metal3 s 279200 76304 280000 76424 6 analog_io[14]
port 6 nsew default bidirectional
rlabel metal2 s 269486 239200 269542 240000 6 analog_io[15]
port 7 nsew default bidirectional
rlabel metal3 s 0 222776 800 222896 6 analog_io[16]
port 8 nsew default bidirectional
rlabel metal2 s 271786 239200 271842 240000 6 analog_io[17]
port 9 nsew default bidirectional
rlabel metal2 s 274086 239200 274142 240000 6 analog_io[18]
port 10 nsew default bidirectional
rlabel metal2 s 278502 0 278558 800 6 analog_io[19]
port 11 nsew default bidirectional
rlabel metal2 s 264794 239200 264850 240000 6 analog_io[1]
port 12 nsew default bidirectional
rlabel metal3 s 279200 98064 280000 98184 6 analog_io[20]
port 13 nsew default bidirectional
rlabel metal2 s 279054 0 279110 800 6 analog_io[21]
port 14 nsew default bidirectional
rlabel metal3 s 279200 119960 280000 120080 6 analog_io[22]
port 15 nsew default bidirectional
rlabel metal3 s 279200 141720 280000 141840 6 analog_io[23]
port 16 nsew default bidirectional
rlabel metal2 s 276386 239200 276442 240000 6 analog_io[24]
port 17 nsew default bidirectional
rlabel metal3 s 279200 163616 280000 163736 6 analog_io[25]
port 18 nsew default bidirectional
rlabel metal3 s 279200 185376 280000 185496 6 analog_io[26]
port 19 nsew default bidirectional
rlabel metal3 s 279200 207272 280000 207392 6 analog_io[27]
port 20 nsew default bidirectional
rlabel metal3 s 279200 229032 280000 229152 6 analog_io[28]
port 21 nsew default bidirectional
rlabel metal2 s 278686 239200 278742 240000 6 analog_io[29]
port 22 nsew default bidirectional
rlabel metal2 s 276846 0 276902 800 6 analog_io[2]
port 23 nsew default bidirectional
rlabel metal2 s 279606 0 279662 800 6 analog_io[30]
port 24 nsew default bidirectional
rlabel metal3 s 0 51416 800 51536 6 analog_io[3]
port 25 nsew default bidirectional
rlabel metal2 s 277398 0 277454 800 6 analog_io[4]
port 26 nsew default bidirectional
rlabel metal3 s 0 85688 800 85808 6 analog_io[5]
port 27 nsew default bidirectional
rlabel metal3 s 0 119960 800 120080 6 analog_io[6]
port 28 nsew default bidirectional
rlabel metal3 s 279200 10888 280000 11008 6 analog_io[7]
port 29 nsew default bidirectional
rlabel metal2 s 277950 0 278006 800 6 analog_io[8]
port 30 nsew default bidirectional
rlabel metal3 s 279200 32648 280000 32768 6 analog_io[9]
port 31 nsew default bidirectional
rlabel metal2 s 1122 239200 1178 240000 6 io_in[0]
port 32 nsew default input
rlabel metal2 s 70490 239200 70546 240000 6 io_in[10]
port 33 nsew default input
rlabel metal2 s 77390 239200 77446 240000 6 io_in[11]
port 34 nsew default input
rlabel metal2 s 84382 239200 84438 240000 6 io_in[12]
port 35 nsew default input
rlabel metal2 s 91282 239200 91338 240000 6 io_in[13]
port 36 nsew default input
rlabel metal2 s 98274 239200 98330 240000 6 io_in[14]
port 37 nsew default input
rlabel metal2 s 105174 239200 105230 240000 6 io_in[15]
port 38 nsew default input
rlabel metal2 s 112166 239200 112222 240000 6 io_in[16]
port 39 nsew default input
rlabel metal2 s 119066 239200 119122 240000 6 io_in[17]
port 40 nsew default input
rlabel metal2 s 126058 239200 126114 240000 6 io_in[18]
port 41 nsew default input
rlabel metal2 s 132958 239200 133014 240000 6 io_in[19]
port 42 nsew default input
rlabel metal2 s 8022 239200 8078 240000 6 io_in[1]
port 43 nsew default input
rlabel metal2 s 139858 239200 139914 240000 6 io_in[20]
port 44 nsew default input
rlabel metal2 s 146850 239200 146906 240000 6 io_in[21]
port 45 nsew default input
rlabel metal2 s 153750 239200 153806 240000 6 io_in[22]
port 46 nsew default input
rlabel metal2 s 160742 239200 160798 240000 6 io_in[23]
port 47 nsew default input
rlabel metal2 s 167642 239200 167698 240000 6 io_in[24]
port 48 nsew default input
rlabel metal2 s 174634 239200 174690 240000 6 io_in[25]
port 49 nsew default input
rlabel metal2 s 181534 239200 181590 240000 6 io_in[26]
port 50 nsew default input
rlabel metal2 s 188526 239200 188582 240000 6 io_in[27]
port 51 nsew default input
rlabel metal2 s 195426 239200 195482 240000 6 io_in[28]
port 52 nsew default input
rlabel metal2 s 202326 239200 202382 240000 6 io_in[29]
port 53 nsew default input
rlabel metal2 s 14922 239200 14978 240000 6 io_in[2]
port 54 nsew default input
rlabel metal2 s 209318 239200 209374 240000 6 io_in[30]
port 55 nsew default input
rlabel metal2 s 216218 239200 216274 240000 6 io_in[31]
port 56 nsew default input
rlabel metal2 s 223210 239200 223266 240000 6 io_in[32]
port 57 nsew default input
rlabel metal2 s 230110 239200 230166 240000 6 io_in[33]
port 58 nsew default input
rlabel metal2 s 237102 239200 237158 240000 6 io_in[34]
port 59 nsew default input
rlabel metal2 s 244002 239200 244058 240000 6 io_in[35]
port 60 nsew default input
rlabel metal2 s 250994 239200 251050 240000 6 io_in[36]
port 61 nsew default input
rlabel metal2 s 257894 239200 257950 240000 6 io_in[37]
port 62 nsew default input
rlabel metal2 s 21914 239200 21970 240000 6 io_in[3]
port 63 nsew default input
rlabel metal2 s 28814 239200 28870 240000 6 io_in[4]
port 64 nsew default input
rlabel metal2 s 35806 239200 35862 240000 6 io_in[5]
port 65 nsew default input
rlabel metal2 s 42706 239200 42762 240000 6 io_in[6]
port 66 nsew default input
rlabel metal2 s 49698 239200 49754 240000 6 io_in[7]
port 67 nsew default input
rlabel metal2 s 56598 239200 56654 240000 6 io_in[8]
port 68 nsew default input
rlabel metal2 s 63590 239200 63646 240000 6 io_in[9]
port 69 nsew default input
rlabel metal2 s 3422 239200 3478 240000 6 io_oeb[0]
port 70 nsew default output
rlabel metal2 s 72790 239200 72846 240000 6 io_oeb[10]
port 71 nsew default output
rlabel metal2 s 79782 239200 79838 240000 6 io_oeb[11]
port 72 nsew default output
rlabel metal2 s 86682 239200 86738 240000 6 io_oeb[12]
port 73 nsew default output
rlabel metal2 s 93582 239200 93638 240000 6 io_oeb[13]
port 74 nsew default output
rlabel metal2 s 100574 239200 100630 240000 6 io_oeb[14]
port 75 nsew default output
rlabel metal2 s 107474 239200 107530 240000 6 io_oeb[15]
port 76 nsew default output
rlabel metal2 s 114466 239200 114522 240000 6 io_oeb[16]
port 77 nsew default output
rlabel metal2 s 121366 239200 121422 240000 6 io_oeb[17]
port 78 nsew default output
rlabel metal2 s 128358 239200 128414 240000 6 io_oeb[18]
port 79 nsew default output
rlabel metal2 s 135258 239200 135314 240000 6 io_oeb[19]
port 80 nsew default output
rlabel metal2 s 10322 239200 10378 240000 6 io_oeb[1]
port 81 nsew default output
rlabel metal2 s 142250 239200 142306 240000 6 io_oeb[20]
port 82 nsew default output
rlabel metal2 s 149150 239200 149206 240000 6 io_oeb[21]
port 83 nsew default output
rlabel metal2 s 156050 239200 156106 240000 6 io_oeb[22]
port 84 nsew default output
rlabel metal2 s 163042 239200 163098 240000 6 io_oeb[23]
port 85 nsew default output
rlabel metal2 s 169942 239200 169998 240000 6 io_oeb[24]
port 86 nsew default output
rlabel metal2 s 176934 239200 176990 240000 6 io_oeb[25]
port 87 nsew default output
rlabel metal2 s 183834 239200 183890 240000 6 io_oeb[26]
port 88 nsew default output
rlabel metal2 s 190826 239200 190882 240000 6 io_oeb[27]
port 89 nsew default output
rlabel metal2 s 197726 239200 197782 240000 6 io_oeb[28]
port 90 nsew default output
rlabel metal2 s 204718 239200 204774 240000 6 io_oeb[29]
port 91 nsew default output
rlabel metal2 s 17314 239200 17370 240000 6 io_oeb[2]
port 92 nsew default output
rlabel metal2 s 211618 239200 211674 240000 6 io_oeb[30]
port 93 nsew default output
rlabel metal2 s 218518 239200 218574 240000 6 io_oeb[31]
port 94 nsew default output
rlabel metal2 s 225510 239200 225566 240000 6 io_oeb[32]
port 95 nsew default output
rlabel metal2 s 232410 239200 232466 240000 6 io_oeb[33]
port 96 nsew default output
rlabel metal2 s 239402 239200 239458 240000 6 io_oeb[34]
port 97 nsew default output
rlabel metal2 s 246302 239200 246358 240000 6 io_oeb[35]
port 98 nsew default output
rlabel metal2 s 253294 239200 253350 240000 6 io_oeb[36]
port 99 nsew default output
rlabel metal2 s 260194 239200 260250 240000 6 io_oeb[37]
port 100 nsew default output
rlabel metal2 s 24214 239200 24270 240000 6 io_oeb[3]
port 101 nsew default output
rlabel metal2 s 31114 239200 31170 240000 6 io_oeb[4]
port 102 nsew default output
rlabel metal2 s 38106 239200 38162 240000 6 io_oeb[5]
port 103 nsew default output
rlabel metal2 s 45006 239200 45062 240000 6 io_oeb[6]
port 104 nsew default output
rlabel metal2 s 51998 239200 52054 240000 6 io_oeb[7]
port 105 nsew default output
rlabel metal2 s 58898 239200 58954 240000 6 io_oeb[8]
port 106 nsew default output
rlabel metal2 s 65890 239200 65946 240000 6 io_oeb[9]
port 107 nsew default output
rlabel metal2 s 5722 239200 5778 240000 6 io_out[0]
port 108 nsew default output
rlabel metal2 s 75090 239200 75146 240000 6 io_out[10]
port 109 nsew default output
rlabel metal2 s 82082 239200 82138 240000 6 io_out[11]
port 110 nsew default output
rlabel metal2 s 88982 239200 89038 240000 6 io_out[12]
port 111 nsew default output
rlabel metal2 s 95974 239200 96030 240000 6 io_out[13]
port 112 nsew default output
rlabel metal2 s 102874 239200 102930 240000 6 io_out[14]
port 113 nsew default output
rlabel metal2 s 109774 239200 109830 240000 6 io_out[15]
port 114 nsew default output
rlabel metal2 s 116766 239200 116822 240000 6 io_out[16]
port 115 nsew default output
rlabel metal2 s 123666 239200 123722 240000 6 io_out[17]
port 116 nsew default output
rlabel metal2 s 130658 239200 130714 240000 6 io_out[18]
port 117 nsew default output
rlabel metal2 s 137558 239200 137614 240000 6 io_out[19]
port 118 nsew default output
rlabel metal2 s 12622 239200 12678 240000 6 io_out[1]
port 119 nsew default output
rlabel metal2 s 144550 239200 144606 240000 6 io_out[20]
port 120 nsew default output
rlabel metal2 s 151450 239200 151506 240000 6 io_out[21]
port 121 nsew default output
rlabel metal2 s 158442 239200 158498 240000 6 io_out[22]
port 122 nsew default output
rlabel metal2 s 165342 239200 165398 240000 6 io_out[23]
port 123 nsew default output
rlabel metal2 s 172334 239200 172390 240000 6 io_out[24]
port 124 nsew default output
rlabel metal2 s 179234 239200 179290 240000 6 io_out[25]
port 125 nsew default output
rlabel metal2 s 186134 239200 186190 240000 6 io_out[26]
port 126 nsew default output
rlabel metal2 s 193126 239200 193182 240000 6 io_out[27]
port 127 nsew default output
rlabel metal2 s 200026 239200 200082 240000 6 io_out[28]
port 128 nsew default output
rlabel metal2 s 207018 239200 207074 240000 6 io_out[29]
port 129 nsew default output
rlabel metal2 s 19614 239200 19670 240000 6 io_out[2]
port 130 nsew default output
rlabel metal2 s 213918 239200 213974 240000 6 io_out[30]
port 131 nsew default output
rlabel metal2 s 220910 239200 220966 240000 6 io_out[31]
port 132 nsew default output
rlabel metal2 s 227810 239200 227866 240000 6 io_out[32]
port 133 nsew default output
rlabel metal2 s 234802 239200 234858 240000 6 io_out[33]
port 134 nsew default output
rlabel metal2 s 241702 239200 241758 240000 6 io_out[34]
port 135 nsew default output
rlabel metal2 s 248602 239200 248658 240000 6 io_out[35]
port 136 nsew default output
rlabel metal2 s 255594 239200 255650 240000 6 io_out[36]
port 137 nsew default output
rlabel metal2 s 262494 239200 262550 240000 6 io_out[37]
port 138 nsew default output
rlabel metal2 s 26514 239200 26570 240000 6 io_out[3]
port 139 nsew default output
rlabel metal2 s 33506 239200 33562 240000 6 io_out[4]
port 140 nsew default output
rlabel metal2 s 40406 239200 40462 240000 6 io_out[5]
port 141 nsew default output
rlabel metal2 s 47306 239200 47362 240000 6 io_out[6]
port 142 nsew default output
rlabel metal2 s 54298 239200 54354 240000 6 io_out[7]
port 143 nsew default output
rlabel metal2 s 61198 239200 61254 240000 6 io_out[8]
port 144 nsew default output
rlabel metal2 s 68190 239200 68246 240000 6 io_out[9]
port 145 nsew default output
rlabel metal2 s 60094 0 60150 800 6 la_data_in[0]
port 146 nsew default input
rlabel metal2 s 229374 0 229430 800 6 la_data_in[100]
port 147 nsew default input
rlabel metal2 s 231122 0 231178 800 6 la_data_in[101]
port 148 nsew default input
rlabel metal2 s 232778 0 232834 800 6 la_data_in[102]
port 149 nsew default input
rlabel metal2 s 234526 0 234582 800 6 la_data_in[103]
port 150 nsew default input
rlabel metal2 s 236182 0 236238 800 6 la_data_in[104]
port 151 nsew default input
rlabel metal2 s 237838 0 237894 800 6 la_data_in[105]
port 152 nsew default input
rlabel metal2 s 239586 0 239642 800 6 la_data_in[106]
port 153 nsew default input
rlabel metal2 s 241242 0 241298 800 6 la_data_in[107]
port 154 nsew default input
rlabel metal2 s 242990 0 243046 800 6 la_data_in[108]
port 155 nsew default input
rlabel metal2 s 244646 0 244702 800 6 la_data_in[109]
port 156 nsew default input
rlabel metal2 s 77022 0 77078 800 6 la_data_in[10]
port 157 nsew default input
rlabel metal2 s 246302 0 246358 800 6 la_data_in[110]
port 158 nsew default input
rlabel metal2 s 248050 0 248106 800 6 la_data_in[111]
port 159 nsew default input
rlabel metal2 s 249706 0 249762 800 6 la_data_in[112]
port 160 nsew default input
rlabel metal2 s 251454 0 251510 800 6 la_data_in[113]
port 161 nsew default input
rlabel metal2 s 253110 0 253166 800 6 la_data_in[114]
port 162 nsew default input
rlabel metal2 s 254766 0 254822 800 6 la_data_in[115]
port 163 nsew default input
rlabel metal2 s 256514 0 256570 800 6 la_data_in[116]
port 164 nsew default input
rlabel metal2 s 258170 0 258226 800 6 la_data_in[117]
port 165 nsew default input
rlabel metal2 s 259918 0 259974 800 6 la_data_in[118]
port 166 nsew default input
rlabel metal2 s 261574 0 261630 800 6 la_data_in[119]
port 167 nsew default input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[11]
port 168 nsew default input
rlabel metal2 s 263230 0 263286 800 6 la_data_in[120]
port 169 nsew default input
rlabel metal2 s 264978 0 265034 800 6 la_data_in[121]
port 170 nsew default input
rlabel metal2 s 266634 0 266690 800 6 la_data_in[122]
port 171 nsew default input
rlabel metal2 s 268382 0 268438 800 6 la_data_in[123]
port 172 nsew default input
rlabel metal2 s 270038 0 270094 800 6 la_data_in[124]
port 173 nsew default input
rlabel metal2 s 271694 0 271750 800 6 la_data_in[125]
port 174 nsew default input
rlabel metal2 s 273442 0 273498 800 6 la_data_in[126]
port 175 nsew default input
rlabel metal2 s 275098 0 275154 800 6 la_data_in[127]
port 176 nsew default input
rlabel metal2 s 80426 0 80482 800 6 la_data_in[12]
port 177 nsew default input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[13]
port 178 nsew default input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[14]
port 179 nsew default input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[15]
port 180 nsew default input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[16]
port 181 nsew default input
rlabel metal2 s 88890 0 88946 800 6 la_data_in[17]
port 182 nsew default input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[18]
port 183 nsew default input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[19]
port 184 nsew default input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[1]
port 185 nsew default input
rlabel metal2 s 93950 0 94006 800 6 la_data_in[20]
port 186 nsew default input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[21]
port 187 nsew default input
rlabel metal2 s 97354 0 97410 800 6 la_data_in[22]
port 188 nsew default input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[23]
port 189 nsew default input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[24]
port 190 nsew default input
rlabel metal2 s 102414 0 102470 800 6 la_data_in[25]
port 191 nsew default input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[26]
port 192 nsew default input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[27]
port 193 nsew default input
rlabel metal2 s 107474 0 107530 800 6 la_data_in[28]
port 194 nsew default input
rlabel metal2 s 109222 0 109278 800 6 la_data_in[29]
port 195 nsew default input
rlabel metal2 s 63498 0 63554 800 6 la_data_in[2]
port 196 nsew default input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[30]
port 197 nsew default input
rlabel metal2 s 112534 0 112590 800 6 la_data_in[31]
port 198 nsew default input
rlabel metal2 s 114282 0 114338 800 6 la_data_in[32]
port 199 nsew default input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[33]
port 200 nsew default input
rlabel metal2 s 117686 0 117742 800 6 la_data_in[34]
port 201 nsew default input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[35]
port 202 nsew default input
rlabel metal2 s 120998 0 121054 800 6 la_data_in[36]
port 203 nsew default input
rlabel metal2 s 122746 0 122802 800 6 la_data_in[37]
port 204 nsew default input
rlabel metal2 s 124402 0 124458 800 6 la_data_in[38]
port 205 nsew default input
rlabel metal2 s 126150 0 126206 800 6 la_data_in[39]
port 206 nsew default input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[3]
port 207 nsew default input
rlabel metal2 s 127806 0 127862 800 6 la_data_in[40]
port 208 nsew default input
rlabel metal2 s 129462 0 129518 800 6 la_data_in[41]
port 209 nsew default input
rlabel metal2 s 131210 0 131266 800 6 la_data_in[42]
port 210 nsew default input
rlabel metal2 s 132866 0 132922 800 6 la_data_in[43]
port 211 nsew default input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[44]
port 212 nsew default input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[45]
port 213 nsew default input
rlabel metal2 s 137926 0 137982 800 6 la_data_in[46]
port 214 nsew default input
rlabel metal2 s 139674 0 139730 800 6 la_data_in[47]
port 215 nsew default input
rlabel metal2 s 141330 0 141386 800 6 la_data_in[48]
port 216 nsew default input
rlabel metal2 s 143078 0 143134 800 6 la_data_in[49]
port 217 nsew default input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[4]
port 218 nsew default input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[50]
port 219 nsew default input
rlabel metal2 s 146390 0 146446 800 6 la_data_in[51]
port 220 nsew default input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[52]
port 221 nsew default input
rlabel metal2 s 149794 0 149850 800 6 la_data_in[53]
port 222 nsew default input
rlabel metal2 s 151542 0 151598 800 6 la_data_in[54]
port 223 nsew default input
rlabel metal2 s 153198 0 153254 800 6 la_data_in[55]
port 224 nsew default input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[56]
port 225 nsew default input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[57]
port 226 nsew default input
rlabel metal2 s 158258 0 158314 800 6 la_data_in[58]
port 227 nsew default input
rlabel metal2 s 160006 0 160062 800 6 la_data_in[59]
port 228 nsew default input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[5]
port 229 nsew default input
rlabel metal2 s 161662 0 161718 800 6 la_data_in[60]
port 230 nsew default input
rlabel metal2 s 163410 0 163466 800 6 la_data_in[61]
port 231 nsew default input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[62]
port 232 nsew default input
rlabel metal2 s 166722 0 166778 800 6 la_data_in[63]
port 233 nsew default input
rlabel metal2 s 168470 0 168526 800 6 la_data_in[64]
port 234 nsew default input
rlabel metal2 s 170126 0 170182 800 6 la_data_in[65]
port 235 nsew default input
rlabel metal2 s 171874 0 171930 800 6 la_data_in[66]
port 236 nsew default input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[67]
port 237 nsew default input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[68]
port 238 nsew default input
rlabel metal2 s 176934 0 176990 800 6 la_data_in[69]
port 239 nsew default input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[6]
port 240 nsew default input
rlabel metal2 s 178590 0 178646 800 6 la_data_in[70]
port 241 nsew default input
rlabel metal2 s 180338 0 180394 800 6 la_data_in[71]
port 242 nsew default input
rlabel metal2 s 181994 0 182050 800 6 la_data_in[72]
port 243 nsew default input
rlabel metal2 s 183650 0 183706 800 6 la_data_in[73]
port 244 nsew default input
rlabel metal2 s 185398 0 185454 800 6 la_data_in[74]
port 245 nsew default input
rlabel metal2 s 187054 0 187110 800 6 la_data_in[75]
port 246 nsew default input
rlabel metal2 s 188802 0 188858 800 6 la_data_in[76]
port 247 nsew default input
rlabel metal2 s 190458 0 190514 800 6 la_data_in[77]
port 248 nsew default input
rlabel metal2 s 192114 0 192170 800 6 la_data_in[78]
port 249 nsew default input
rlabel metal2 s 193862 0 193918 800 6 la_data_in[79]
port 250 nsew default input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[7]
port 251 nsew default input
rlabel metal2 s 195518 0 195574 800 6 la_data_in[80]
port 252 nsew default input
rlabel metal2 s 197266 0 197322 800 6 la_data_in[81]
port 253 nsew default input
rlabel metal2 s 198922 0 198978 800 6 la_data_in[82]
port 254 nsew default input
rlabel metal2 s 200578 0 200634 800 6 la_data_in[83]
port 255 nsew default input
rlabel metal2 s 202326 0 202382 800 6 la_data_in[84]
port 256 nsew default input
rlabel metal2 s 203982 0 204038 800 6 la_data_in[85]
port 257 nsew default input
rlabel metal2 s 205730 0 205786 800 6 la_data_in[86]
port 258 nsew default input
rlabel metal2 s 207386 0 207442 800 6 la_data_in[87]
port 259 nsew default input
rlabel metal2 s 209042 0 209098 800 6 la_data_in[88]
port 260 nsew default input
rlabel metal2 s 210790 0 210846 800 6 la_data_in[89]
port 261 nsew default input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[8]
port 262 nsew default input
rlabel metal2 s 212446 0 212502 800 6 la_data_in[90]
port 263 nsew default input
rlabel metal2 s 214194 0 214250 800 6 la_data_in[91]
port 264 nsew default input
rlabel metal2 s 215850 0 215906 800 6 la_data_in[92]
port 265 nsew default input
rlabel metal2 s 217598 0 217654 800 6 la_data_in[93]
port 266 nsew default input
rlabel metal2 s 219254 0 219310 800 6 la_data_in[94]
port 267 nsew default input
rlabel metal2 s 220910 0 220966 800 6 la_data_in[95]
port 268 nsew default input
rlabel metal2 s 222658 0 222714 800 6 la_data_in[96]
port 269 nsew default input
rlabel metal2 s 224314 0 224370 800 6 la_data_in[97]
port 270 nsew default input
rlabel metal2 s 226062 0 226118 800 6 la_data_in[98]
port 271 nsew default input
rlabel metal2 s 227718 0 227774 800 6 la_data_in[99]
port 272 nsew default input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[9]
port 273 nsew default input
rlabel metal2 s 60646 0 60702 800 6 la_data_out[0]
port 274 nsew default output
rlabel metal2 s 229926 0 229982 800 6 la_data_out[100]
port 275 nsew default output
rlabel metal2 s 231674 0 231730 800 6 la_data_out[101]
port 276 nsew default output
rlabel metal2 s 233330 0 233386 800 6 la_data_out[102]
port 277 nsew default output
rlabel metal2 s 235078 0 235134 800 6 la_data_out[103]
port 278 nsew default output
rlabel metal2 s 236734 0 236790 800 6 la_data_out[104]
port 279 nsew default output
rlabel metal2 s 238482 0 238538 800 6 la_data_out[105]
port 280 nsew default output
rlabel metal2 s 240138 0 240194 800 6 la_data_out[106]
port 281 nsew default output
rlabel metal2 s 241794 0 241850 800 6 la_data_out[107]
port 282 nsew default output
rlabel metal2 s 243542 0 243598 800 6 la_data_out[108]
port 283 nsew default output
rlabel metal2 s 245198 0 245254 800 6 la_data_out[109]
port 284 nsew default output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[10]
port 285 nsew default output
rlabel metal2 s 246946 0 247002 800 6 la_data_out[110]
port 286 nsew default output
rlabel metal2 s 248602 0 248658 800 6 la_data_out[111]
port 287 nsew default output
rlabel metal2 s 250258 0 250314 800 6 la_data_out[112]
port 288 nsew default output
rlabel metal2 s 252006 0 252062 800 6 la_data_out[113]
port 289 nsew default output
rlabel metal2 s 253662 0 253718 800 6 la_data_out[114]
port 290 nsew default output
rlabel metal2 s 255410 0 255466 800 6 la_data_out[115]
port 291 nsew default output
rlabel metal2 s 257066 0 257122 800 6 la_data_out[116]
port 292 nsew default output
rlabel metal2 s 258722 0 258778 800 6 la_data_out[117]
port 293 nsew default output
rlabel metal2 s 260470 0 260526 800 6 la_data_out[118]
port 294 nsew default output
rlabel metal2 s 262126 0 262182 800 6 la_data_out[119]
port 295 nsew default output
rlabel metal2 s 79230 0 79286 800 6 la_data_out[11]
port 296 nsew default output
rlabel metal2 s 263874 0 263930 800 6 la_data_out[120]
port 297 nsew default output
rlabel metal2 s 265530 0 265586 800 6 la_data_out[121]
port 298 nsew default output
rlabel metal2 s 267186 0 267242 800 6 la_data_out[122]
port 299 nsew default output
rlabel metal2 s 268934 0 268990 800 6 la_data_out[123]
port 300 nsew default output
rlabel metal2 s 270590 0 270646 800 6 la_data_out[124]
port 301 nsew default output
rlabel metal2 s 272338 0 272394 800 6 la_data_out[125]
port 302 nsew default output
rlabel metal2 s 273994 0 274050 800 6 la_data_out[126]
port 303 nsew default output
rlabel metal2 s 275650 0 275706 800 6 la_data_out[127]
port 304 nsew default output
rlabel metal2 s 80978 0 81034 800 6 la_data_out[12]
port 305 nsew default output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[13]
port 306 nsew default output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[14]
port 307 nsew default output
rlabel metal2 s 86038 0 86094 800 6 la_data_out[15]
port 308 nsew default output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[16]
port 309 nsew default output
rlabel metal2 s 89442 0 89498 800 6 la_data_out[17]
port 310 nsew default output
rlabel metal2 s 91098 0 91154 800 6 la_data_out[18]
port 311 nsew default output
rlabel metal2 s 92846 0 92902 800 6 la_data_out[19]
port 312 nsew default output
rlabel metal2 s 62302 0 62358 800 6 la_data_out[1]
port 313 nsew default output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[20]
port 314 nsew default output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[21]
port 315 nsew default output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[22]
port 316 nsew default output
rlabel metal2 s 99562 0 99618 800 6 la_data_out[23]
port 317 nsew default output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[24]
port 318 nsew default output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[25]
port 319 nsew default output
rlabel metal2 s 104622 0 104678 800 6 la_data_out[26]
port 320 nsew default output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[27]
port 321 nsew default output
rlabel metal2 s 108026 0 108082 800 6 la_data_out[28]
port 322 nsew default output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[29]
port 323 nsew default output
rlabel metal2 s 64050 0 64106 800 6 la_data_out[2]
port 324 nsew default output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[30]
port 325 nsew default output
rlabel metal2 s 113178 0 113234 800 6 la_data_out[31]
port 326 nsew default output
rlabel metal2 s 114834 0 114890 800 6 la_data_out[32]
port 327 nsew default output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[33]
port 328 nsew default output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[34]
port 329 nsew default output
rlabel metal2 s 119894 0 119950 800 6 la_data_out[35]
port 330 nsew default output
rlabel metal2 s 121642 0 121698 800 6 la_data_out[36]
port 331 nsew default output
rlabel metal2 s 123298 0 123354 800 6 la_data_out[37]
port 332 nsew default output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[38]
port 333 nsew default output
rlabel metal2 s 126702 0 126758 800 6 la_data_out[39]
port 334 nsew default output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[3]
port 335 nsew default output
rlabel metal2 s 128358 0 128414 800 6 la_data_out[40]
port 336 nsew default output
rlabel metal2 s 130106 0 130162 800 6 la_data_out[41]
port 337 nsew default output
rlabel metal2 s 131762 0 131818 800 6 la_data_out[42]
port 338 nsew default output
rlabel metal2 s 133418 0 133474 800 6 la_data_out[43]
port 339 nsew default output
rlabel metal2 s 135166 0 135222 800 6 la_data_out[44]
port 340 nsew default output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[45]
port 341 nsew default output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[46]
port 342 nsew default output
rlabel metal2 s 140226 0 140282 800 6 la_data_out[47]
port 343 nsew default output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[48]
port 344 nsew default output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[49]
port 345 nsew default output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[4]
port 346 nsew default output
rlabel metal2 s 145286 0 145342 800 6 la_data_out[50]
port 347 nsew default output
rlabel metal2 s 147034 0 147090 800 6 la_data_out[51]
port 348 nsew default output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[52]
port 349 nsew default output
rlabel metal2 s 150346 0 150402 800 6 la_data_out[53]
port 350 nsew default output
rlabel metal2 s 152094 0 152150 800 6 la_data_out[54]
port 351 nsew default output
rlabel metal2 s 153750 0 153806 800 6 la_data_out[55]
port 352 nsew default output
rlabel metal2 s 155498 0 155554 800 6 la_data_out[56]
port 353 nsew default output
rlabel metal2 s 157154 0 157210 800 6 la_data_out[57]
port 354 nsew default output
rlabel metal2 s 158810 0 158866 800 6 la_data_out[58]
port 355 nsew default output
rlabel metal2 s 160558 0 160614 800 6 la_data_out[59]
port 356 nsew default output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[5]
port 357 nsew default output
rlabel metal2 s 162214 0 162270 800 6 la_data_out[60]
port 358 nsew default output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[61]
port 359 nsew default output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[62]
port 360 nsew default output
rlabel metal2 s 167274 0 167330 800 6 la_data_out[63]
port 361 nsew default output
rlabel metal2 s 169022 0 169078 800 6 la_data_out[64]
port 362 nsew default output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[65]
port 363 nsew default output
rlabel metal2 s 172426 0 172482 800 6 la_data_out[66]
port 364 nsew default output
rlabel metal2 s 174082 0 174138 800 6 la_data_out[67]
port 365 nsew default output
rlabel metal2 s 175830 0 175886 800 6 la_data_out[68]
port 366 nsew default output
rlabel metal2 s 177486 0 177542 800 6 la_data_out[69]
port 367 nsew default output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[6]
port 368 nsew default output
rlabel metal2 s 179142 0 179198 800 6 la_data_out[70]
port 369 nsew default output
rlabel metal2 s 180890 0 180946 800 6 la_data_out[71]
port 370 nsew default output
rlabel metal2 s 182546 0 182602 800 6 la_data_out[72]
port 371 nsew default output
rlabel metal2 s 184294 0 184350 800 6 la_data_out[73]
port 372 nsew default output
rlabel metal2 s 185950 0 186006 800 6 la_data_out[74]
port 373 nsew default output
rlabel metal2 s 187606 0 187662 800 6 la_data_out[75]
port 374 nsew default output
rlabel metal2 s 189354 0 189410 800 6 la_data_out[76]
port 375 nsew default output
rlabel metal2 s 191010 0 191066 800 6 la_data_out[77]
port 376 nsew default output
rlabel metal2 s 192758 0 192814 800 6 la_data_out[78]
port 377 nsew default output
rlabel metal2 s 194414 0 194470 800 6 la_data_out[79]
port 378 nsew default output
rlabel metal2 s 72514 0 72570 800 6 la_data_out[7]
port 379 nsew default output
rlabel metal2 s 196070 0 196126 800 6 la_data_out[80]
port 380 nsew default output
rlabel metal2 s 197818 0 197874 800 6 la_data_out[81]
port 381 nsew default output
rlabel metal2 s 199474 0 199530 800 6 la_data_out[82]
port 382 nsew default output
rlabel metal2 s 201222 0 201278 800 6 la_data_out[83]
port 383 nsew default output
rlabel metal2 s 202878 0 202934 800 6 la_data_out[84]
port 384 nsew default output
rlabel metal2 s 204534 0 204590 800 6 la_data_out[85]
port 385 nsew default output
rlabel metal2 s 206282 0 206338 800 6 la_data_out[86]
port 386 nsew default output
rlabel metal2 s 207938 0 207994 800 6 la_data_out[87]
port 387 nsew default output
rlabel metal2 s 209686 0 209742 800 6 la_data_out[88]
port 388 nsew default output
rlabel metal2 s 211342 0 211398 800 6 la_data_out[89]
port 389 nsew default output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[8]
port 390 nsew default output
rlabel metal2 s 212998 0 213054 800 6 la_data_out[90]
port 391 nsew default output
rlabel metal2 s 214746 0 214802 800 6 la_data_out[91]
port 392 nsew default output
rlabel metal2 s 216402 0 216458 800 6 la_data_out[92]
port 393 nsew default output
rlabel metal2 s 218150 0 218206 800 6 la_data_out[93]
port 394 nsew default output
rlabel metal2 s 219806 0 219862 800 6 la_data_out[94]
port 395 nsew default output
rlabel metal2 s 221462 0 221518 800 6 la_data_out[95]
port 396 nsew default output
rlabel metal2 s 223210 0 223266 800 6 la_data_out[96]
port 397 nsew default output
rlabel metal2 s 224866 0 224922 800 6 la_data_out[97]
port 398 nsew default output
rlabel metal2 s 226614 0 226670 800 6 la_data_out[98]
port 399 nsew default output
rlabel metal2 s 228270 0 228326 800 6 la_data_out[99]
port 400 nsew default output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[9]
port 401 nsew default output
rlabel metal2 s 61198 0 61254 800 6 la_oen[0]
port 402 nsew default input
rlabel metal2 s 230570 0 230626 800 6 la_oen[100]
port 403 nsew default input
rlabel metal2 s 232226 0 232282 800 6 la_oen[101]
port 404 nsew default input
rlabel metal2 s 233882 0 233938 800 6 la_oen[102]
port 405 nsew default input
rlabel metal2 s 235630 0 235686 800 6 la_oen[103]
port 406 nsew default input
rlabel metal2 s 237286 0 237342 800 6 la_oen[104]
port 407 nsew default input
rlabel metal2 s 239034 0 239090 800 6 la_oen[105]
port 408 nsew default input
rlabel metal2 s 240690 0 240746 800 6 la_oen[106]
port 409 nsew default input
rlabel metal2 s 242346 0 242402 800 6 la_oen[107]
port 410 nsew default input
rlabel metal2 s 244094 0 244150 800 6 la_oen[108]
port 411 nsew default input
rlabel metal2 s 245750 0 245806 800 6 la_oen[109]
port 412 nsew default input
rlabel metal2 s 78126 0 78182 800 6 la_oen[10]
port 413 nsew default input
rlabel metal2 s 247498 0 247554 800 6 la_oen[110]
port 414 nsew default input
rlabel metal2 s 249154 0 249210 800 6 la_oen[111]
port 415 nsew default input
rlabel metal2 s 250810 0 250866 800 6 la_oen[112]
port 416 nsew default input
rlabel metal2 s 252558 0 252614 800 6 la_oen[113]
port 417 nsew default input
rlabel metal2 s 254214 0 254270 800 6 la_oen[114]
port 418 nsew default input
rlabel metal2 s 255962 0 256018 800 6 la_oen[115]
port 419 nsew default input
rlabel metal2 s 257618 0 257674 800 6 la_oen[116]
port 420 nsew default input
rlabel metal2 s 259366 0 259422 800 6 la_oen[117]
port 421 nsew default input
rlabel metal2 s 261022 0 261078 800 6 la_oen[118]
port 422 nsew default input
rlabel metal2 s 262678 0 262734 800 6 la_oen[119]
port 423 nsew default input
rlabel metal2 s 79874 0 79930 800 6 la_oen[11]
port 424 nsew default input
rlabel metal2 s 264426 0 264482 800 6 la_oen[120]
port 425 nsew default input
rlabel metal2 s 266082 0 266138 800 6 la_oen[121]
port 426 nsew default input
rlabel metal2 s 267830 0 267886 800 6 la_oen[122]
port 427 nsew default input
rlabel metal2 s 269486 0 269542 800 6 la_oen[123]
port 428 nsew default input
rlabel metal2 s 271142 0 271198 800 6 la_oen[124]
port 429 nsew default input
rlabel metal2 s 272890 0 272946 800 6 la_oen[125]
port 430 nsew default input
rlabel metal2 s 274546 0 274602 800 6 la_oen[126]
port 431 nsew default input
rlabel metal2 s 276294 0 276350 800 6 la_oen[127]
port 432 nsew default input
rlabel metal2 s 81530 0 81586 800 6 la_oen[12]
port 433 nsew default input
rlabel metal2 s 83186 0 83242 800 6 la_oen[13]
port 434 nsew default input
rlabel metal2 s 84934 0 84990 800 6 la_oen[14]
port 435 nsew default input
rlabel metal2 s 86590 0 86646 800 6 la_oen[15]
port 436 nsew default input
rlabel metal2 s 88338 0 88394 800 6 la_oen[16]
port 437 nsew default input
rlabel metal2 s 89994 0 90050 800 6 la_oen[17]
port 438 nsew default input
rlabel metal2 s 91650 0 91706 800 6 la_oen[18]
port 439 nsew default input
rlabel metal2 s 93398 0 93454 800 6 la_oen[19]
port 440 nsew default input
rlabel metal2 s 62854 0 62910 800 6 la_oen[1]
port 441 nsew default input
rlabel metal2 s 95054 0 95110 800 6 la_oen[20]
port 442 nsew default input
rlabel metal2 s 96802 0 96858 800 6 la_oen[21]
port 443 nsew default input
rlabel metal2 s 98458 0 98514 800 6 la_oen[22]
port 444 nsew default input
rlabel metal2 s 100114 0 100170 800 6 la_oen[23]
port 445 nsew default input
rlabel metal2 s 101862 0 101918 800 6 la_oen[24]
port 446 nsew default input
rlabel metal2 s 103518 0 103574 800 6 la_oen[25]
port 447 nsew default input
rlabel metal2 s 105266 0 105322 800 6 la_oen[26]
port 448 nsew default input
rlabel metal2 s 106922 0 106978 800 6 la_oen[27]
port 449 nsew default input
rlabel metal2 s 108578 0 108634 800 6 la_oen[28]
port 450 nsew default input
rlabel metal2 s 110326 0 110382 800 6 la_oen[29]
port 451 nsew default input
rlabel metal2 s 64602 0 64658 800 6 la_oen[2]
port 452 nsew default input
rlabel metal2 s 111982 0 112038 800 6 la_oen[30]
port 453 nsew default input
rlabel metal2 s 113730 0 113786 800 6 la_oen[31]
port 454 nsew default input
rlabel metal2 s 115386 0 115442 800 6 la_oen[32]
port 455 nsew default input
rlabel metal2 s 117042 0 117098 800 6 la_oen[33]
port 456 nsew default input
rlabel metal2 s 118790 0 118846 800 6 la_oen[34]
port 457 nsew default input
rlabel metal2 s 120446 0 120502 800 6 la_oen[35]
port 458 nsew default input
rlabel metal2 s 122194 0 122250 800 6 la_oen[36]
port 459 nsew default input
rlabel metal2 s 123850 0 123906 800 6 la_oen[37]
port 460 nsew default input
rlabel metal2 s 125506 0 125562 800 6 la_oen[38]
port 461 nsew default input
rlabel metal2 s 127254 0 127310 800 6 la_oen[39]
port 462 nsew default input
rlabel metal2 s 66258 0 66314 800 6 la_oen[3]
port 463 nsew default input
rlabel metal2 s 128910 0 128966 800 6 la_oen[40]
port 464 nsew default input
rlabel metal2 s 130658 0 130714 800 6 la_oen[41]
port 465 nsew default input
rlabel metal2 s 132314 0 132370 800 6 la_oen[42]
port 466 nsew default input
rlabel metal2 s 134062 0 134118 800 6 la_oen[43]
port 467 nsew default input
rlabel metal2 s 135718 0 135774 800 6 la_oen[44]
port 468 nsew default input
rlabel metal2 s 137374 0 137430 800 6 la_oen[45]
port 469 nsew default input
rlabel metal2 s 139122 0 139178 800 6 la_oen[46]
port 470 nsew default input
rlabel metal2 s 140778 0 140834 800 6 la_oen[47]
port 471 nsew default input
rlabel metal2 s 142526 0 142582 800 6 la_oen[48]
port 472 nsew default input
rlabel metal2 s 144182 0 144238 800 6 la_oen[49]
port 473 nsew default input
rlabel metal2 s 68006 0 68062 800 6 la_oen[4]
port 474 nsew default input
rlabel metal2 s 145838 0 145894 800 6 la_oen[50]
port 475 nsew default input
rlabel metal2 s 147586 0 147642 800 6 la_oen[51]
port 476 nsew default input
rlabel metal2 s 149242 0 149298 800 6 la_oen[52]
port 477 nsew default input
rlabel metal2 s 150990 0 151046 800 6 la_oen[53]
port 478 nsew default input
rlabel metal2 s 152646 0 152702 800 6 la_oen[54]
port 479 nsew default input
rlabel metal2 s 154302 0 154358 800 6 la_oen[55]
port 480 nsew default input
rlabel metal2 s 156050 0 156106 800 6 la_oen[56]
port 481 nsew default input
rlabel metal2 s 157706 0 157762 800 6 la_oen[57]
port 482 nsew default input
rlabel metal2 s 159454 0 159510 800 6 la_oen[58]
port 483 nsew default input
rlabel metal2 s 161110 0 161166 800 6 la_oen[59]
port 484 nsew default input
rlabel metal2 s 69662 0 69718 800 6 la_oen[5]
port 485 nsew default input
rlabel metal2 s 162766 0 162822 800 6 la_oen[60]
port 486 nsew default input
rlabel metal2 s 164514 0 164570 800 6 la_oen[61]
port 487 nsew default input
rlabel metal2 s 166170 0 166226 800 6 la_oen[62]
port 488 nsew default input
rlabel metal2 s 167918 0 167974 800 6 la_oen[63]
port 489 nsew default input
rlabel metal2 s 169574 0 169630 800 6 la_oen[64]
port 490 nsew default input
rlabel metal2 s 171230 0 171286 800 6 la_oen[65]
port 491 nsew default input
rlabel metal2 s 172978 0 173034 800 6 la_oen[66]
port 492 nsew default input
rlabel metal2 s 174634 0 174690 800 6 la_oen[67]
port 493 nsew default input
rlabel metal2 s 176382 0 176438 800 6 la_oen[68]
port 494 nsew default input
rlabel metal2 s 178038 0 178094 800 6 la_oen[69]
port 495 nsew default input
rlabel metal2 s 71410 0 71466 800 6 la_oen[6]
port 496 nsew default input
rlabel metal2 s 179694 0 179750 800 6 la_oen[70]
port 497 nsew default input
rlabel metal2 s 181442 0 181498 800 6 la_oen[71]
port 498 nsew default input
rlabel metal2 s 183098 0 183154 800 6 la_oen[72]
port 499 nsew default input
rlabel metal2 s 184846 0 184902 800 6 la_oen[73]
port 500 nsew default input
rlabel metal2 s 186502 0 186558 800 6 la_oen[74]
port 501 nsew default input
rlabel metal2 s 188158 0 188214 800 6 la_oen[75]
port 502 nsew default input
rlabel metal2 s 189906 0 189962 800 6 la_oen[76]
port 503 nsew default input
rlabel metal2 s 191562 0 191618 800 6 la_oen[77]
port 504 nsew default input
rlabel metal2 s 193310 0 193366 800 6 la_oen[78]
port 505 nsew default input
rlabel metal2 s 194966 0 195022 800 6 la_oen[79]
port 506 nsew default input
rlabel metal2 s 73066 0 73122 800 6 la_oen[7]
port 507 nsew default input
rlabel metal2 s 196714 0 196770 800 6 la_oen[80]
port 508 nsew default input
rlabel metal2 s 198370 0 198426 800 6 la_oen[81]
port 509 nsew default input
rlabel metal2 s 200026 0 200082 800 6 la_oen[82]
port 510 nsew default input
rlabel metal2 s 201774 0 201830 800 6 la_oen[83]
port 511 nsew default input
rlabel metal2 s 203430 0 203486 800 6 la_oen[84]
port 512 nsew default input
rlabel metal2 s 205178 0 205234 800 6 la_oen[85]
port 513 nsew default input
rlabel metal2 s 206834 0 206890 800 6 la_oen[86]
port 514 nsew default input
rlabel metal2 s 208490 0 208546 800 6 la_oen[87]
port 515 nsew default input
rlabel metal2 s 210238 0 210294 800 6 la_oen[88]
port 516 nsew default input
rlabel metal2 s 211894 0 211950 800 6 la_oen[89]
port 517 nsew default input
rlabel metal2 s 74722 0 74778 800 6 la_oen[8]
port 518 nsew default input
rlabel metal2 s 213642 0 213698 800 6 la_oen[90]
port 519 nsew default input
rlabel metal2 s 215298 0 215354 800 6 la_oen[91]
port 520 nsew default input
rlabel metal2 s 216954 0 217010 800 6 la_oen[92]
port 521 nsew default input
rlabel metal2 s 218702 0 218758 800 6 la_oen[93]
port 522 nsew default input
rlabel metal2 s 220358 0 220414 800 6 la_oen[94]
port 523 nsew default input
rlabel metal2 s 222106 0 222162 800 6 la_oen[95]
port 524 nsew default input
rlabel metal2 s 223762 0 223818 800 6 la_oen[96]
port 525 nsew default input
rlabel metal2 s 225418 0 225474 800 6 la_oen[97]
port 526 nsew default input
rlabel metal2 s 227166 0 227222 800 6 la_oen[98]
port 527 nsew default input
rlabel metal2 s 228822 0 228878 800 6 la_oen[99]
port 528 nsew default input
rlabel metal2 s 76470 0 76526 800 6 la_oen[9]
port 529 nsew default input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 530 nsew default input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 531 nsew default input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 532 nsew default output
rlabel metal2 s 3606 0 3662 800 6 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 22834 0 22890 800 6 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 34702 0 34758 800 6 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 36358 0 36414 800 6 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 38106 0 38162 800 6 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 39762 0 39818 800 6 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 41418 0 41474 800 6 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 43166 0 43222 800 6 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 44822 0 44878 800 6 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 46570 0 46626 800 6 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 48226 0 48282 800 6 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 49882 0 49938 800 6 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 51630 0 51686 800 6 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 53286 0 53342 800 6 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 55034 0 55090 800 6 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 56690 0 56746 800 6 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 58346 0 58402 800 6 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 14370 0 14426 800 6 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 1950 0 2006 800 6 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 41970 0 42026 800 6 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 48778 0 48834 800 6 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 53838 0 53894 800 6 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 55586 0 55642 800 6 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 58990 0 59046 800 6 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_o[0]
port 598 nsew default output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[10]
port 599 nsew default output
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_o[11]
port 600 nsew default output
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_o[12]
port 601 nsew default output
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_o[13]
port 602 nsew default output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[14]
port 603 nsew default output
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_o[15]
port 604 nsew default output
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_o[16]
port 605 nsew default output
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_o[17]
port 606 nsew default output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[18]
port 607 nsew default output
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_o[19]
port 608 nsew default output
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_o[1]
port 609 nsew default output
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_o[20]
port 610 nsew default output
rlabel metal2 s 42614 0 42670 800 6 wbs_dat_o[21]
port 611 nsew default output
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_o[22]
port 612 nsew default output
rlabel metal2 s 45926 0 45982 800 6 wbs_dat_o[23]
port 613 nsew default output
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_o[24]
port 614 nsew default output
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_o[25]
port 615 nsew default output
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_o[26]
port 616 nsew default output
rlabel metal2 s 52734 0 52790 800 6 wbs_dat_o[27]
port 617 nsew default output
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_o[28]
port 618 nsew default output
rlabel metal2 s 56138 0 56194 800 6 wbs_dat_o[29]
port 619 nsew default output
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_o[2]
port 620 nsew default output
rlabel metal2 s 57794 0 57850 800 6 wbs_dat_o[30]
port 621 nsew default output
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_o[31]
port 622 nsew default output
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_o[3]
port 623 nsew default output
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_o[4]
port 624 nsew default output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[5]
port 625 nsew default output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[6]
port 626 nsew default output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[7]
port 627 nsew default output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[8]
port 628 nsew default output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[9]
port 629 nsew default output
rlabel metal2 s 5354 0 5410 800 6 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 7562 0 7618 800 6 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 9862 0 9918 800 6 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 12070 0 12126 800 6 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 2502 0 2558 800 6 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 3054 0 3110 800 6 wbs_we_i
port 635 nsew default input
rlabel metal4 s 4208 2128 4528 237776 6 VPWR
port 636 nsew power input
rlabel metal4 s 19568 2128 19888 237776 6 VGND
port 637 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 280000 240000
string LEFview TRUE
<< end >>
